// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 02:45:30 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VU22x9Qx9dSYErajB0Fx5s+8mM87dUzuyFi2MXOUg5YrEOfv9qXksVz/bChDj9Z/
KzQ2eLYZlsLWnHUV7lQWfShAzT2m+JU4bQonRuim6tTbP67ZJrPEyXLpPBtsfr/+
8ZHxrthfxpEG9RIXUQTncZ0VjZF8jJDNfEoT1pqa0m0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1429888)
W2sGDPngcM4YatjqxgKuSHe0+caDagMIrLN2O6xwoyx0VPiOi2XDAH5OYozpponq
bjjZxQCVYcVCfw6HuQ5moWuWneB7IFxZe+d7r9LZy4Jne2d065Z92YQqM5fZhMe+
FqChCc5jfOqL7RSG+jM1GET19jmbHFWFY2xSVEmt32kMkuPau7cklJHDcnw1vDep
/mg6YypW4+sKhPMIcTldTIrxFPEuTHnBF35oASrE87sKnlkUTAn7RN/H/zJbkpfR
vG9LLAoUUnuf6LnHuSzmqQFEr/HRSz+UBeL1rFmiRKIxDUiLzqYXtjHstf7sYy9m
v0yseE2ZA0Sei1I/UVYOfNu9Uft9nnHRsUeWWEagyUpzvTjq3HWsV5OJ9zHJMQVG
wRogocivARZGj0yUlanRDIT3iDyE3shbc0AF0JGBnzwD2wqG9y5gJlQQtqynrRfr
XLGtzrU6wIKdp0WfUZbP0L43zzvy7nodva4GO6NZpVLDG1Eogx14xk3AgyqpDtev
vw+SH3v0wjWo/8TPi9Z+WQK8UtqYPLnBo4jPC6U39n9lP26Q0QPsffsv+hWHGTEt
1H6Q2kuXM55oeh9Li1ix6Voe+SaTjE8aVEyiICimdMQh99c/S0+q42KOsmNe1l6G
pKRBZ2i4cL8j61/lr2hH0b1yBgSXhrgC00AJRw6rzEchqpOgw+NtUTGRNz1d9IGL
T2XI/c+ooFbonOnBctw1QEOlnBP7sjePm/5z2tkB/GsEfc8/vndJUfDrtWddOsbL
tamSxaQ8n7dqGoWGT/5NiNiq++y+NIxQkVCFybGYVJGstyf4y8cLokfUpxONq7MI
oWpNxqLXpQAizxO/5LPiJ8qWMQ3b7fTjHeiFSk2PtnkUdgiF1gC9XcA8Pto+6XuZ
WsJHKDI37BR7CVQVg+GzcL9F/s+rxy5J4DrETVvkDXoZ2KVh6GxvlBtupY7MxQeZ
hMA6d28uW6rjFk1YHOIxqH4MTzDGRf0zQVlNfzGh3C2JND3SUPNZBrkLxijZwPdw
GekFH2PW58dcSQ/lkQroKl2zk6iybxwzaXSGEtYn/wBXL0vkPUhAhxiOOp/fGnwd
kUDKQawYajcDGj3mOt1U73G7ow39UvON1/dWbdgVJoboXPbNflE4ZGLBafKDl7yO
pcnvS69JGHRqzkq7wf23XV0tFVL1b3Dt9dDItRfvF40JsOAQQZJzUcLD1a7i89Os
iBVquPZfNrb22C9fw+6x/82SiZxi5saoyL4KDnh/5HeXw1IZqO6JUeq7m/zflr8+
NZ942oyZSWOt6pX5bI90t9HnldhcUSSvBt5/sc7bFz8Kw14cbKjjutSkBTjr45+s
XcgkmP5Tl8k0N9Fv+UNBjPSfgSTN8OfD3E+x50fHfNwdMhHCMni+ok1qswCgYdU+
Sq4KejeZWP2ovbLpnfRO58Ezty+V4Kuf3lUKrh3L/zxXBew8LaiqqfzmmF5R583m
dVkw6BM91j7zc1QxnpQbQg822qrwMexHcLprVSZg6NCe2QdwcBsFsjcaHozIUvSH
NR9coiYtndSgMj7oK4n45qW1FplTqJZ/3Hocj509D10LqCNyAd9Nxi2YDdkwYjON
qnhr+/Nc6WyV9qVEH+dtSinXVXfuqi5EkWAmVa+OPoWN/D3QvCzQoiC5C4+/ZDk8
ZA67XQUwP/GSHpRkQMHgOIkYonJ5OXzKRPaW3cxrFSM3yA/mhZaVGudnoBWlKQjz
Knn3V8IrijhbjqnNhNe1H6AlsQXIp8wOvHUgtldI3itZ12emC6SgZsmpOUgNlrTF
UPKDpJ0xKYvdyLrFmB0qFvCCrZIsu/mDB6y/jbSoluzeyT2qBdqD6VlieSWFmBu0
VVv31EScVDl0sOYpJrWCEKuBDnFLGqMKaxoquLYargwlKboGVP4H2IuDRo/TXQnp
fB5IZQE/yQD5992I6356Asw2IGOuqlAEB+FrJAC4Qlo66U7RkFBS6Usl44PngryD
Uk46GSJIqOY5uK/ncmEUQtn5McfncCQPObzTrXcrC4VNdivtAGwtcC0hTQqKXyak
jyNwvFnJ58jji1DQlKnJgY1vikWAWUsCdTIWiOo5UKPwTn7w26uuEE015Kz88Lt0
b+suDYYkRfh8qQO8D9U9IdTSkxYrEZRkIohC4fvLYcZAJHEwgQ96q6f4QoZM9FMP
UmNWNMZXQA65SQLMYwX+Q+mv20oF3wHma/8NqU7cOHYsYxV+KRFisJjbiOb3a+ej
r+NV5gVTB4L1Mljlykswr7a7JYVp8PPXpN8bh+7n0PY4OpTgjmAV7AwpWWtBm3qE
0GTXZgBEPk27Dp0qVahTRqcq3wYIJzAPFt79mlwCY6ZJmc7w52c4IlNppwGzrC56
+zxM/1hSSJ9UQWj3CCkkZF9tO/ESs2BnKJ9ThVenudcxo5rG+kxhCVayIixW7US8
J6knwfRe//o38D+LUdEnfCUGoyM9RcuJ4V19Nfpu0Fig7/BFKJZBXD+rL7A+rPDa
2X2nkRcH7hYZ3DQ4ekyAILekpX/t0LB8vCzS8APK7lgdkqh1F5BRCp5OWPWi6xvG
q9/fkRJXvwaKPFLg47CRN2U5KYN06G3B/H5XgZ/xSkHJSW+LFG8BOA1hSXUe16Yl
amrNDQJpeqSo18FGeF+sS/qxaNthOM4mbCgAGLTRfISVveoLHd+1NeUTnf7tcILp
zl08iiyHipIThhFK7g7R78DX+qg3jLTAp8yzTJK60wfWPIAVOvfExSkI8AsZbD5X
D3ZiVeTpf9AwGmAEO1l9yeSZuMX7uRgtI9TwAD5QsMUJbzmGWBenoyUI6PYnaYSG
ChG+1hhfcPArd627aX30ie78L23QxgQl6L8eInjNBdzD8ZG+s7r7Su9XbBllZ3CY
bxtsDsrRC/XFaTpmHVtTkPKgqXj8rMFRTqczhggDU/liYQUaFP41TyEj2Q+EUa1i
YTz9gra833uqb9sIyuuga+jWxEhuwoth4qvJYXGgiMPgjt7NyfWG/JTFGcHXqEqo
GkhdaXKlShnUGI6JdFbbVGiPOOK19jyJRneM0OmZ8jz7f58A+w8SeDYxWybl74ak
iUf7SD23giO1hbFJW+zcxGmi99kmkEb5TD3xClFuBMM+EEoHgM/8HMmC8p+iCy9s
qL7jgfnSHBE7NDxHI79EeC8OzSLCHaXzrdb8dQvoPDWYUTD1RCYvOLMpKjVmqhbZ
SNqDf1TSDtlMK9pVZN5ONm94L3AdEGsJlF9ZQBoHGo48U7tBIxyOn5JYDM/3hrEo
ZR/sMrU1C7hceYtglkNeyX6tajSrFJf33rO3ZfHKyymgn8u7AbUJ1kE9NBRWDsrj
iAhbK4uuYnnujRHbQzej7dEKTDQEiH5BFcXxshF7zD7kbnHbtDgnUGPhgEja2HjP
A4xYVL0bffYFlFOLpj8lHA6T8YPtfnFaialDnpseY8/tdSzCjL/bDtyzRnFMpn8j
nCHHAQIJLdQeISL8aVyEoFsMHZLLzRDnQwiZWRsthCO+vF60r+aWwQEkyhmWZ6Ch
U/koyuEqYuWipDxBptrsSOvsfmEvdsNiCp/5GxByo8hTnHne/UjhGuQLLmF0agkR
yGIipsf4urikuArmfP/iWaYOxCKsHkV6yU6bOd4MKrBQ5+p+pH8tLfm1wn/TyPPX
o/Az56E7JY7jCLR6X8U00aP1IkBqADS9KPTM2VBRfDl8V2St2Mq2etxaiPGVwHtJ
+nzCJqVCDhzUdZgw+mNjZLlcPq/nSOA+sWukdaCS1+A8sHKQC04bxxw2UaADk+8W
skHT6hKaT/U6YITSw9i4IVDZGBatpYDo7uFABxrhgipKFMhluw7PR5l0UxJXdQHp
PfPPleOTOZdX98v+oHPdhmjYpRT7bsAiU8Bsp/9BogJD7OfFtYH85Dvba4Xaf60x
saJUi1CdKvx4H/3NPGYEj93XESzS4O+LNBheos+h8tjKIIv0B+hqAAz8J/xQu5d9
OYDkziSDksqLhhz30KovCbp2ts5CiwhKEVxA8lKngl30YzT5PW7HZN7Yvyd4vzjr
Q6QKNd5vhazWoE276z7pZHqLZdRlluvXj/idGBEby8+48F0g3tuIuaU2Mr149Gwl
le/c/KIiEeHISC7T1P8X1lpgMGYMtUupcN0FTGIDx3z7nzHoN+TVweccwHg5fSpP
EBm6vKY3pRSkEjvhfGfUUpGX65V0XIBIrh5rpvAuG+52CHvGbUxjW2vLGgaNcilI
w7CScnuyObc9xoz9220e1TSaTiya78mBP/v4SYCk7iohQlu7AYcDvp2+P88fRCZm
qQ97Z4zjaZXlHNVJwuybuazzaF6M0QkDYsIMpXUC1FQdpQlO0q15vWoL5nhgog4X
CLMpxm4ojxFjbnmNrQD0QX5zKkaWW0FLFsNhc37tgRubnJkCajcq4cczeTdYD1Hu
1fDYv1RCeu+h/AuZhg9GFFKNP0xVmn+Lgz+RpeiEgHPGqnh9coqQQmiCU6v4pN49
s4kcgId++8IqRaZQNgJqEfQzUm0jyAy0F1+lpU7gt4DnuHf6zhXq5Tg+2gNbwAJa
0/TpQHUFfpK8bGo0R7yGptaItAYVvqzoV1H01aks9HUMCm3krO+QLaPWGgfiOu65
sbc48sHmvjjrfFviMpcb4ugcJKm+oEaieWbfxZfwuleaBjLdYeixlnvLJmPVzAvz
iGKo9dJ3zdYQ75GE9VVF4MPWsNxR9IqB3/Y3XF6zhYuXFFeZK+4e/r9tFtsYJJdU
yIyIIJwnIl6qOSDaosFqn/dOwgRBY8KJmIz99+kC1EvUbWMiJrieu+uPwKLJSzkR
Fw510w/xcPsa/XOreIHxm+H8rD4GTLdQcxj95pH66awEb0M6IcFGXXhTdeyOELWW
8LKC5KoXJJ2P3RJlWWWBzbv4I7tb+dYSmL3RGNbxOGDF/lHOPUgSuCUdvpSYNrZe
d5XCOOCouQaJxmmHUFauA8quoZgRESmBudTYVCh5OXsAiXwkzX92fxeR+7qgvYXL
bdXjsJBjRRdTPJUXWcUEJ8Mmlhf006JFaNcRNXKHkdSbUZCX0jULYAbUbKrScBlc
PXCcSFTqJHQFNFeU/lhcNN1SAmZUmsV4vVIyfVZY3vyBRTpd89dKRK4H/BN0o5eQ
IzjCCJOkt4cn7h4btGuwOJaX2lhn836KnCHrE6Jb72mhWoPmm+C4mIjM0HrbomTU
wYGtYdpvbfa7BPa9BtSRG5mzLicRore9yRlgadkuu8P0K/lc1XRXJMjnkqmy82kJ
gxJPWsjZJGpluyuO1M2wp9HFgQ8X/vVmx8OhEK9jE64z/LMSfBhm8zBglmIm3ADF
fXGm3YClms1uzUw2RUz8RtPIPzb8NPX20wOBL1YjdR5jQpg3cHvA1Sbr2ISFy8A7
6/b/Auhh9cSjwGJWjT7fu9DmrCrI+/TiF4XCBej0yncrGP0imgA+o+zBDgWopyss
Ktw2V4y/5ObZ3KmOR2wZKuHofopY56eMmaLNV8dTGWvEna1n7OVcGB+KRUDk4fnw
hLwas+bvEqwz5cfMhpqKZuz0vSxz/yJVyHJ0UUtypRvg9en5DlEZCcCcHVjHTzCt
yLHf4ooLg/B2kbYdqOLQUiEa8Mb0JGtJ2sYOEtT6aGIP3P+iVo1qL7vj9igbqC0q
33ET/FerLrnorxYf/e49JpiPPNeR00T8bILVwQIk+B8OcX4bCjo8pK1XFv+Bzxl4
ZqVhQW3vuMfShLWtICQgw39d/D17KJ2mSo1K7dPIsFSs7qwV1pGhmxGgmR5tUmsu
1NVmgHkXIT3K015KQ+1aQ7FG9+PKZzj9Xjkg9DvgkriAO6FzEP0j4LtH0oMZEcn5
jD/g9Bj/Zl016hZIZuzs5eEb6hKdnxZCQXRlEu0hb66ic5EusHDJhYdCMoPrgNMf
y6Fg+wtaW8Uy2f7Y3DMQG6FcKRU5BdQIO+moBcXsZeV6kPsx490kNcViZdqNNP6P
67f/Ujk+J8ArbwkESiFTfrAShQkgKUgOutcRgM5oIqbTOH1H3zlNEktJP24Zqrh2
o3wH12xbXPBEpPxoCEAJyoFZcxZeSMRR2bVfCx5NRLJu+vXhdRi+3lTXqcugAJVU
OXPn0+6mhgQ/PrmErBItHkRQKdaL2ecjeHs3bbKLeS/r3+AzZ1sWx/mBrE710L4b
FQlnQ03XEYJKORUD6RQxjctFh9FlKXeEvi5zHjGdfroXlEuVyVBb2dNjMX1/6FKu
FIFY6HGsNv3CJTdxmhFJ4nGSBPx8hVMZ7/H/inArQ8YiHBgDAWQvAHc9IiqyWFe/
aVOz3BkKtTHfqarnfjgYhSd8lr+VxrZ8+Xz47EsFECoNx0+/3hxF43MA9L1BJs0k
HXkHIwE7+El2QR2BkSHwzuHNs2gyJ0wTJSlxxcgfTCzor+SRQa5E8dmtNCKYroBu
0hTk4c986Wjzu6xMJ6BKN6EfgivSdASeVoI+70fT8JdgVooDMkWXQB7s+hb+2NLG
kc9ROv6OUh9Ybk2S2TiMtgfk57Za5QzEXB/MrlJaqdBotKUZhCaz5CDoj2oPCAia
XGoGa8PnHpTBAp3Or3Wtdygm8NvPbMfm+a+1FJlXyStU0nJCrHwuU8VQrD5m0gxL
UQBCeMS8Rym7TpXOarDIHdx8+jZeBTnn/7orgubcy3XWkIgjXRKJPym5+t767DTk
ajnG51MTLxq1hYbbh12P6hxNA2XtzIAKyxCNWO18A/Rvx6iI2UjidksB0Lk//vr2
4fSFeKqCE9rOIuh0KD2YvoyeLb1Vf430nWKNl71QsO+oO9t3iUPGlU+nuhMQ7c7r
O9fJUNnJcGp/QpBc9IjPMgtHiMz1q5uk8bSlvm7PqzE5XWZxR8wMvrigRHJuRBKo
bTTot95CPY9ygdPNXSCKTkugD4eCC7/JGEWH4w7mMyoM2hwtJAQtAVhNlyR/4p1l
VheA5ZRHV+zCMDFykRUKFtQCmfS3osWgu/4znWdhdSRXaq5sUT2/EYBPRo/aLVQK
f75C/UqCwso9fogJffdhVdf7xM4PgxJqWNDPpquntDpXSDPNQAlcrmIKCt1ONfke
3LqB26lJAmdQ07RDtp9CSG5ftuSQqt3rQj3YauENkd1H690z2MY71LYYDEW9S+4G
+EgiLjH2tqbs3bRZN7s85p1A/tU5cJ8ShQfD2L7hcFMjnTjnVT4291aS8LzGJpEo
/Acr91FFMVOiD4QCltmjA9iKlNBopeEEumNk7EBvhEld6cjwja6/c5tYVb6AfZyW
qCgfvXjFwHkbfEJxLEOpzZ66b1nnJAPUKKvQ3KKPCjsf9YsOpy3UQHVndSmVdr5u
96twtx6no7VqigWN+qMRzydYmAFfi0Ns+2HlUtiIUf2/7ATagHeeo/16zRojT74R
AuhiXoMvadmJBFvFg2xQWVuzeiAyRzIa4b8Rbhes2T5ldtHQIUxVkyfwmqwW7z90
IJ7Fc+ExPwXCKHlSUlsGMwoU6GvtTrRX76YaoqyzaZsATWsfQEDB/7EAPw0OZXlq
pz3L8wvLWO5PM8yLA0uzs1gWYx+IF/U/KKeep2SfWvdPFWlm5UBkotRryJAdX8Jl
3qd5VLoYrI8ZZiSu3KUDamJ2F7yhQ5jZ3UvmyBEqwOp9/dF8DknX4+k4knpXsiZr
fV1UEhl3qe+CleEVJ9t6e3HGUVnxVzZ+6F2sRu61O3Pk+e8UzI7zqRU0TKmNxTsm
LRR6+REMNLYNVWipIdn1zvpQ+BK8qkjLeSlNcCoP8jFnLuEsOMxr2XEBH3bri+W4
xCRSV3G/y8yMgsXL6AaEIkl6SUrPjNkOnhTaQDPBlVLLXAvWFTc6wXTzCDdzpJGZ
hfZnkQc/gR6PbOPwK7xqF5nTisA8kV0PBomTA+apZjpj/akHRwR2OuQnETGQ0mEz
QsYyxkcv3ccfPJS3Mh/Q8rHmPRcpwpL0MQJbhuXbn+RIRj37MZ3UEb5r6NXj4rQy
bAY8bM+T0+5G3QujR2JuWWa52irlWiCP7ePLwbYmguzQY9DvoqxBWWDcV27uJYNz
Di9+rS6F887QfzSbeRoZOXPk76f/3bQVrZ13rj7hOApq/aGLjYlRStWAo+eVfl6x
PkkStU861tktaQlo3+0lGfiMUH1oYMKmd0VmFWVtoDs/X4RMikdj8adyotC8xVLg
2emK9pVv5ROzHpgm8/0t4A1LKaNHh4OD6QF0DHg+6q9nI5ejlYN9FqpBrGPCt6ie
mgg8v/cX317mvBBmUsMLZYc8mNZo0aMcK8CRBJqdqD5ouRr7edxrwbnMr+gTK0SC
2qLLoNx+SE4yEW1h5C/wpv5vW7hb0c5hDD82mUdks5SoDVjXpc2jHeP2UPStfLxV
j1pKyBfXfyZT3/ngNDPUnlVB2QR0CJz6s673RSlZ/tNciYYUBkNhbVbcw6SdbZ8B
SA4c/+rZnlKam7iHwDNF0Ti1CI3CXsfvjdiLds9GeOGVyg3RGcBthUh78pkVtlPE
q/SLqz4GLoPoY/yESuZt5W8d5KMQ96BTQecuUBGO+MUJHV1E6BKFJ9lB4gVX3vAI
FkQc9k4OwkK0NHsLKD0uMBfiu1Iwvik321nx+fmkDj8sM9kk4pFa5z0Iic8dPhBU
KcV2/9/8OjS1uM+s5K0VV3qcL8D26IX6NADlw0rBwHEtzZZrnlxr8LX2AVGoTp9t
2s+/KQX5BNMS4uhRMZaCsgb+1WOlSWr4zl3/Yjoqov6FEo5/0+QsIYchIw/T1xj4
WKuVqReXz29tzymDedzUTJyhAhHpA1Q14ur0a9mSLna3IWFBMCnadkyyUyYp1mlx
eLy0gFo29FE7G6Tlpf1Puf/mC/KHcMuxMfEz9f6qDrEoCZcfiyJnKwI6WkWZEmGk
vTsv32DChoGBIY42YZpNzeUtojm5ALYCYpMtbLA5sYYlOuPOFZuMzLoIkDLCzniB
rZKk+uymfcgizUIrCF9HptRcoZvtxX4pKMRG+mjqzm4sLjRd0YWD9FRZnCbt5QLW
+QalCe3ai+Nf69gVJsRpUBZC1JEesNQ7Vy05RQlCXkIGTJcWQGZzPHumW7KolLpi
TJI6SjO54ehu/koR/iBjyWuYtenUl2TdSSfumBGvEKUuzn1ZUTXyFHP268G5PF1s
H5LOS3zm34cqGT5MOW9lNfmhbO2CdRKQgyb6k6ogdI0YgZEuQjIKWg8vBjnaHCLB
7c9cwD/SpABG7xe0BAzIDDK9Edn1NAfQwLLYFQr9ra9nFXwKikETauGkMTGpVhfn
uo9UstgDdPassMxZLBkFrE0hK4f6Wp7dIgXQVu142om6lVRo83D6uHMUiuUm83FV
rSQCCYDDFFbeF/XlrE1038yohO4NZaKg0eO6p6WT4CnVb84YuJLIzmLnw4Q1SllN
f2sJ5ok4jGxLYoB9PHAvAAFoeDPMksZKBHx5cohdTRo1U5aFyRF8ReHgomTL4r0f
Yh3IghpvHCCnsdvhgkVjcs5rLZyykI6EaZqNpJiYK77g3DZXL1SKHZcrkd0iIFbe
aY23r1cNZmVzcm7XHGO8RNHh81onSBQngBgdBUAsEzlpXu6vfKaZnPtiIyl93A66
Pbc9hHRnkgz+5+dbwI9LT4/Z9Vcu2RazQX4OUNd5E7mIH+qWbxJcCDn2i1qkBksS
KAc/VbNhgoDcb74S5sOaDs5I9f1tkoWAGWmeObGuvqd16Bm3T+2NDPSR0ebG2bPz
uCe1GFNGQhVwTxszrMGvY0xgEAd6pKQInc+7vklMyRcwcO0c0kaqCzW4CAJgKVm9
yRJYVHrxZZ+NKFdJD85lci34ulqoO3KStxZjueYGqAO9WGulk4unfC3GyLnD/RwK
9QB3iqZR/0sNdldZHZk3zPFck3TYyAt8ZaqivOhDUMZ5omUloY40So6I/jVQwidx
GZB0lDDFnEJ2bJ2659G/8kq7TF8ICwcfF5N68R5rzs/SUJ8uAtzyH3pb58YaxIrI
XlX3MY9TKF+ZaxrxEKKBBa67REgDDLZPj3ZBmDajvP6tieZYUxlawpO/w5gzHC2l
2ySA7OOUUy2qqLSM6Lf8wBvzpQ6QvmGElZLcp0Bo8GL8ljQKwqftVPGp7kG//rZB
0uPEkQtY2dBPwOJr4/F+xCYrDSP1mkjiF3JTs8DjwoFGRr/CSHejszxJNUoyN1Wj
mrDzbePuwJ+011znzMYXWavEqVHURtRl9xBbm7BpBl3dLTazlpbyuGptRunP67KY
eSIAYgmohkjP9RtrtNkhVnomGqMXPv7v+tCc1lEq4gqXAeLN8qMLP0vBEXTqLE2Z
m3S5kpP/RjNHsG2P58+eflWTQPyn7oUnklaQJwAhq8bigcDBEVZ4U8cWGK7lMmnc
dqKSrt7Q1w+IJrwQEqqcTXoxDmiP/INB3rruHBxAM/cDLOpxbCergvPXtViFwBxk
ZNc2ZEKq0lNQUjYY24b80ltRtQ+rT4KW/QGzHpNj4c7EZspeoHtbzrFhECl/5+tq
QjrOmO3TU71i7iDfiWwSBDA6qtIWjsz2RviWvcO0RHBkBMp4tx5pszOe8B7z2N4l
DjM2ys1Oe1FJClIPLt+9uKfEPkuyjHk78j+LOfsEUkzqxHysaY3B2to3vTIduZwL
is02YuiCw0VNYlmrxxKti5aNnElsOmlUR89Al6glsVUnulGHhKsON49Q974Q76Gn
yuBjZW2yBY0PgILzVr5OP5I5KS3SqNI0RXztDsfzQA29dq6QGUkO0f19cj9EMGFI
SkvyLX62+nRQaKkulMMIOWAT1jT9l0N1XCCYUvB7vCaUnIH3u3ub/nzU7TRVs6wH
utAZceBmxgeH7T1vRpZxQvalxzOwsmw0suJm/U1lMnVEL86lZuZ34xhBececMKQ8
r5sfG26paPnEUo9BHAajfhvYrPBP88aOvyEyYDjNUmjP+94zEMqsXezThu0L1geq
NMVTDKjnb1S2GBB4iOL1inBfoV2HI0onhu5B7zqf5klnF6UDfg3oDEvj7bp5wk01
cq88/AteA98N0g8UXCEFxIoqccKDuWyZ96DIyGV49OaC17MawC+vhwPPO/hnUE0U
VqpZX+Vpj759wWueB3bv2gvZV2k1RXeJE9uWk9gqQxyLPrDxpti0NdzYki2N7ecE
y/rry6jGaJ7fzF0cpShM1crxZnu/s3I5M/rDQvI0YDjGO3XoAWARfLkAwdP1+jfF
sLUjfU2Z/8kgN2QRSTkONqKh6zfntHvY7lOQG7xdwoYlB31070lwKylYkVhLAZ+7
NAgNuBfQGsfBSWgL8Xhwwd+pA8h3iFIcnESydgJM4N400vsLdIGrNzAo0T0bsJVh
dC+cg0/kOfzq+xnl41imcwP9mKTPP9caTwb2jmSviA7omD853DqiLs3l9ed/BEFQ
LorB8m/c/wdGT6Z1Uu3fj8ZNrVUDUs6HNufHGhv7+2WO6oJ9HBY9SmrqE3lYm5rc
6Jy6EDKmyvGDhYRxOry1lLSmxOSBlHUUGKyxQcwQ3vKnyxYTTE/sBwYURdQ8I+TH
qNt7TW0QF83eG/NyAT0dSM8gJ+Athxis9Hr22eoU4KGRvOlJHXY0+5nNtGH9dqgI
6c6ZwKc+hOJhlr/q9sV7INIRXJQMfqSSJ4TDPbHKeUKVd9He6VDM0tx0YNa7JC+3
Y5QEE4RA8RlXE6/JMV5u4wgP7q0/oH6Ksp8Qexopx5jso7OrpAvbWTK311Xw/VLd
/L1gZaCeyRnwwsEwNSGPm5zDhEH6N8gBJ0z58vMJ5+VVRJj99MM9neitoNDK5avI
bBcoTd++yp9YoofvV2UAbt45zo3cUT0jWfdhw0ypEw5mJDIFb0TOZdoDeCmb04SQ
Erq8XHNp/+hqJUDSfO6iY92P04Pbe++2XXfxEn62FowgQpQ04YC87Qf+XSA37HIE
dj6kl5TKR/3B0OzPkjEAf9+4gYXb2sqNTArhzqbvVJJjo3Laemj3kE25OuFSI0i4
DMG5npVDySCwvYU8LcLRob+pS4XMjkUCYhu0zmC/LacKkxxMY6pcMhT1dSBpS0n5
6q+BRH9DtsH/feKfJ78ujq6nf4Kt9YbQFy6PbJ5ysFp03IyHKefj36dGQS4EQZ+W
9Serh2DBOeHLxHmg72FCtM8Qszc5SUBrDrWLoQIIXkZyabHOwHSnxcudUyDALxUw
zKt9yOIYyDOzuTfRhaC5R2Sc6rwJOA/fZYqfdfqwALksDpEcwzA1nV3gVtXdjrnY
U1NvhA1aQVDofjzTW96L1JqeoJ0Uh9d0XBORyIz+2DX0a0k1ka9yH15iDbcNPn3X
xskN4Llm/TibBzepqci3cVQpnoNOi0FKA52LfEyE8U9UjkFXKcntKVF1f2vCuhs6
ShRO+qGeQhsx0nOFmfaxOnqcw4LJYtouPyhAKP4QpHTgoNskl4wfl3GkfGFKW/fN
TrQ5pu/ZUDVHhPD+MRir40vMBxt3duXgsvJak5ukuHVK5dnK4xAVLp3PUZIaIK00
TRvAPllsbUyc/ojQh76W8V3qS6dwlQc8QHbI3Vo5HlN+xFUR0qbAOIooGkdd0aOC
1EpfO9ep/wuApysJoQAN7XKA89FfJX3S3beNFRkA9DmWKe3cfEgpnwyeK9AB4/9R
N3QG17DMX/V5K36gcOjCq2WEszu/4z1Io5wZYT4Kk35I6NusU5yxEdn8z3zUlFqY
2M1Va5Rx3F8FiHUbDzvA/uXOkePXmxMckRxuiAwTMuDyH7QcnRCG8YwbEPJBRz/6
/oVr46XIIX3LtkNniABGNHIcVwXwc7MBgjWBWtvWz+fnWrxAQM3Wf5y+yB1+VMYG
ZXnmIy+K8wPPU7vBQ/UnbCtgzerumOq3pjbUQLVGBdx9V6lp4YHot3tk7qHMfMeD
U2lB+yr5XYfNqodD12u3VCBPjVy6oVdW+8/FIY/WEc5vkkivHliejvaSEBXJWg/d
0AxVd751vWemDZ9ijtfe/K6Cr88M9kQYH45U3kFOlrJ+Ay4Yy/P37kl/gBPOSElX
aWzBkfjDd41sgDk9x3zkZMlKzBnThcjbOw0FoJcDng1LnWFq1MONIsll7JWMYMLC
WsKo+HGL8UHHoey8Raj1VeDDva7ZpU+sruHM2qsjjTU/RxM2uOjWTp6OlhbNJqJs
UAmJLXgfKKXQGhOhiHGHFPcKK4HaKP4OzQxSNzyStIEGFO0yfCBy7MdgDfsNUMUs
qGyOix02t3vaxhkkiKY99arAL0SGP7RnuXEn5MCjf7zve5o+0FdTdn+7hm72iaJ8
92Rrvu+1lp8avwyp9v24fl6TOsR87+/fueaUf/pT5p3QSV9x/ZexqdZeLZJ2IruN
r5BJBz65+Lca8VRxaFwBtofvskgaGSoYDSctflSJA6uCQ1SteupEVYm+xydNQzUR
pzOfmDRavdByEZ58LMcidHvhOQAYpp3n6DK4/LHNzaxo7CW7KEAn+Mz36jEXvTj3
1L3qVwqIPx4vOwCFmvivi9K/fcruFeT5PTmvXDNyhSEfwxAFa2os+2p+Nd+skRaX
o8Of/++9DhOLoCD2Nrw83tjoyD4b5kpDUqMqvJ/D1k+yAW48bMl1llFHX78qSzTF
BRa/qdm8sRad/iCEPhuaBgv/OlzJECHMvLRrzVwje3WL/h9MpQAyMbj5lFN5RRry
DGsghQkqRDHEB6Sg/aOomNx4whWBWWpNOiwCqakLF9KffB+4fckgTvz/nJBYmAUX
JRwU3cPnDQMZZvO6bAy6f7J2iiTFTbzQHas6F4JsrQV+iQijyuduuRInIPU0g4ar
uWJohv3E9xdVVyAiuzxKnip10p6n0kTfmtigQM1IB05EoiuMfdNO/buP/Gx9Jlc3
wEw5za+iz5ZyDxHvEhgeNA0NUZPXIKgTXnywMAtuC/Or8OlA1al4gvw1UqSMoVZh
4VJwCw+MBoKprufwpaDd/C+kLF2Wv9hr2PiFIfh7KwuamEevIHRUj0oULze8dZtB
XEQ88/titvUkE7K9r618aNmey0Euk4ZEIdbwdIn1SEFeqvOyD4yDisLHEbD2h+ml
VAJvVsNNWIFHJ/ZjrfLco0UaNbN/EaxWIy1U+Q28c74URtUB1KlCM9X//2cwkaOS
XH34DeFPsbqkRZqyAIt3FGAE1kS2yb5AxFqxab5Ti1N6SG1WDqclzIOzlH/gqWvX
c+YWfJizNfVxBeD+6BdNNWT2SRiB3K2f/vmg4UwkZgRwU9+k4rSTdjg5PC5FGgYK
r/5IT9KZk+JHwfKvw7OFaV3hWiXowpggJlAh6ZQ09e+Qh2Y3OTjx1sABkpAr+3+G
jfucRSLWf42pTLvoWbFdNJCnuDn98PsRtDfgSJ/j24YpnPrinyjNVBh0GGlbLQ0q
QYiHnuY0ipNEMLCq1GAtQLyvs8gmhecz8qcFwOE5fv3unm9IpmFOsGSS/g9Bmbwq
N7C6xNctJyikSqdfMCzN3SRby0Zkr/C06WHhVqS3nudurivRIXgtoWqkXdtyEF5d
F8JO0y0M7GA+GGR/sVsikcHzI8OauBTxXupCTCmcmvYzJTnIIVhX5GIT+4ESS9Ye
tm4OvcXcI0fNy1Hz6/ulwPBtXEaHVUQaqSolOyDv04FdbIYaOH38mgwvdIoaVDwQ
IwCfC8U1sDFqRdtuVaUcH89is3bJyoc9YDYWgSwzXfjwB9sz2uU6tpTIy5VB7Wbz
IPhs84QTT3rbinOqhwZZFKANYW36jDiqpfdFcPV55y/KbegpLzygF5JUW4bB6WBM
Ipv6A1fwWy5mmGP4HeCH0HN3uRM+IPAgySab3APqm2SKo0HEbmN3lvz1wVzkz7pA
jiLJwq9+1+IT7Zw7n0rSAqOB86sVzxGYQU+rLfdX2cjD02wtWLQGQIbWYrY00ESb
KMRxqSyWiQ/LRq0SE6IhmB0MiTevGtPmfvFlcyxe3fC/0uhxRcScvc743qlu8F33
nhdr12+EVHyEAMBz+QIY1Q1CAPm/gCGJC8ly4pTNpCTetBbcDkjx5+G0KRc6B5BH
JSQWq4odvEirgkbQT8Ii8dSHRCzaxTAGqSa6/pg18SewXi5nvqW1xlfhG70vuaVu
9TYpGLxd+XAlo3bEY/4ihmyuD15g+MrKeuNXKzIBu6ZGHJeVknOYqfaufIl6VINc
MW3YCTXihAZuer+F9j9TSepbTgA6fJSfeGwrEkgrCgr4AMBfsxVBrRLf7NFxax9e
AE9iBxtRvOHoNR6HAZBG+zA9barqCDpMsyDvjFbhJ8Trl6STKjAg54dsC63Mrqp8
IhTyJSkIdIGnBGhlDlMXL2/HqrQhx7QExCZ1wB7Nh+1nSk0MBT9YWVA7ZogtRQvp
rw0IPFTj1kzD4ZWjFey80916dzA02hwqkYwf1lypv1wVaPKNhOJSibK69SmncuYn
dugqlRaEo8pLts5J3KgHRCU2oCYLqHLDxtzE+77pqozLBQtvOfhaB/nPPhLtdFUY
d28mirW8wp4+f2PPLI9ZNkmzRAw9+WUkm8Z4CALJ8J+DEvmpiydrBeY62uKOqD8Q
+TFznJ7bpXEgz2xrW6GNRFNm+fxCjRHF7Mg+260JkRrwNHm9EvA1L/Lyk/4Vaq8P
56k24TXtKN+K55TcKNN86p1yudOk9F7ZFvvXAr/otc+I7AKEQmrOXY6SDpK4XGyj
9OBBN7ML0cQOfQYX8QeqjWWAAgR69aLdPs1lhyyQL3Wv2XDdphvQhEkfBkq5+xC7
2WHMdLWGHFhhqQfvA/NEHJg4xm61EL9ouIJrsLTRpMzpO1G9q50atLsKN3VM+gHR
BoXxx5ln/wsxIXSLed18oySBTgmyORrr+0oSdjdC4nemcDHDyd/tTk3uqeCSbYwz
qz4y2uwSBtBXPe3gxFZvcuCSrF+ueRvgRmdkSS/F0DqLGS1feAd4V9fTR4/s4GEG
nmX4VWJeNOvEP3htO4hGRDJNiFlzWwb4SGlMEQOHs1LCVH2uyMnjQhSSICYdWeX6
2JsSYtAe5tVp8jbC/xcx9+bhB1DMos5XSHF0t5J3kDsqdVtUwBoGFleL78MacvMp
/X6V17hWZLl5pDY9Y35upi6dHRSBXO0yWNX+oBhBaI6poT367XOXnzw5S6czM1gp
A1FLC8/r2DkUVR3dpTNodqrbx45t/BY6e9bBOuy7zGaAxsD8uVWe03PHPCyqqIvw
+EqfzVeOdheSxfMFX0UlYqnIVGwo/mbasVthPHBoPYGnahw2fHsx8Y0v55FTa0yV
HvWTGzavuPoJd5nlJtjE0ysV8G45Lw7K2p/CTCcAWMRjSnMGGIbrzusGYc1vsiXF
FsCsTrwz7kI61sJaFCnmz/RpIotx0TK+R0Eea9lO/Z7zgy9G7gIDZwD9JkQ4GF/N
xQc2I2SK/FzZsMsAoipehG3otGmiLP3ScE0m4ZdVx5hWTrqU2UrOgyBHyQY94rCz
Hpebws9pboJH+M3dv4agppYViplARcZSgxfeoVGjR1wPlYCBKM85204BJeDV1R6r
Rr5s2YBz5HhcCn1SaFmKstGntcEHHv4rGsbZDErNm9bUhoqH3AeaeUWCpnH/AqiE
C+mGFwdpqtxMjIrs9D7lKUbTpvrjNmUrQVoX901kpBAvtWc+vOUfV22muyD3r6E4
mzPvyzLQVEqnF6b1cHQelqhgd/+b0HQD5pgC3Q2fnXnrdgEQF/URofH1BefuVaml
+978+kVNiZMTbjzwWoOsCX4QiIg8UUWkiF39j/ChxxK027f9NRUKTuH6OzhcqlAQ
VJGsMdywn49EZVG2AhnXX+rpYjVjnfMOXFvKmxNifFxYACppDd5etBpn1nHaQGzJ
E8q5lmWb/jBOfhmfh7iCphrMfQJ/YhdtoV6hn6eesp7zSXARZQZN1DxqMY93ox/3
SZ8ah3XWgk0mCejrv74RgfXBg7qwfWzG7Qre3235rXKi8em8EAcHv1IAu7vHLmIj
fdn2o2LXnD3RDoZMiL2QXJEMcsoCdF6OPYLgDGufbwXlJXsaZBPbKTKzId/bb9n5
aOh8ZeVVaV6Xk0aqAdzo37rSklHttJuHRHuhko2fArBjDGBs7YIySERJRLGhQMAW
7uEzQkk9ruKMHe7DbQDJDSHHSsvT1R0Ewvq5BoVteFvy4h+VWayWYCQZmWPbvj5T
JItPpJd6EmkR47gILBjOn2AuW79NV7/6ozX+qmygUpMarMxrGyZVLvQpyCzT1bW7
nYkB+zhGXr73uQfitN/icknzQxSlO83/NQMjhuZ64SFnkkyAVJfJn1D//rQy6moY
gp8H4PZN3Jo7I7A9oQACLRsAISCUEefq6v79n53oHyq2Ip/TdYHLufUjHlOwnacU
mfqpXoCnQSMt+9dL8DvmBg1FmKXsfKIp5naAfKJ6pPLcidjkZHg++15uBl4wiSMX
JLqWKP7C5IeIR/i2Ixoh2SuTJO97aHls3ejH7Ig6qaHpRgxR2AQ2jTUwA0AZmouX
D4WCfyqFNGrAf+ijY69q4VTk23/DXcjklvUYYRfuxj42vKeezOo/2JCvp3Z+qx1o
9n2va5oe+tXRU+H145KvL5XQ0aHqEk5gmBoz6Nmu5/v3jWRtEstZD0pPzI+/zMJR
CZ/XsDuTNtvSHPeJxW3SOFWHREFUjOUnuoN2AuxODb0+/FiR5le2dP3atJhlmk5h
amtIx9n0P/Itlbv1hkfzAKYE3tkqm1o7pW63L/9Pd3nEJJ7zUvk4vpvCpxNeOa7b
e7ygTdGsS4qh+jnVP6/5n83APNMA6Vr4X1HVaeKaKh+rQGpNsRn3+ibp012LW99F
M/BeeFF0ISQsU1eOKavfVx+19TLg/Y46rT0AyPlt43L5uXLi20ojS/wcwOhzHcVa
tmNZtF3hS0eWWAj7ro6LuYBfCCKlg+R0zUuKyYURQSWnlGcma7qXIsZnstzMAKmX
eVNDDxYIRoKx9lxnkAIxuSbu863qBTM3zf4SuXNJUyKKuBmN1pvYwLXi8kNlX8me
Y26AZnsraMGQNe7dOsEC9dH22QDTSmpw7syZR10By3sJbEzrEFRARim4marg0+cc
AvHGZGgCBqbPWcDAGi9dtLk5FBgjB7briUfzyDLaePGqCXsKJMSlMDoTjNb5C5Uy
YHuI5r9BTKSZTc/uB2oetFH0RW6zqSOVp4YR9WyLIpYnVq8VHkI+HPmCnOSVP7jn
hAtlCRB4NPL/QhQLxdHj2nuJQFE/FImTnxaQtIR+bK5Gv1mcMMIysykr1gJFKUbZ
g/nUCqUJpqSWjkxekjL3s/zqO11DX1AkqnKmjGaMrGhcEkjjH9PeHVvim40YZTFe
kP3EOXcutv1ZZ0sTZdZEOK8pYrgu0R3huiRvJlXEcFxZWCsjdh2XfFiv4sZTQU+/
zrr3Zg6gx6Nsv8Lo/Ce5zh/4caYK0F7VR6aCLwRW8gocuUpf/33boz+s4pvilLwe
aReLx8mTtCD15pcxjJLSkIA5fghfF13rwXr2WsduDEqOmZKhWfmwGaT2lZxagLII
wvn01EhCRQPGinXO/wAvFpQWqJnCE2jMLtUcG9SwBmuLKIhzKoyGhc8VW/lcSK/t
vUfggPo16zueUdwWCnAu4SxY+PKtH1Y0e3rZ/y7z9U+bAbFT9LsyNKNeqHGThVVE
NmpxKG19ffVlc4+t+CtqZeO7uh+UkWmVcsez1foxvHapeyN1cmUh48hX8fFY2NEd
lkUTxclLOt1y2x9x6XTSHcNuCxayOIRVhgL7u85ScHExDrlg1TzwuEiymuQ12MDd
KX+rG30EHIcEMjFu49zo8ZvrPDiUjdFmD3X8qWx8fiv8C7jnvHh5+5lV8ulfSEbK
Cbj4/B4DGO5DPchOU9b4BU6xckjP06mlLqmGgrvLV3H/w7Ybw3EDm5qlapz0GJ2N
5sS+6hzhyjTIMzR0XNPdZ3LszkKuCSkE+HuuSQDIt8+NoFV9yEjFBaH0HmvvR8DJ
h6aYslGA3f1F/bWJDLyUz+fnAfnXZWucBvhxsFrRvqjgu7R20cD4QGIVOAfvDTXe
ThEBB6pXkrz1lca1RMkfXaEjtuGdxepFrXrVPqwdHWyZl+hQa9zpfZADgOGUSpgQ
ZT7gcy2prUVMppWQ4Agx8PbCy9iC/zeA8S+xcM1u6hQ6c5ssyl3xmWGTBSHg9rvL
qr4cLsjza+4s1qs3NGy/HzD2CjiwTXynHFiL9gXvWaRAfwN3/eFBtimvLfCnqRUC
tiRZvUIrhuBYEBEFGPrY8FjcWhoT4UDiFADvHbZY8C5tuYzve0rIhFssefjMDatA
6m1cUj9VFL1aPaos779w2jipSy+5KKRLxOh4o0VAyrHKcelVfrwWprqKfUFP+usW
WSVJr5cjzg2b9V4cvjPxE7FavdSnZN+TIakKDiqatSZFuQ8YgwWpBUdgy0css0rr
U1iqtoH+zP9hJ+lLPeNuGYaAU7boqwSA5bfP9d4gzvToh1xaWVyvdjrVf4xrbwaH
VtZr/iJAzVgcOrhBnTtZjn3Mw18OwOu7H5+t9e4h9KMTKhOkpkPSfy582DYsPpLG
Y5DakdQUf3nEkSW1oL7VMAv+SEGwDbVsx9xCzHEeRqxadF15N41ymb54x81fcY/u
PxSoiMjGWYmSdg5g8uAR8SRzerfuuxvjx69n2DyuuCAclZVPYBKXdvICDNGadLGH
TOpvxE+6xpPpzMhqBxJnSVqZZmN/flzHiR8iw2daP+UycRxYv/Z483p7B+nAu829
zJxowa0qrEsLs3k4/x/qvKFK6kgQ+q02NmRvWa+Od8P5MiBSHMisKWhbv39Sr9fs
j+UZqeaLBgMDd7VDr0EXy8m2snkhJ7nqf8U1yjUKPsVEYWVv0TYfTvGHWSQ7T3Y8
QNwUNd1eMF7ZFJ/RGhuAMnPCFDK5jin/NxzqtJM68RJIKijBIYYlU3RPClXou87k
qJez3ZVANZXM9MQjdxzUc/qugXRA+9Mvku0qlYWvqyQseeh2tCLGxxOc/PnkO3II
KipUPuI/hlLDvh44Vil1KHNsNkhTqfxUbgM4te02HOqwHffiI1SJfYLoRIUAx4fX
KuReZwlLkrxq+1SYUtjhkKBrNNU0uZ6c+GkMomTPqfuR+LUsKws0HSC6JWZYVNQg
pXmW9IosmXBa32iJm+S6OQsA32vNzWASW2pAgRw4L4oQwpFWHsx0mT/sghGtnxC0
RU9kirrxeuJhpb7Eb3nVMXEz877w8N94L3U/1EnYJyK9wqAib1CVWBbRJKAJnsfn
OacDkzFWbpU4xeGE3RlRhBuemK0XQYAPeoEYW3KW/6G741eQ+t2DrgX6TctCpNRg
8BQOQ0b47Q7LSBaevMsRCcsCR8NCub9ZEX2ix9ch6XG3PyvHQQiUE+MIOkyWjRvj
jdGI7ieVYcPlf7+v9fbRGg7XGiwtcDjZdr+9/kIRmwB87LeXLQQVrJrbKlV/tyrp
Z7by25cd6dfhpc1n4c+7cUoijqtTEYzVlPYAUR49jkFGokTeEULu2rmX7sYE22wT
4pwD5HY+O/eTsk+TB9fKtTyMznpvStZFvktS5K1IFVNx8XTR3r17EpvxwZQKYhQl
RoJcXLenO1gDm0d4UrRZPoPlXQPLMFvql6EbypXKGFUV69BzMEqn/OGXSJpAnAn0
JppwGL18rOtUALKDhxOZ117BgRgCQub+k18aOId3pMfMpnYb0mHWsoPVfXWOsdpg
PelqQ4FoGrqAqDPhOtWqT+6ofqiN/yYwu9l90Wc5XAQqPwn7yynTvRPHONXiZ0VQ
AuMn+hU15pJ0cSDNU7ukZypJvwO3g3x+52wEsbcw5ZX5Nn7IvD2qPrXlkzqD5+bX
3nK4lYsO27aRO22ol9r9nkaZ014+HNhWu1XAYbi8rMMor1U62Cx6sQJEl55E1Ujo
KyjexSGNbj3eh5T2CIZ9apL6e9flD4blULYtzLkh6ihFy0xt4m93EGPEdtoM56bk
LQqQQ0PBtXTucP57iWKk7EngI2+jqOh+/whMT95kweK2VFpABayNspNidviYZfFb
gb2jTOYMpppzlWNrVimE/6+eWNu23hilq45HCBGGnuSXZ6pQZ+rujTSxH8N46R5h
cnY+v5J8Mc/IIV+dkcFB85mEkaIuVxVgaXTKDn9iLTm4DLGZZPERHay64O02TxOj
0ZsB6ejz6GTQD7HjdyL8AXE5uRyzWgpzyHFa/y0A7F2wEXakqDxULRnItq5jDFgo
b7l83yM5DZS4oyL74wBuwQZsaHhaGKeGCyyOF/djcicpE3lp2LjoOzyTXJ4fHnsw
7pT9/3exG8OQXqoLkmIisPnSmjEHKoJeq4Qzry5pZ8sTHEZNPf7yoBbbtDJ0XIuO
jE4MBIa6IKUMDBTNkiLHdRwLqHkx+futhH0ETsLAP2xE9XmYLIZges4BqXBQYoN0
Oq1iEManHCqA8Ln/afBEweODYiGGZkYKvLvghibY8cSrmtzXVFR+hlE/4X4uFwxz
AhXQTCw8Y8zEZYi2KRNemsnRacdWshUoNsH/orsbl+DQ1aB9FRjC7bGTws+AOgc6
Zc6jsC2kMpxvKKSPiZF+pmf0kpDZK1w9Ytlayv8cwYPoAqVns/EJYyB31QMh6Ri6
5DJcJcDjGWcV8Ht3nR9OWeFRPgUCId6Qq7m4xkeWzeI9AkGJR86RZLevdUaiV2oc
NLJ02uc2uGOQ4Wn5pfEItPe8U7mAf6W9XyEo7wvmy7Pi2TrH7iqWvQczoahtAm7v
SwWUlAYl1/kMOspoV76WJR0ZNcIW3b2Hotf0e1PqijZIE1lIA0oSgZWnnEGFBJfW
mTAPz0ZDfLOx6zc1HFLWfAOMc+FG6Li3iy5DRXIMSbM3Dg2eeHBVRgzjOWKkaB4K
vuLDVpwsemg7AXPbHnwNkXQcMfd/OMtC8AYkp7WuxhrXSSgoocDGkUiGfylY/Roq
a41MYuq7x9Fc30DP+s/ysKcN0ORzTgrz5AzpXCiugeQwHKBTky8TPVMc9hdAZ1Et
C9QjahRtGMeJmUZ6us9B3vrzxAh7ejxutfMcsDqebh5CiJvrycL6RKx1e0EKOotA
SUxmWd+TOGuyWm0tgMWryHNJOvzLVZWAJ9MWtvdpk2OKGw5ad4YOEK6UYLzb0aS+
1AB6agG7O0xL14CZG0yfnQDtWMSm6P9ZkTo1AWPYcvqKtGaeHqqCU9adEhc9FnJX
zK7wcJoAPfucjHPQ/XuZttR9/6EYKgW2T+eDkQro14vR6MBwM3/BKf+7h4yrKHTY
ENZo3EUUxg4lJKC09RKwsQmrsAbu0UEeXYP033FCt99eBgQqAoZNdwiS4sRLX5+s
BbRiQg1Lw/iStLWsV8KAZDl7594Sjg8ViOc2FQ4N7hktis1+6ov43GtAQ1GCgPSy
rNxsFHG0Jn3YCcGEwwFcm/numi/w9BeQ/SnkTG0/t9yxlWsfrQ8tg8LPzoI4ZwZP
WQgTCisSuGddlB6mcAehIXYwDGkmPEIkpRk/t+9PNUjLL8WC4hf+0rsc2jDSR/Jp
ufgILHR+BApGR5NJAstEKK7HARqR2lZjq7EZkHLqDxlX2s69yy+biLJKF8TiCdVe
1PSEqm2Vw/UWPwW2ynbWF+YLOFuq6Y6uA/2DooF2c5/YjqwBFIGmJZBRD8grVxu4
gJVAZfckhTmXIOPYSCBTsZ+sofHjVP3h6DMo2I27gXeSXAcV7cc4DP94G3Us9dnA
qPnco+U/DyWn4R1FrCFPr33FqGloC4nLrpbqTmeaN0bPavG2+3RFIRexwsBLgvnG
k/x30m5Ok6jSW8Ql/1aprGRXvPc/mXx2pOVoaJmvNqh/XdXfCfYsayWrM0gEZDDu
kST1DqAvMn0fT++r1TSEUYYjyoHj7Xm33gHAdsZLCQ+tsEqLYT4zjjh/32lly1y8
O/NL/JTdnf1nQoClXcZiviW9i92JJ16Ht/yBX9XvmkvynK6jpN/wJ5vn8CNk+aJd
Y0AIbeAoEUxPeX7xj7bvesWoO87na2zYIhjHubU0ohICpaXGq0H++4lIhgbN0FZx
SWc/2jWxchFkkIEk6PjNwsC0s8AVfnbeoJWSSmMQiWIqv+9BRUFYEX18hW7RQh6w
0y3P9/+iPvWaVNkh9WABgOvSXvaSM7xIJMl2d4/zVtUpD+egFX5fvMDabLObrar0
pKqOZmSw+6ADLRSb9KrOmcBYflg8F/8Rl1dY0lYMTUWYCPwsKA2cXK1vcpp3e3m6
NQ2EpMUUzVK+GgEEuQ1IucjWEDJKEzfwMAzC5LRqOuVpTuVv6T8qPX3nz3tEMmrN
VOppZi+//YcRGF0BarIAPI17vcN4z3N5L5WaGO/TOSe6jYbhwPBzbGTCUATDpCL1
4rTk3SUyaBzA6wGaSHxXyPMak1skGCXt+P+/ZGX0EKu6Wq8eur8Fxm+S8/wUJCjR
bI9yNQV2n51Sw+srFQMyX3NCVyxcFkMJyaEQFu9izHmdkMx4UBwd4RCh5NjTh13U
t/+GV2k0Hkp2DKA+D3YRLGTFfuuaO+k++F/mf87siGsYeq2j9gNAeXC9bLwbjqz1
8HlpIw80gIaoqOZcFjScfHLLxZJHWkXT/wi/aLB39+4C0ju8yThq5Wbxmj5zC2as
YpHVnMsI8sqtjHarOlyGoSd+1Yq2Zn3OMOUy/e7PGN2JHkoy/W2WMnSkEWhNll4m
YYbb8gKL6rAnI3245VCGMI6Ds5cqTNvda+hLaUk30dBFe5lrMylYPD/xoY3jHgvi
kq6O4jIuaSTcfT/fqL4o/odNSC3vemLfO0hP6rwfutcGuhDFLLL0OsLhAL8W5o5v
Fi0VlUV6WLb4EBbxmogKusl52+QJJ1GBHE9bzqwb7f/6w1DtyHnvnMWrc46eqA5V
Shtg69MpZKY1BbgBDZxkksWGXOPyqJnxWVT6DSUWz7xjf23SmkQbxLutxevxmnJe
GjgowRFOCCGhlXZxgqdsTNBA7vSEb9Fh0oQQZj2CtGD0MSMHn/GPkDxhOXDGLWuh
ir+NrbVgWV85Cb/tvhdjEGRdCJbvnA4KLfgzaDFmTeMR+sbjNWD0Y03GlUM7+q8H
60rt1takL+OJ2iwBULDidWwVsbnoO97wSy2CLkqGIfLth9c8D3FHqT68lIzlQ3Hk
zcMOUtMsCS+DPYjSc/s/B3AdkegHOTGKoYtHxiyZ/ItwcZ9uFjVH2zLNh/hLZckP
yKUrvhus9vC6Ij7LboROlH3IT1mkrKEpa3mKsnBWsbCc/ZR9FXio54+GF+0ta0Sf
/rSWwddXqOvFtzKi4hIb1ZLnOdfhuOsYkSqtGZUzyC0hwYvdrtAnHxtX4YLDOwaJ
B0PQQ3upVLJKNPDkKJQptamUkvdYmdtB+kU4G6WXA6jQkzFdd7XJg42osaAr965x
vjsAXNzF6HVWJSIidfSPV1grG3jM54jReCeDl4+P++/jxt4nsCth9MyWoyUdja52
IH+DO5uofHT5ItaIzx/6MCDN2wqNbKgCqiu5KM26A1lzYzaxIbFlA6mc4YH8QvCP
d1uF6SVcvBw2uhhkSX4aQR6DxZKCz9BqCSvO/o40ArBsfDRNS38ISxIgia7eVrYP
BZ4j+jomGi1ZrOaPoUBOa8kUSVNm+v4jBkZ44vcQpdkr6Mda+3NrbrWmTHnxevqF
qnCOTQs7+ZtdN2LsSnvZkNpjJSOmbE32AckWDdUZ/hLDiSyY/NvPh0RkXHYwbBEh
mNlqniL/JO+BG8nb42XDC7WtrP7qJiIvarKJfFydmyq9upYL4aXgykwWEJjGDpzy
kGxP6j/vSlu7jyEcXx2JSBAmcrrk5+XQx/Z9E1Di732oeO/9Sr7REVRUizhIffP/
gxZgFHucA51J6qrZKXlOjroTP4nXWAVZ0y+9htiQNzIekiuXJiu07xdhTsIy0Z/v
Octkbu9rfK5ne0C+rcoHLN7CWEccDQELQgBc9d9HZybvqmS09vUpVQhVd893lMaD
Wa0SY5MDUbpxF6RzLVec6Un1C1goq37mDwxljCnh6vs/qGCl6WEYYZpmD8IWErqY
c5lr8BheHMCd3NCsDp+UahCl2xojA1z0HD71MqozBFNsinFkbexv+TgOqrh8V4PV
CxfKsujeITwgtdve76KqC9T25D7EP+3glOi0W6jpacHyUYXG97mKE3/WjfKFN1xB
M7G+8/3ReHMis3/HrOTSqqpHZFuTwCitBn914mh4PQFdZb0fmU8Fe6mm8ZBoZnA6
pJ2FpUlYBKAmP/bRo5L/CDDfAuGDiKo1qbxluxjY96gDnFHnaZmTHZqgkk72yIkJ
wZSIBAH+Xflmn0iTiIsoNKBWVYofk/gfLh/Gd4yCdQ9BU/uTg8uJARhEPjAgIZJG
sKnbL10i0GIsraoZGsYGeHfJd6BQ5utDbciWDvz5sJK3Rb7yNLg8RLJM1/hWnxCZ
W3cmdq4tylN33hnCgayQlQFIeFB899hlaRZDrVk53xzyXTFCkB3anqelFTHxsyeC
a5lqa86Ge38mSZjhPg28Mgwoosv+q6xeQv6rZPErmEVipMUG+ir9XxIjLYv6rO2S
lpXk5YxfWQ2Dj5ETwUyUKRDAQvS1JX9X72JIWj8NBYe30sOR2xFXZUea+90wLGJX
rksy794fH56zPh/ZaEkTvVBHsUw4RG1YmaGmjCgKbeNpewjKI3juZKZELq3iHpyx
i8C8zqYHHz9wk5Hgdr91ZyJoAKEQAs5j0KEH/QevVJVlnWd+Ynos3qxkhMSK99b5
DgZOTeOGPQepaBXSmEBAlmAbGFpdNH2geBu07KpDBunoan21466Psr6kvjRgyOdU
+6RLdSQ1vfQDhuq1cUTrLFvlwoxMjKtybPIfLDO+/ODV3z3dZ/tU11VGBWekSw+X
UqtDug72O/36m0g2jnFbTWOdDxCnYaXqRsHozNIWyZ/bjrCju2p773GGPocaq4GE
msqSYbQcxQYxPe4D+b1ebMzDolNhfDMTZvd0J48SKTiSXwZT03dpKqIxOX0QVgdx
zqqOfFmDt+qIYOq/VcgrcNnSSNeiLI/rZPr/NxgxaBLLYw2lfmXaJHzsyQponLGf
h2r81tCPlvDLeqdX4PXYfmTmM73ZsFTOyMIudtCMuwv8vkWvD+8QN5ZDpz0ewYkq
e3B0pdFDjI0oBoMB4y1MDMk9MTxgXH2FHU36yJerb7UO3gmk38sPrEc5SI291gPx
P+g9liWrbCbULR/iZA4nlbctVKk2SsYCE5cONdNBa2VpZKop9KxMQ7E+3aFg07ka
aTWIQxzMISlt8p8lvJFjBPdtFULay0FqwRXv6OolGWS+n+IyDPS17QYTFMHjqVXY
zLXNgP+zDxrhceeco8KPBJgdbLapGVztz+72fG+d/tYVdPujojd1U2VdOXWPvxkk
CVXbF6bsdmSATBaBIaNNDbG7NzoD7oz+yOmmDN8Os5+7HQ0s+mBsLLRJ1QLYcu2s
wtdN5/06sktHnUD+vJ+Oldx/XcLbxaHnEkpJ1ygDcAA7LKd0Afpt0r20QDqereZX
UWb87WCITYdL7pCYoc50biMP3zXXSX4o5p/Wjl+xZ2aL2pprjEBAKG0pBSJp9du4
fHH5llmPs4WzwYAiMRz9e+I8TT25CNurlYgawLlxrBaNbOjD8eFhcBmnTCaTMFWV
ZMe16AGeZhztU9UJx08bOqBjiyp/X8y/SOVGYNBiYi2WS2SLWGXdFxQIrULrDEFh
E70JtfOu0gxi30W8ezt+N8fBhLWVOBI+UpYZYd0OfuRB15DO2FLcInrf5jpOcmpH
eIt8knJAeTsMSoIHkljSxLSOYt7iuL56hCf5O6fM3KlwKFLGh3pXm02NqH6w080n
P7GOQ2AN4aLESzAOw3N6iiuLq5872SMKgUW2g96dIYr5QiYhMvA+Rhf0JB9VaDLU
jsURrjn/RuY2/hnvO67D49K8T8MghAc5RUk2lDSlc6PvileGrYSvpNIrr7/TQMnE
9xIrYAIwa3I/OIPXgD8cPLtmV+7ud7upBH0EcvYGHS/nBCUXRWW1CbN2etrESUUV
jnfSDgiOtD2XwW805JVb+HdAN41WAeO3jqTP6/IPMemcCG4cHDv5QdGZX1IekOac
HjKd0QZf4LbYY7xaxDtx2s4iE1eFWAdEL3+5oBZtjLirXtLqaFicoNZOoEVBfHf6
yOIPxdBY49IPVFhR+YvoLhnMjTwB8t/bySr0qqlPnb3Xe8RxEoKphByf6SCvmO2V
pTPNxZdYYUDQl7x2h73hRLuxS43fUR+WefemhVAHUxR8dyEctmEUFQTacaFvQ4HU
ph0Iufs4C0XfyIpDM9K0d2tUN8dW60S5pbQ05qYXTcRwjLVnlYvRg83VesLvEby0
jCxgYiIGTYdImYjyq55WVc73a46qTB869qEAL59NPtTOFxxM9KwRuYyQ/GRcsXY8
F18Aj7TwM/C/VbTyCq40UmdtPX15e2QWDu7D7W+QHi4baKnqE5um7oUu+VZkuYih
LkdYr1Bu0N47sQO40CeHZZRkR+VoN2AIRoU0wYLkXZcajGZDzSZB6YzrsIi5eVCM
tN0BjRN0OCOfrscYJL4u4RWz3rq6jDrkWFb6Dh+EVQJmjPi1thBM3eKs8GkuNnM1
lm5xOnZJ5YBb6pjg8hz4lln+tY+UXGL0CilZBzRVPOPa7luNs4jISsSKNExOnP/i
2uC4n6RiJhmVqIFoCCoxBXTpoIIRsGqRdBZEK37pwLdozo8/3Fld1iBAmvD9/BUZ
7gtv3oKQehH79cNb0FYzN3kqZVO0EZpMjN5IVl9QxCpJA7EA8aTQOrZ/ZQWf1KNe
V62k095U6UkvUd/w2MLGY1F00jSpTGx3tfTXzQC749ShrzyhBOguGSm565mVM3Ne
z2vg6pX0WkIZDI/RysZIZn2IBf9wh1ELaeuRPCsxluvgZY5gQZ3zUxflV+jT2H1m
86PdXVIniguFYg1CpTgC+t/Is2M//0ltTLKEn1PUtwmFfvsLaLgQoDIJmODy3cZh
4W4ZfDLTjhlo6xDrwUVPnt+cCSarHBtMoa7fgGhSjg9MUx0t8ugzQKmHMaJ07k4Z
a+VqfbpzZJwzG4+iWmQVLX4CdPwV4wicffiKF7ktfVAM2WKQSacnACW4Qaz2DDAZ
qSHfRLIO1BRClOXWmfPVUcugiQRqOZY85A3PFffglJ1y+aEqsGnDZZ4Te5Et2PZh
mKlbIjvkSEDt/lmD7sDev4TfOOqE8I+Y55pYzJk0V7zO0Oonp6Pj1XucTeD53g2s
+gdU92cte+pOCV23JXvDWmQeck6nU/uA1evS1R6OJ6AydoGYsWCAoGOmIeblZ8Rl
gg96W0poQUx3a9yBYZnyeXk2jHXR5mXXZHRKaPrmmAJjElUpElYtRSrkj0dVCEVT
tuGbtikzleaRIsHJSM+I0IfJqONKqkK6NIofVUcUhW9eLWNKXQwqCwRwUOgeJXYY
obw+KuuMq208N3AJtQgqq17UsRWCleOJd2r/TzjGK8xz4bKvY+ANVZ8MxRi4nlxc
nj7fkW5awDgVkLj1v41T8FHj/+VqsEKeBuMk0lZ31RQaGMCxctVJ8tX9qDM4NJFx
j9J5Fx9EKf2D/hW4YVHiYXyrwWSvvmWNgRtnq/YVTpalqsSeR40tqb3RrFKFp19l
2p2q8gHDyFw/Q8yLa4ALOklsScv7BRihF4hqHroZeC9pydx+lHlPQuJpdZKf191W
JlgNQUNYNzB88QvXSq69PyBor/WwI7DNsd8ZnZ/8my4TncrIbo/Xuxa/9hCCrHgM
4GjVXJFePwYaFp8brPL9wKYUpnrjYULWtYEx3eI+/2NedH4+gdQdUSm+hXj13eUU
/zY1fHEswNCNwyuNcvloXwX0CUEDpmP8doKBHc5H9n+a14PMiK0hEMM/RjjcM8DK
ZJYyxgfYcIOip6PYX4i+zhYlZBOhmdg5qPBfPvHf128vuqwoUF9P8QacwuXWoAuh
9G6yiD7vgcmJY8Z4XKaN+HlzZfiIs7Azr3rqb5od/BGxDQuXfDqQCF8NSy7uNvgJ
OeKsDPxcho6atzfis8ggwTlYQ+Bz3XvFXk9m8RrIE2YXl5rETvIFfW3X3VAS3TXG
yboEEQtj6Ea4GOtUbtfN7AqbS74vqjosE1dtnDv9b3BxnAw8R8NQkK9Cm3rux9kb
BFAqJ2h05I6efQrLTNOufrxoOjHlu3GwRSn2bzyXmZDrMCtV0yNQSsyQPn3NCTHP
/WvxvJtfA94LMR7pPsjB61VwVzp+jAocu9GG3+ZJJ+/yvXwSLoowX2nfkTekM4Pb
m2d6X958nS8OlhckRHG334AoTHRTsLnDa0jQr+v3oOMXP6Mwn7Ngj173SBatVhba
ozpvQcC/7C01j+aV/+nnfME88Yj+7vgX+dtrq9Vknb6GPknqA7lIyL+VDNfA2bct
BwI4whyXC5o6No3mn4H1JMrz+8+POqPEYXff0r+zXBr34px3JkzaXOXseWo2AkJj
PdbGjqtXTiSVtoGESQ8t15Rcxs4+481MemB81VYbGC/fgCLNTZfpP4VBkFowwHeE
OOqtk16qpzW3+98oRclIm3groIp7khukS4RnQc/flR8WEI0AMKETi+hMA40R4Lv1
+0bMoG/+rIN9rDFHn6LQkzlmxooRSC/rdyBd6Bc6G53THbaLQFDolr/WscFzZVqr
uD5McZqtTsl63wVV7FT9iKcPZnDvGvFfgAz8cHgEuvz3260gvrqa7VIcx1HMiKLq
Do/JjfHbmLqsdg3WhaHRNokPSwlUoaN63kP5mJ2VYPUQ7qHUSbChkurdHF8RNinW
PTJQXpsjCNwvUOJVh1jEIUz0czJIEgpAFuEQv7Ub6LJlSCEnEM2CtCatO9WhWfm0
REoVCljDUkU3b/uRuiP0/yhTo0mlobLDE4TZDLNIk6bb5/lHzu/NdOZvMOaSFKFG
V+AVTp+iKfbwY7Kfk0mG3ux7LSAAncBR8iqmx1Lxud6kHNSmbwEf4SSzgUygmQJ0
2n1atW8sXLVuKYNt51LAFsv/KxP6Wqc+71PaM4xBI4TP3Y4/6PcepNcjGuySMYs8
+qFibYjbjsXUlq0LXj3Iohh9OI2ZeQO5fN+GN4Cd+9Wytr9/Vp6h5X/A3jCYIkbK
+7xJayOMKaLAWMr47fxRy2nnkwx7fYrdlDwt+w3AlvxXPMuqhweAmRuS36dLkaLV
QdeTeFFlKw6Pp66aXvw9nsJyhiYySz7hReYqW6JAd+AEEg8I3rmcJBwrA2hQQ8gB
jpbT2g75pBx4wgAHlx6jAzDvauT1CaPBs/AMlfTr1sDn/6Qc4V0KH1bEJccJs0k2
XVyY4qcRBiK4Uy/umnatIAZqBrGdzuvm2saUn03kEIojefRXF4xXmkMLM76MO/Fb
QbTbvJy1f9LAFR8IUPBAjZH30AtEK2SzzNAXgzMBIDSScKc1+VkvIvDuy4m96eYy
5AJacjuxUCjuXEw0qzNqzShFA2VctStmcVP+riLnCj5Bjj8iT6lPfBgWcGg189I0
ClzG34pNasBgldeCIQXyux31UuG0rzwzGcJggtyNrTAtU4fzWjKFsewjK7VDT8CN
gWxEx/NiIW0Yuyb/9GAYIuqENGU+0Yr2bLUzn1v6CqpED19+uDyXoaUz0nZh1wbP
42Im/oQr5343zbLA5tRiaJ20zW7kuNOjKfZqM94XZjr9jjLMEdVEBLZH+dVgNVer
+cGeX4gWYooo9M9kkhjj9yDwVhDMiccpY4e8ap/FF2kxh8citabQkW4189EObyCB
xhadxYSUHK0ypZOowamW7XtnZpN3dZ+xT8TkTAlQxdDW7P3hH1ssmxvx6SzU94dg
M9zkGIuZoi1BQGq8//ib6gLN1XAFtIvdVe5d/tXLi81AiaRMfulq/xcRAvUb61TG
DWKseq3kxEuFaZ6C7FXdWON5ns6IcEgb2J2F5qlWXz4y8Hq67HpVdbUdVD5Gyz+k
Ajecr/aVlsiXGdC7dHLsdjdxaeoV0eb2NLJW10UrAcw7PxNuBGunFKRBzWO8Kxzh
9VcL0OMQBA5K3T7Z6N0nnH8WLqOSAnX5KUU/BXzsqAU8rcURnoPl7Irnlo+XTmKW
I/APF5UFe4Q9i0a2ZICEvZ1mopFkRD4qDnmZDey3wDx2HjmAlGGdTNvwNjh+k1OO
05cBGfNRajhNNAPcpHUVqt8Fb8HPkSkZ89QVtSW3uvhX4eCT1zdQ5uecRxbiw88Y
hGn+Kq675BF0BEhZqbfz9uMs5XcYIT31VzxP9LYS0JIZ85OfQoM4eySX2MbS4lP/
fjKh+p99OvNB5s4/OQM8uMwLp2BtPhGAvleyE8KuXvjwn3/l0dycDBs+c4O8+WM/
6u/5ueez43KRqlzL/+/vlNfXj8eYc/PE4B70YsqwyMY3KpOfITefFMlM2pRFBVFG
jnG2w4TKXxnIIcsdxm0M000SYunwcLeXQyBng0stWlf063uNo4z/AnTSzlND6Bit
y5hErbFtqCh+kxeFG30/o8NFPKPCL921O8ufKmProd/HqdqFu2WMCkzh028om1AR
VXpgjRdWcfb+q0TSqz/3vFX+UyAAK9skmZrBTQyUN3FjWJ39cp6O1MoJejfrPjDj
a4BxvtxbMKg2g/PvAleUn8m72Km1seX2tO6z1/fKxrCk90GfWPDVPDbB+D8kZDmG
kgQv2Zs1kSqmDFpGbh8r8/sBIgBnqauEYBBFO6ZHHMznlxmHxeKcloSKsZfYsbuO
XzymPFgzkCeIJbunxnQTHDlnLAm1SsMCSIWcWDAhrvUFO+L14abcnZk0zehFfUSE
Rs/iPCDbmykoafp7XGg7V9wAE229JIKr10kqYI9lfYJxIIH1mOxJNnywNm0ycPDB
eC3JqLwy7AzOmkey7mJ8UDTk2jS3lNkJJbP/vxBWfZLzI2UyXFL5U3GVZhvqS/Ll
KngwBCkXkAlJrd0rP1KAOSHAsv6oTVxYVHDxb+TtI+MQZPOXqUeoUEALWcBlY7LM
b9FpwhMLmn8aLqP5J4RY95kq27/UfYvSXS8WehrgX3opwkIT5Q5bEu/KkQX/swcj
diMp0KUFqpUfYI/EIqHvliFZ2VShXPUV+LC23JHuwQDH6S1xXVji9xrX+PmQbAj/
N+hCi6XlHrOn8u1ETsl2RVqTwbqeTK/fxDc+rkBWB/OQ6rSPC9tHHbviTfOUaGCe
phCkWquJTVk7L4l/esEEiQOnd7qBFxHp7jqUhZPFePvLWTJXHwLxMh81oKe+SXc4
h6cIly38w4n/sygt+oQMEI6VAbMcuf514fegsFZQSiQhcipmELZ239bYxtGOkf13
YfRXdMb/uees8ZWsTZbwA78RkYGjga9GBJfXQCvk6637EwA7fSq2EXZ6xK+e3fDM
rKkhUiuU9/2Ut9mVoGgEEMK4uUX+xZTQB2Hhar6DcnzUOa6W3KLDHr9i+LLe9CqP
EWLI6dijU0cyDDi0FgA7sE77d3IJIpmCBiqNU6NlRyoydJRa9nsWYwVgUsEcrbwh
SwXYiT4XOuiIDhs9LPI+rf0n5wEobOfbgjcUukOEttt7hyjoRN+7BQ4O6OiR9zh3
lKsMCFhOGzsC3XKvUZfezvqQY/1/7BkvEqTOqdZWRrbbZrLmDoPbimzGMW9cmKuD
PnMsU/eghrUEeMo85eAIiHmXDpQoPUc9er0GwXRS2IYfpY5eW3RZtMVFrOI3HljG
JCncBLfanZssXf9OrZJ+c2ApbrfRGDQAhFzB3EVdv7gZhiyukruxGT3rs4rDq1xy
EOcuP/AoI3QSQxstQXQat4voCACzmHMsMjBmTt94Eak4xF7vN7r8WKSz9GzGwxfK
tqV+QAY5F2Od/Cpo67vw5Vxg+yKxQzm/leh2l928YdXURa+y1pMndtEN8Ykc93SV
c2AGLCWJxDYGQrEEXKgijIqpjnwuYR6RZjbzQ1aYbhOPj4LemZmgEdxstVIsieHl
ozIW+ixNtIXx6TDDdAJsCLstyosdBaFQgvYRyWtlPjwRxc2zSJ4HoBkx+Px+nVqp
wRCjBf88w1VRznIAXHb0Fiuk/xPK/qqBYZgPeEDvBo31Ye20pm+8j15Hxgqqm7vg
TvpMiOc2XNQg0gPD8w2VaxPPXf29h+h/nIBCBl7TeqEusH2UJ/uvnjclTR6cax7e
uPyQXVOZ1pqdQ/lMUKv0PqFl+lR0zLFA61htaMpwfVY1+D26EDtWhwiciISUzZVm
gO9W6W65Vx7Vp1+MooEKu7MKXmeY9ubZ0TXXJE5vOg61a1836fwVzKASe2IVS8NV
yL1e4tJn/fM9PTDX6zirJXIwNnYTBCMB/nBgR/YOBdTOONT7avHRpFYPsBHgu3VZ
6A6SkCTRE9HnqCmkNyR5vu8W9UZfZSXeLrgJJ7hoN7CK+7DRwdIQX9tyr5nJbnM3
yYfao7xDDLpqWa6GUFVEL8WaeaJpB6+pfiRTZMQMzkb4bUpII8BOvnA8RCZQ47qy
lJ9haH8y7ewWTR37jb47VTPB3gX934rQZKITX/+I1wKK1Vh5Pfa8HKadxalC3IaP
4nPP+QDMca8JcGCuDhLy2+VZz7I4vuidYJ+X3WHJgV8DNmz4Bv+0Ww1Bm2biRFyk
i6UEaf79XJ8IG7mgJm500QxP1MbEOmpaDgZYp1YFb5T2zUGHsEDHtlVNe03jvBaU
Gdc6/iHmn1xrtT7MHCQCPU10+t6i0oXfkzZaP14/qzwS8N+j9Y1a0DjSlBqhjVTU
IxAupaXBoWoa4UHMVnLxjMr7W3wb785fVuZdU7cme+vo3CAPq4SJfCwb4ad4DpwT
NYG9IaWtyiN5t3ypjR7tz1bvS3/XfnkuSjBFkxiaeo7fFToR4HCjBoRhgsehjndH
/X4xP4Q1uHHkhANCD3czxatZUB6n+Z4gA2D7p7PvNqaPCtdRfjKsI9nyMbovt4Lz
Tu6pWuqBuX1U7PnrdZG2rxF0xCvw93JX9CW1pYiLkDlrFZ6W+8zJVHkfpl9gk95v
pMvgMMYI4tprH5VTKH9hBM00vgGzeR5KJoFjmX1U/fB7uEpWHP6/POtZZi1f8Vm7
X3gVPr1TKM0QZnPTfIOeKzXDKFlZhuWmjWBcqa5tkOqPOC5U5M9+04kcJk7V5QvE
3lBJzpTTJe70io18zxYaq8HANQO84wa0o57dwXXx0OkhY8ZE5K9O0IM87Fon61kq
dYJb65kJStzGo58z4kiSICneWsI6MhCvH4PLx2bqtlY3iuNy7G6IQtg3gFhk0YPa
zhEUE3DJSs7hZQbXoiRua2Igj0dCXB6a66A3+rchCsCXNXPKj9usfwiq7hahL2S9
GocMJUuPId6POYjzp26OZrsqnqInZSP/UOVwyMmkEbbO5JJPz7yCbp9XxOI9ZZJj
Xi8KwLM3etbrWQ4+JxbbN/2E/xsDr5ABCZXcifopFrPL+DrpSNN9YKNLNiYmnUlj
luphb5bJ1W2dAmUUxH8xcahczSu2fhtesx8aSLK0VnHQJYJOL3vH6kdtHAmAeoLD
1Rs+RcD6lMQu7i6beJ5IsvpvywetKJiKHFEafAqKNYF53SeIObF/XVjKXvFZdDTU
PIb7SbnYQ4A0E89t402uRZXOUWQICNhMXMB0HFK5OW3MccNOqlvW6imRcw9P6S3e
ZK5viw5fEUq5rqBic9uxzCDlr0HqbhttIcHkyjGOE8ZSBn9uys/vKLb1LOdGLs1g
agDWA6mZzJEss8wjt2HMegFhh7wWqeAIyD3mA0A/MIBRJFtazK6PXhN5wLB8sZSa
eG5g2M51+7tKJrycItetqIR1nWU3A4kysUxzh3D7TR6cCrSpORxiMFfZQztxaXJO
RA4cB4Qvc6n1SRxDnk/OXkO1wncvvg9qGwCZRD+/f0cU3PeyHFgjUFi3JWXkwxfz
IzHu0bSIgl2YFToZSLY4o4xB/uaDk0cbYZ5SYxkxtxgS193S2Hv8K4hyrmZvqQ7H
CUszJkJI/aNswU6NL1qt7RqC9ZjQ61cKN1zZpQY2P56vDD8jt82DN2Nm+ijYX6DE
yueIZKKbtkEhg2rxTi3u9tkpSqiRw0N5oUJFOCq3hjtgXeWzYO0fwg+jsojtfOgs
zci63ccD5dV6Ohbm8RmJ/wzLQqSGOLDvvrTdfOdrS6OwZGSmeaoYtfo30UzR81LA
BTKrCFUVYcwwxJTMZf8+MzsXZIQ9gndaNegzVIIXlqobGOQlAr4/YeAa13XsWDy5
CWANpP7ewO1iynFKqPLXjq3WQBL6BUUWfm+Wa+5ch20EKfHcFjYzSRQdtlg+uX/A
IyD+bENq5jt59OPqkHMt4JNm4U7AgKRmaaqK1phE6YAhHHsFWFX6SiPl/o33WpWE
sz6Tj5cbhKMoo6kfXg/6aoYJzM1JOb3z+MNHNU5e3eWEccTkjPPNhC/V1mkyaoLO
CnN8Zs8ikZkuM95Bdz6zim8oECjfNLtBf9ELkmi4q7cf8cGLCVZavRVVKWDCC9Br
e5kJJhPpD59FxLnehjJMs1fGWo10oAJF0fikH6GJKIVenyBXL+y4oXE0bgxKOOnm
oQoibzjssGOsMEvPh1239CSQ2TMNW//04Aey0Lhgu92zjVf3FqBBTdTpNxdnTkc3
6h3qjEyhVFdXEhiIRIIJLFYiDX47i+9wg1Ck1iT8To7hbrU7etXkpzRRl8I5IVl8
gopCRDQn6St3obZi4xo163uUWcxt3yOUfIQR4z/sLAbCgsSBeVhhJ5EMzjtjlRKy
SR7rqsse3ZkSJ4LPJwEUw3uRCicxgdIdnIeLI5Z0/5iiFCbw0n+n46e8XlVw0kys
2zisTLgqWEwAggL7BoE68BKjQ+3kqyI3BksFdHDCsKjwPq3Ph1ymukdSsEsEajeB
sl3Ed2w7Pwn4VsyJF7tIHC5Fdzi0KjbAifM29VcMOIobiFghOCvmaZo29pOKv+kb
Xc3j0lteQ8/fHSCO8UiSDFNZ4dSv6wDWKt6EXsyczOU/PSoGnVH/dOEAwGkQ+WvH
ODaYNltwsaNqsgor/E//tfEPfHFAyRpvs4F8lq807bgEKBFqm+X7azTxtoy3QX7X
UcHYBn4Of/XOB9fwdLDG+DVxKwHBqGEeOx7VR70CPQ1aWgv0xW49atAwWOYG+av/
ZlB16e+H/fAGTu4gidz474KwXSNlwy8edRr+UHxfY8MSclAibPSxSYsf+U13btV5
EpiFp5M1oCzsQfki/qKa1QLv4NDxHSn48gNntBMnt59oW+JUXkDpkpef3o/6svmy
nUl7lz0dGWmVBNLj7kQ2jPC5E4tRjB/DjiivbYqH0F8CK82KuEDSwSAECvwObrYT
O20JfgzsFJ8V5976LWxSQXL/m4am5Q+Ht07iKmB4s5+THWJOQtnlv3fsLmboCZfI
kDDe3FQy7uoOBf2GD2IudbfyO/U4rB18m1uHWB5d53iC0tYbZcXe8WomcmVOjt0z
ahHp/A63oeij4S0RW68r2VN6OgeVOW07ffHp8xmMRx6CP+YfDIcmUFUyPABDQ5Zl
yLZB4JdR/6XfzESJNtYBX9YSogm3qBARwWvb/TPNnDJhY2doysYzNbu0vO0M+2Z0
C+Ks2UQJIz7LUNBiXqsoEc47pN1BwSN1dxJqOGENrHbYCrOB+a2NSslJ/LBg1WA/
pY/vRxnHM36cjTQETuUtLEdPZTa8QX8JCAJwF+/SWtaNlT0TZstDxuUv6oZwdgdL
DED4hXvRA17Vcu7FrlnU8dpIez9Z2H7GAxR04/E1UB3KHRjkzTYo+5/EOxbe7wxm
LpXxSj7Ye6nOaQFtCsXJd/4ji0JWIbkJZgslFwCG0YgM9n+vToGCy6adxcrDRg9M
sHeCoaNCXqxqVJCjrPr808P4h/54mBjtdMzdLqpE2exOWV/fAMHNCZwhNwrKzc30
QdAW0IKJUVs60SkEs88T7psX6EpnX61fz3R80qdxsoi9ufZL0zdphhghzAakGMjJ
ZketuMHR30rqlSE5YMU4JVcpBX2wJsf6c3Et6XwMXmZwYi+5FyLETccsMCtVofdF
jIHFyBUMR9mXarZeRJSBwyVR6I1JyXHfu05jvnrCRyvt28SQVWqWhH/dxkqGoFN3
pi3IqfwAL8xl8ubQTJAWMe+WwZJaGKFPG9QpIoynIDeco3I4/MsIzaRDZKJXzAgI
Yfz5ePxni6hJdN4HIH/V9QV4L15YmqSAsW8j/ZOs4WRcicGWEkHNRUCyi4zYVU9M
y2hVHE9Ctzc3NWrWqBDoASMzjcAQSP2J7DJfc3O3DIwMIfRd5Z7kGE09VxJwTfHu
rE4ZyNwd6InPcUP5/b0EvDm2OkXxQAeBR4nHK8E6uQ6ct/Blwdy++pnAr3/C3I4d
9UksVkHTVxWaEoXK4AnLeNTogzCvlu4G7aDsGjsFTClEHWEIF1ckIMrh1EuwTvcx
fMc/ElCMRuAJP7GCGblpcnR66PiJ68vpyRwMUyZLNzf4yFaNz2Wn2t8o0RbpFVX1
glcVQ5LqodNCCugWL+chw9tUNndhn0ibcrdu9ZJlfp+9FGdPRXHb5wJI/4/31qI+
coqm7qAW3b5CU0kCmDvldmhl94E/HX4B2WA2UFzLeLC9yLsedCLVcGphieOWQRe4
HCT7O6UZRR9gQ3zJzofOo9HFQVpUl8+dqT6TUAXhv7OrU2rlXVfN0ZXsbBjDjp36
VIeSzyM8we0W92fQwkD9xe6kpmcJ5RxzpRSgL1OEiAEQt4B5DzdI2cf+8xfI2ZbU
8KvmUdOqKa0526Cpd7D5YhnTlCuH5WJXnVtX5gTaU2TO2yMm8CkNbMmPVSKgrCaH
ZWCVVKFPKuAPyt2lHJCqXyEgIYj+chciKSy2A72qPNTDdSJREzFQgoGs6T7llSk/
CD1qO9RkoSbvbU0Gnx9kRaADtarx36nlyuvDy/QI/iFhLoFwOAA3ObfLBK9VLDH3
fBmXyQblF3bnoxoZYXNjOQaDSxm98kCzRfT/Mk7cvKjK/iG/5zevFk2xwBAkVzyD
Om9mqZQ4Dd+n2H6nZM2D8aZaxnRgGmbRkB0ILVrhR8824YWhlc8Mei2UtadtlFNS
esFdQ86PGNNywqkuiMRAWE9tb2MZFEcpgzJuAjAlxoOdj26ySEi/bbx3qliwJh/u
219j5nZmyJ67ycwUWkU760iEZ6Av3QlhNXUVV2TbOM07uf2PRkSDSWBw/qkgBX/Y
GnA/FrurKI7hSHY4UrZDsPHzMJHy2umQUtWrsGXTsCmQdUe1BcGBI3a0WFHHtUeK
pzIbn0rx8d12fQ1Ff+XWyh+lZDGSygy0I8eVz4lNiPQ10Ym3Dr1VeisrJ5CsLmXf
cZCUmIKWj9ufmsgw7o+5WwrjkwINK3dCRrCLSZAUVbrtgUOkIfz/QCrh5dbz6VAe
NbavftWZc5jri+ICLlyp3FWTkH8wmg2KNvsHqjfkp6vx0plKF9z7soiXviCdFJGn
cFNBcXW6MZU1qwmkh0e1kjSvGmMFQho3GKJWApzp/2zRe8sn9u8htXNL9IA7kp1u
nvt1Ec/xpXP1rqlpIwrXMZc9W1vPAC3UGaA3ZtNhOl0aW1i6X2kM628v0zdjHnJI
lAve3HdrCSfGKidrJUz9hU9iG4moMNQG70T0NaBDwi1VqG7FoVjaA5seBRUCGYPx
YGGqyMbArVxAQrunLVnRht36Ov+QB79Mg+1YdsYfbF/M66OtofhsSWzy0hLOZtpV
YhfFfMX6XmsTi5RKBf5yjxSIafNlRGBm0Mq9zAjCWoZZwjZ3eEnd1og9JLH/IVTj
1kKaT5i1pCGovBWJiPFKWIx/HN/ef8HIMtv8fRj+dWeWBsl0ueq1b8Jd8d1wCEdZ
rKzwZo6ftvCntxsbJWzcnmXztwJX4A6T3GoygHtyWJ/0WBTPte4iwIAgz2lbs9CU
gHEtYNePPMRj6UKn+/uSrzIQ5QoM4rjEjUn66YT8TYSI7zb6Hee4uALsWuKYG0OR
bkba39PuyjN54uzZLOE7QV3sLQCO4zYp8y8nNOiduogALnlMzJE0ITdyqwmSdIeu
NyzL+liAhGExfx5m+4SYG96flUi3/R44eJALZxdbUPLZe/JAtYtbwvb5gYRdgKxB
iQ7mJeD2o5Ax1VWtCyZOnSwE6w+/xCx3epYntYq2qBYQ7Z6i9BL2t7pTvGb2kUH6
kc5pkDruB16wDu2XszGusLV6wtJfOz9wUySrzBAMMYCTgeCch5Q/5B4tfRY6UvxK
u2UEY0M/jzUZYRml3T/0hdfDknUvx1ujBYetRTTHFZr0yRRB5LjOjhlhVvQU1+Md
NMmZas9eDu/FPuuw4a+cyERmcJ57Q3gTFCLmXtwzEuUY+OgrErNhUza3rWpsZIuO
ncQxHb84iDcgbHHSWrs6Pdsngro4M0h3wcRRZv+OAXiW3rNeFGridUu71L0bAfTy
Cx49oJfU8WqY+jK8upT9GG/6U81+4ek38zwhFf2ZlsSSi76LsMPVOV3A1ojiHKqv
xYBc/qXdD41Wuocxv2+3rrh6wC4Kk4hQFJ7r6gv2Z2cyB1rSXoL3a7jrRTZY31vv
lRDwSiHSMc9QPq+Ds6YN9vUbhH4jH/l0iacuij115IO0JvEPXmySO29VCdXejbTU
HTSVVO0Vz4GFEAK/oXhHKUc6czt0X89sn2mV72LD2imhzOdmu53z8551kxES9N7c
hoMON5TULvHqX3v+75MFldficRYb+Io3WqrUvDgER2Ygd4loa4k3CLYf3JTeXxCP
+KFRHNYCsgzY3Yq0Nwpw2XOaJm0UO2CtpzuYFcvRH0xMmrT4JA51erF7MXkB02HC
Lyu6QoEk+X7L+6T3LACYYD2Tto1QzgVByjtaMyIdnlIRG0uP+9oGznUIcWzfuem4
oFD8B5mbfp4N+TAKga4npADh7Fnx7uXb8KVxsprcxXyB6AxaKS72asQhOX7n6m+R
iREcWr38VhUXiSwBRR7puYCKjEdSxhOxt4XPp52EIIz+EWPPGQKbysPbV8tLLtFa
dLIGExz4MjPX9Cix70lq+2XG/XGQNQKSKti+kkcEgScRC6ShAxFfN4eIBAjbsD5d
uuPNBoLYCYN5znqcuYPGAqheCxs1aUDD+1irMZHME4QjpDlmUm+jQbHoFcLmzDUr
LMDwcEbn8sfT+1wmwXegPml8Do8JLLDd9mq+zHd71sHg4U5mLhEK4kF+BTVC5jIq
S8ZBu7N+qLbTzWTk5eRSVzrzNH/UvhRSTw1N2YkfpA5UkoywrmtPq1rddV2l9tBZ
lXR8lW6B9RrdQZ/kla9hhFZz6bIIPF/9/5nWE4f3GgHhSwJLBAfN7GBjHEbEmFe5
8k2HSOYecJL3CYLM06nM6mksnaFIQMwqg662hl9UoZ74cPRv653Wdgon+qhd0k9s
LlvZ1DQJloKeMaNdrcJmpx4AY4oRtYAp5cDgAwbRmvhcNumcEF7HVz2UG2ZJOJ7H
S8k7luSrhLFTv6m4p2IvXZkjUXf2fR1t+ubNVZcfOTskIKl/W9FtL7O+JzX18RRq
odqR1dDwiZ+R3z7rBCIBW070BtA7XoS5QdyZX87/LJ/uLOHbH6jjRhSzwDGidpk4
KXTvJPFqpfjB6TAhMci/QwIrk8Fp9inJYMm6iSzv2YvYI4y9kbEiDQOHqVBt0jK1
n+MN//JKQOqrxlMloFUHb1SbZP66p44AjnfJg4o9KoeyyrQw0FFO4rN4mW2U6vNp
R03xH3fQWoAdNA6WvkHD6rsId8AgAX7MLH6SqleK9//xWA737xe08V1xRNjZBerO
EZqDkh8nqGcNi9NPfYXNGOtRboejvhSPSB6gRCwW4khBApKZaTyAamDe6NUxyK6z
+GqzDRxxwX7e9BrNgA2D5F+QFob3YPkmDMUoNjiUOgDwJfkK6nzwBR6ZUa0aAbka
Uy7/vqUDISg+KAUxARLh2RDL//kxHwBO8gaO/doiz569FiNK4z3IE3iISpTwbtq6
rkctnRqr3LJVlHT/4QFSQJHAh47m+Zeh9hpywL9aIkM+GY+4uz4TtKlus1QTYGqC
GEY2O85DwT133ZAH/3rN89r55IYktMuv5vdBQiPmITtoP/ttlYJJcwdNmRgXDaj6
nB/emvmIoCZDwS/xufgQG5jzo3b6EPk+nSz6sw5CNbJLb+8VGK0d4Mse/zN6RpNz
DmokvW72BTINSpCxVkleEO2VHzM5Mq1oVM1O8EWiTDu/kCknCLyZmrmuvbh4SLd3
O12Jz1Qg2f3/O6LhvvW7WNNRENxlqkmZ2p0aVeSk5dTl2xRmyFVrr99iaSOEoqCj
wR+CrQLyvOc659oPgyjAuRkBrV2UOOdYG6HGcxeqr4Ua2GD2SrbCge9BK6E3fb45
4CqHgNE4r9ZRBc8C8G7gt0mLquFjS9ApdITpD3e04WWKy5Skh3cQ0Q4Rk9Akzx6B
TL9ZvtNEfRxioSVB1044pgEJlMM2V/2as4bMpgyWHTd1DaiguqIVyUmDOVmVtjiW
GFETDPsPu7X26gl/jheh83YuclYYS0cTat7NXByH74n/CnEREnOqFFVmglYhif3n
3cdfVfX7/l09SfUBGaPFvarfwVkiwMcPCRarXc9Y1CRtifeK1pYzJ510I7ZU9l7S
Bhf3tlyZBBOh/BKe5YG2w7DOuDVMc6kDcPVdSX1YdK1dStTf2ZKDfz6N8azs1UVT
wbSl1JDnmhii+caerdhw+qWn2hYeW7OkOjxdG7HB8HHSFU2FvlWC1iMWSzJP/Bzc
40dfTnVDjCQIYJFrTbMsOSgEqmnWVYaiMoVpE+kPG+rAvzFSihNiQQWdwc/y4im3
8WljHHjSrH26pbX7Vpyz6BqTocSI4HPIBT2P+zv7USl+JmjyXUDqnQAzljl7tBm6
quS5eZxLTJIkXmBm9m6iexNtRi54Z3thFE50J7cyq9trVI4kScf21ghkaca1azsN
e7asgkFAYnOT70wKHVuNlMYEQIThNAjO5MM23E+gmgWK6fUItSR0Y7rqk0Jep8fh
rbMoHaFgtHsrqeIbwIfQnuqAOfvi3VK9HRL0P3zeoKxxCCx1EOTm9XnNzfBUcUT2
h0UvGMkIVFihfnDihUD3PvFKSsjE++u/3zd3LXPBVYbt59xWxL8gj1qbnBLYY0rl
3aE32TIztNxx20cRylrFmEKP3dz9MaKnKPLjPfjpYaKv+qO5oLl7Szi7iDgfbSfR
QWgK0egADHIFxXKiRctHJCaSWAIC0ELmbvjWdcFv0MqlXgJyIiNJYSzW+aG2Rw9c
Fy2cb2Z6FK5ZyPOh9n+cm8rEAgdd92bsa0U5KegJvxBKh49Tzol7bRsszTbp/RuI
utvVJycgYHCJrVkTPADC/FdYwxMoeOucJf3suSW1apWUEcE1TYZEhfNK3jypDXXz
vQGhwy/CJ1AQiVcB2ui/1q8s+AIHBLSiNxe0Te3WZ7NhLsFosrD+vtkCtsmaxnto
QE6g0iG/hPbpwcNwUfizW+ZF9VgBc1PyIFuCCyHKN6r1SYmG/D2IqXaBON5rrXe/
gLcTEAlvtRUmMxTRYGfR5njQo6H83oa8xS9GCahnNkArSB3SPrmteGdwsrmDtHcW
d6Z723ONvZ9rNJlPD01NYidAiqMRis+eW5gCcK5MRDgacfMdaJLvXNdmjxxUXDdm
T4cacmjpa484XeX72Ikm+ZXB8SRtpMwSxXXRrd7IX5artYQ6C3OvP6uPEG5Cpan7
cYu/sudIDKP+R9VWU+cZuIv42tawvc5j8kC+ZNHO+La7G4chsSxk1gy2PmCBBlfb
Imqmz2CFjSTVSLXrgbYgzX1zbCirNSb14t1MzxA8vcTQwf9G/eBxlQ7fYasrhs5H
UsgrCw9c6sR4ITyeH775vih1VCETsfuY7tQATq6BxenEMC4doib17F/CWZhvPutn
4UyjsQ5rZ9QQwkxkfEpg/zcoeGkx819qM7OJ1bESA2I26igZcug/bjleCU3QAoLC
Wvrtx1RYWhNO26ZS13THO+/ySZTspk8hqBknvJQQNprej5uhBX0SIqNZlmpRxrgL
r3/j8pIS7znTRFB1XZ+kzH/vY2CpLQrFRY1HWgTUzXcw0UJFgKbJv8HAGE0pBG5A
iTBIVlor8ndO27p8DUJwVBuYJ+Maf8/4QJVvaHELjLhbdyhWfca8TdQirpxpvG8n
sYbjV+HQboIFreowzTGM9/9xZGUuz4Fzh8aDQg8QSSOcqJXWEROoGXbf29NWR5ID
c69bs7pKpmNEfyprHCouTu6aRkNX7bbS9ixgJP7CN7hOES94aZAfbOm5+xhffifP
ckmixVjjqN/7ICMO9OVA+8JCzz47q8jNMeESbp1UPr38GGnLceZtc4+2XJpLkoKf
fon/SsSSrM17dlVnwLhqg8iMD3DcrueErcNhGKEXfjWEfY1qJIwX3oqqXW+2ae5O
sNhNKUg7aLCt1l+Sm0WPSXH4C+s+4qxzt2Pk/o8K9mMbrlOr57ERSS1Fp05MjcsR
6AljFESIYUl7c1MlXBCnQwxHJWzMVx9SV0/wUOWet+BE6RQdxcNy3DTHOC1F92xC
Sxncs1YG7oQLeQgqhpd8dpjuQjWaZsJ+3JWhoUnKesJihaKuwoONkyVP4J8SQmc8
hrTtuK+1P6RQm+4NLNwjinRo2v9YdyUXpxKRn+/jOP/4gOuR0fBtW5Sv8/+jQ9R4
JOJ1YGylF1JxqclR6uutvC7K0LZDe2Y/hzlxaUC8yzPTwq67EpIOIOXITiDTfr4z
/mmN/+Zlm3rv1z/yFY6VLGtN1BwbgGKWpzI3AFuQjJJy8GIEY2u0yEagrlAn+4rQ
bAp4a1AFJdbcUoUZDSZSLamctyuSQnTop/ssfpJPNky3kx5hCO8Gp81btUsQWwYm
yZ67l3f7ICEi+0RQMFbqnJWAEXEVSDAsmZTtBDqXfilg1G4MxgngwlvupNsLomyz
yb9hj6assNe646O+OhMBV0pLSZqW0dW+zyE8Wm7+PsFlUfOakaY5tH2Y7UwhSR+8
eREshBeXrm90beD1l5yRel4Y7cfSNkigB5zSEU1KhbePcnAWZ3q1/pGuctT61He2
RkrZa2pgGMmKmneD+k5o4rEn5bnX9WJWA86PMdCfXFcFbrL0sXPbfyyo61BoE6UP
U/Uqk+wlkoU/OC/dKAQ0QLrUIlbkWIsnQg5x8LsBvl8jWhXaT3gu2eRTizQsgVX7
RNLKMetCE1Ytv03lzHpDtGUH41P5kRE2NeghakatKjbFZb1XpR+KFvpmCMHjExcg
w5g+55+evNQp60ngo+JOdV0I1YS8OhxdBAbPqJg+XckeySXSspNh2YW24fh0etfN
35kXABLEWeMHH9Sj+jo1Q3usO4DjkT8Tyxy61lwy1kjLadSIvIikTRMsa+kK0dey
RTFFjYx6xfK3UtN1C+0IPQeYXIYuzxjdXHF8LXZyRhZXm+2bJHtxf0k2m5JTDQhk
YBteno7W5KUjTYYiWg2hHqJOmLku4nyDJlztdCM0SgrKzavRPMaCe5L/ra04yHrE
acLm41t9EynzXF9/fM0e2/R1i+GknI77lvZynijl4Qt8KNdeOQrKSTiJH8cafgCS
sZ6+4YNBPjmdkoacNrYjT7SaLj/vL3aNXQ00qv0Vx/CcQlvuEzmM/qBS+LasqQXX
gdGY2jgVn9Fs2hlTE6kqEhAGusDpNzLDmHJ9DUsmi2vpZEm7lzGOZnZ+3LUY1uWD
BIHX2cuzeWJQHJbqQOlOEKOk7/trJQMc2E5li690Ou1EPL0s5QGIbyDGlZ3ZjmxD
2feBVIbTMBRJnkIsg5SolmEV7aXMzvcNzkWKWF98U/x9DMMG/gaXhoRj/gjcFJoU
iwWj6YCXnYgosfXoF7DBYfmNgr1QfeAJqi2FseWtMNopnqKNGx9EysmiUkggPqV/
LYo8/Y/jvbzguJPdFK+Yyh2UfuEve3653IAcstKD14LopvIn1IXlACggyx85gfke
wFFFidVyyN3ocGJg4g4gEah8JEd7Guv6wUpwwn0XdvfM0tWk+3YlAHIn8pkS3Kf+
NWHhQWInycI6UAV9RMcWLJYw7pqYS6+gZU4IJc9i/2QA5Faer9SOn5KKwSJGHXYv
AYM14QjvKIYLqCGAyDEOoKvRnGJmdzIHW8lgQfLBdI2rLtbb2Rq8P7RTLJ+rLfku
2oKmiEosNYEZ6Y11fE9BxzX6Hfl1TGACLT2fiMKSCiFkrDB+E+chDVHiQfhhtVOn
xdLqEXOey/KdC+mouNWCDXdn5yhvoo9J6SZdTpp+oTybdC7ndzD3YiwvdukEGty+
I1+oHu2gL/gG2Y+xanV7OlpbeqcHFt4hio990Jrkb4B3SjVp/fNXYIrZ7WZxg3ih
9rBJOZyVOb13lHBtuUwgWYkJTBNcoDWPIdWzOYqZJjVO6tskIeklfCBnjhCxA90L
ZNhTGAf2JHNe64YWQCHDaY7iDdJH+i6AIu/bs+hB02bBykBlIs9YnDutgj8q6DXP
9m0fd39byHfdSGVb3ZDt6fJ0b7B5eYZKCi2EAk1pk8dX1/hrnkafTzwCrt/BtvMK
xpfo6pUanKtkJ+uBvtU7J9+reqtju+TPSRDaZhVD/ARRiXjTrKSe4LCB86hEWyNi
yqfo3T/AUsxYQn4s5VkDGCFUkCltUi2mLdBSUPmHK7hDlG83SvVAesKeIij80Q+P
ACo/T7R2L1QfwPsdj3bpBeA9m7/ZKZ9+7L6KszHIULK+hHiVn7v9wvWiFoXHJmKN
Z9vc/UCNJZMyJMx0sw4pF32HP2LfWn28hdpi8tZLBhbJfB91usumUhVB2OEx8kJO
XAJPFX/KGR3MWFf9Acxy40ZgHqBn1Emf0/eq4nWNRvR9k/TK8zhzgLrm7y6e+D43
jOuuNoVwg4fLcQ8i0sfQD2zXxE6onWaSY0HuGvNS94ytlVh5roFkP9BniVkLgh8N
3p7oG7YvTdihdSWppfxfG83dXb/LyFK571W4Um53Y/uIWSkOheo6egkFmiFvmkeu
OPOq2E4slvhaxI+D35khRb/ZylFrYGiiwOo7BkHDfQ2oah2ccGcEPhGQttNs23yO
jJpW4QaI2u4Wjw9tUWU3FVcb1z3rmMi/658bIvxjbsjbFBEafouwf+I4alQlXLJc
a5vJUHPwyFUCOcVS3vpYnr6UA4/v7LGmEavkTG2gWBrMC9xQf7g9ib4DGBC0dnok
s/gtO3iK9ae0wFRaY0F4CNywAjEzy5iu3eFllP7tAifLMErYHoK5hG8DsPYQAji9
2uuzMz+YTGrtrcy71sYg/ZP/SbFrwXuMoP8aw04MYHHsJgS0GlxH+3VIusLNHCRa
nNWFZYPL3CcAfCSpZQ+ZYDguzKm05vUTKrqTVBydOq7Dc6aoJaK0pVfBl6moxCUE
uatrClPIKTnMOGuXDr8AewWc/5j1vsrCjolr0SsIt7SRnbabRa51HJ69J/mulYel
UeegDpnND4V0cOKUdvVdf48J8sjbAznqro6etz8vDQjOgPGq+5ZyW6EKGXmi3XkW
LuAxs6Vbpcrfm6IYptnbAvX/cGIcEyCyTKuZ12xxKkNf7tOGWHBPipOb1GfBhtho
Ma5Q4hXPefaI1Xkno/3fnoNzUMjzuN3F3BsVMNwxkcccnPqXMyQ2v4E+zQ3AgNaf
EBLBM6rFAZAVB+90CUl/PuFnm9iGEq/KXO/UglhkLocJviBHZKkw0hbvepSUd55F
W20G8YsvQYFZBscb4HJL72slM1ZWSIVzY4EDoW/7YlFrlAyfYNCwq9jheJxNQExj
gDoUhdzcF8TbSbrEuGCwBzJpKpxWC3jf4yY4bH77Z4bM7FRWRQIJlieSRB72+vpN
CRaDQJykadgOMDWKd7IYDsAc3D2XXlAwANyveGVhn3+/P/2QHax8TD5EoyfI3Xvu
d3O63fvhs1uc3En+4t4sWlVpDcEWGg9VraRki4PzBe+Nl5+HlvjuL3Zm1C8L4/XK
tnWql+FxpMspAwlQf7MJZbTYuaW36CNXRUQL5bi0ZX8vyqcG8SnNaScgc1S3Tlh/
ZpgabCW0+LmTIRVP++MdCBxALczfvWRfNblmbduab9/24dsLMkbV5pDo+4+F2SZS
ITKU72G8os7A3iFsxsSgpe44BPSPm6EI7sbc6EO7TE3Egpw9bLEkgCdcchycxw/V
7nXWBPRrYTs64gG51qLoLxJi59whnWlSoho3OJx5/S/3c+A0KMQFP737tXZszRMU
dTPddE3EwUFfTvXBCX7j56WPWQGVQ/cMxHFdFzGn6GZDECQqWVNaUMk0NBiO98m/
RB3ofzjh/UTOvMJjdv8FVgAJnXLTkgKdl5S/2Y3NgkzZ0FOegibpd+ReP1eRs5f1
YrfvDY7EuWsHahfzQp9Xlb3LHkk5q3zdYpNb8NuWslDuQmPTAtAH6YltZFslSn34
0bK1g6XCwWl6hNu9nIMtRq9zHTCngaESsHvNEAtjG8cIPumltNnGpugclbEPvJfY
AqYxgOuN+4o0BKqXgT73xJN8WOLsT57xQVAOuGlZDwXMQ17l+oEvmADUgE6FvETC
XhrgQOt1MZnG7+3b8DojSEkIuc9+mxcbpXRm+9eLYRzOhFyBCHsse/8K1tV5329O
4d+EX7eZyMBF3Mn4y7zh60vBn1QZrWsHytw3Fg8AvCtGC6DnaQ/tgx4bNLHPvXvw
E355vDsrP0CeM3eMsBG0XhC1zB1BKfQY3keJGELAHxC9c/7F0PTdTU7grnWTz8JD
BNIpOtL6x5lwM/WTpOzxtU4iQ4YpDYv67XVN2bQ3zgumk3L4YCllNa7PefJuqvVL
raxEHWp0FQ1BHunwdIyXmceYMYM3eMW3grExf/BgO391SDxNQYCIJ7Q04fzGp82/
3ILFFOrkIkAy81LW6UUu1pud/UMzr2cmB9JQDONVfrSTr64l38Nfgizvu6XFaUdw
BMjrv2QdlS8ZCnsNsUlpm/rwwwIaa1TCyuIGcUmAIrSpRO0Tvn0PryEHOza6aaON
hjG75JpnQLTN0vXvsKb7XyLfMCd55ta9H4rnk9Ik/x2QOs3tx+TxlYBltqRsqyTS
3oftt83DJjNA7Sy8XdnkETUXPzYNQdxEDiunwdl9bY2w7w+SrtwALXH1MKSSPZu6
Thkn4phEGyEm13t0CCY4D1VdoZBdr0DMaiQXyiWzrGON4JU28oWrcZjfVaibIyDh
VALkGTv9SNUQPOlxx7KQpqfdVv/0l5OVRaTOMsMtIHeJxi+On2W5TfiXl+VOnbOZ
pbwqbXBgpT4gOsBawZbt2zwJG8EXLjJZTkKB7O3GUSHPd8447s1zbMKy5txs7g11
B8Nu5OftbQF+iXukPgyTnlammamDNtZ2wCx+0w6hBeHguY1a5LH0USbbP1JOPAMz
W11zyO3AYGDVJ+vIoPpTxKEDE/DPWBbmZZpW08tKRHgnzYd1gLMVJDAy9cdSFInL
llr03530iUbu8dJwpSmmdnBvdvp4x9g39wlXJqJDzhr2ipgiKy4324OWf5XXbZ+x
1LybC/bxdJdhwdmOZ8rrvprMQpsOmZjHZ8KWKFZ/KTLcPXLu46qd7/aAeRYAzUoW
7fFWyCLbRb73XHxVSwc/2EtRXh3jQK68MhEuOKgcIOVuOkZV0MxhgGJWTSB/D9e/
Fb6aoG49Tr+DEhMQ9+LFQGiTqh1NjuMMkm1Mn3kqQi5l0ohYAgdHADqB7KccwiNZ
eKmxYRl0kd+Udm5ZBV/S8F1n4SeH1JmVlsBXBEqtxvw922T9v9wiZOZZXTCN2cCM
KxJnGb2nC7ZSd9FLjyGqlo98ZKoehLGRQB3Pq264/InCV4NXj6WvDQ2muPZUvBGB
B6qRDE6cwBK8c2P9A5mkQtrIf/g7hlIUyny4dRfvSe3J6EMIvcgQRWaxVxwzFgeR
Gxp5UknoxNTgGmvo65ltelXqCbA7CVeyInMu2KSnDqBdrhSl7+NzOi753eYUjmyx
cyjVp3FvYvj8zKNpFMVqQcs78aJqOal1m84dgDXMFmhcUFrof518Vx9MWKwaXBjr
9ajochbnt70PAgbzI6vcz/LD1vU0a6uhOboXaxOA783SIp7S+hCW99qd7F0OBsXM
vPSvqChrWOn+0qVGT4zdkbtKJoSfAnPZJpM/WRNXVhI570BSjmiU6TtAAa5rGHuU
FJl08FbJd/rGCR0NaOW0k3Yd64RsD5dqVGlRWANnbsfUSbCZO933+IQnn2HSL9NE
//7C8SbcZy14kVt7vXnSGew+AfRhdkXhprnAT4IHhaLfSrvwqjsZB7SsE1p1s9Lk
cwna0i/EploMAQsq70JQyiAzOOY8fV66X3i5qmFvvfSLYZJpecJEDKRHjCuYiDfk
qqkjyPk0opNXszSkH64/+TGBshhomioh65P0YW6Lyni1fapzjZ3RPNY5x7Gsuc8H
WgpCMO7jcDVPFUfyCZlYIVXtojPrtro+eWz8mDDIw4yaZJR76Sh0NW5uAMMJqfPw
GeNySlX8PGbAaUWnpLFrPhql1vyYoyU8lw/R9VFxWvqik7J4VX0mKiKVEmqiHds4
iqq7zOJO6ylT3/TWj83waiM/qU/RFg0dPWHGmsHNSUocxBTgGb7pvSVJ3uLhoTuC
84XSOq8xcoDUb1POV/VByGxYO3AvpgqhFp4lIS04Hb9vcsM65XExbAXXW3ybNlIP
kpjGDrR9yULnJAHJoK++XlZRkENaysTKRd8q2H8ARc0oJFRgvG/8ZBp2rbWTRrH2
rQeMBdqdigcafwwkDBC9bZSbt3glg2vhYFIujIpVWagWLHUbY68przaxPjc3+QTe
vrgpFbjrhr2ECeBbrBD7Dl0yTmdCcdqrAOWo3vj+Vl62tNAb7npg/IBwkLJdeedm
ux22w8dggNhsLZunuw9yPSthCUP6S4J0/7mDUrLA5f0maekSlRAusTbpIN24n0aI
LhSFwrKNiu/3q4y0zkNR4n7VqYNqIldFtHTV5fSobd0bURUWSui5B6yOzRgZ2iV7
fxH0MojV5mgc9gVaTuCVSVG7qNyD5/x7E8VHkRj878cymrFoKGUpjmlBYscs9XFC
FiqV+kKm3hUb7iXkxC1rEI/ddmMJs10VNFZite9Z7qDm4ioHayCV56EQ/7R2MP8w
vmtxGzlFZizAeK5A28XuubZzZLn7anRaXnOuUG07jiOYK1gMHpLvm3Xju13RBq62
TEX5wYhOvlxpa5qXp9IxgejF6CtRCWhUry9L+kWNkGRsPVvzJ7hDk2i3O41inXi4
7fPgPMkIcuH8mhIM11OaTbnL79O/w4pboBy7u/W03nd6B3YKH4WN6723cd9+dQpo
WjejqDOHJA7GAA5wnTlLlHLGFaZKezKDt9S14bwXlxA1x6j72LUCwjsRe7bSd8Ck
xKPKN7EReWjplWNy6/lkZjF1S82WtVtaPdnajeAlvUI6BpZn+gNi6Pdw8rVJ7aXs
OqifeC43/gzSvEKhfgb5HNHeNXfZGSIdn2vraC9F58K0evhQjkqh2Qk4Ac3b5Ivo
+XWC6xL45KL5AeALOhq7nteaVeysttO40EXCnfBWkZuq4uRgDurTLx5hbb9A+JSN
7l3Oz2aPz7eaiPohKSnV0xkkDbfYTMmbgkBM1DGbtrZ415sWOL2hzAM5BTERqetx
IQrAbqky4LEw+oNlgTN37Db45ah6dae9AXZmD3H3mvDSQyJxCDUJYcE0BL7iY6+1
kOSZcSaRQPpSgegC1lR5L2JozDAQXvOiKbAEuYJE8d7s9pkJOjknGnpbCLEemGnD
QT9t35jkUbEtnkkjoysxUYtjCnr5lQEObdQ56CfxIEl6vhhZyC5l4aK1VSt2vS4d
810Tose2HaESZsXlWslrxvDBLEYvHoE9i1pRyt0cWIOOtywps37dS+cIkLCFirHZ
7BH7/coATqwF/cAZez9fiAU+KBO9c/w/fC2rxdmKA5Zg60zEHCgFpob73VCLfBBe
GGX7tppzVDsDujAYUg7koTXmVS3fw1JdgArJJB7GOIGJsJmxk1Gws1E3TFv+DCot
+rT7VqTfqfsHHWsLnxsPLdYPthl7HpFViXdsh+NChOx7q/P21JDKGSwETvOnWODY
o0XhRvl6n08CAzuM1LlQ3tP0Behr2XDXBPcXPDZk+2qqDOLaEVYaVlceim3AZoLp
aD34BM7sbWDhZzy3NbMkN/lMrKJCdGRTOmmyV9pWBpyP/1YxXwOfE2HNSmqV8/Q0
aH2IR1TT3t+9YczSUFgoZt+Yi+isCxeRFWp1aAR3PEZnE9eLEeqoH09TWY6vNs1C
Eia/OjOD2K9zXc6yEot8XHS65A3gHodwlZ3sSXE1ZgRY2rtPFsiRoWg/KtJ4g5Vd
c88x91CEkOHE8WC5I2qy1/8SEH8jpqlTOA44/2mTN+6Lt8oFxgL9Vj7btUG9WejB
r+XMSHhkTCLTT7IiAf12oYmYB+6tWQMulitDRsJ5gpDPZadki+C0H4iFkg7iJ8Iz
pLtfBzpwjObJpwj3wtTxsTFgH7HWyuc2FT9zAXSekguLCfnCEMu+PaxFGoNaWfls
hRFEtlt6SVisNpvLUHmJZ1Ip4cn/2hvp7kla6NCF42f9nz/47CBgfWF/6Ds4FzEp
+cCjPVV5WU9Zdhgp5h8tAwWwHyXwC+EYG/F2ANaU6B0bsC2ezEEZCfVibWpRFmVz
sYDXY1iS+mxuhsx17PBPdE/ngkYbgcJaFL2KpksiOGX5cLkfPbB/BT7qHs27N4r3
Lxek1KnEcG9GRG3V517v/ubZO6nft+FSjOhT/0S1Tax5Kv1E7kLIwPvyxC1OWG2K
4gag5Xu4WGSRoH0C/F8Af7TDYqoM3+cytMyI37OzMaQHdBZNqnZzliR5GVgJ/ioe
PublNV+8hc3B/pN+WyjS6i8kSkwJMUCTmQvzBEwjvSIjBg6GzvKlyr9sesKKzMnE
UofHC3ujDVLEzuKBAuMWMO768D5uXRn3sWNfhgkqhZsqhVzpCPpXc/xLOulsU1Cm
fp73+uHlITRWAuyg4+T09UbIeaJiAhwh5z8B4L89GcGaHzchMlXzHx/YDG5U6Vhb
GE1Y2bldKNbKR0gWVK89Av07gBfsFJovN5omphuD8hlhkuwAK9MMIbGVkWxTO9A/
Bk43UKgXlWga0OLHnQa34Se+RzETs+v9pdTchdG/b+kTpk/UGKlKGl2WCKnUM3nl
qHujXkWL+TLiQ1BtD43ulW3DH8lB0Eddjozrux3+9j8qxRB4oqwtSYWul4aD1Qvt
yhZTrWUQLbaVhDJHdTUneZKikOAT0URwji7sjnvYFI77vnuB7sAlCVwPXVlkOsQl
NKQm6v4g/1WYh0vf4aByFkd2gl0T9O7S+y1S2dwKhQ1Sv8isWjZFIupHKQlxvc+4
YApgBdy0kymlgFeG7MC2Zog36sPRPtyrZf6xvmcSqFpIVwWlRrhEFbHky07xbB8U
/D3uYC5RuFzhW5hGxqEzyxGsoXyjp5K6lfWpNd3QnjgAdLaw6UpgKToQ7Eubql+4
mF78TRXE7Le9k/zQqftnLTnliW8zezkjcs+7fPEc7VLhvv2PS+6pcWNvmBI/ThMB
BnDq3TwKpvj7h16B+xw93YBj91ivWVNbPO7qU7zKI7XiDMTq7iIbKNIlqPsjYhgf
jd1nbUnd1Lz/lnmMw2BvFjBPJmm1YCXVVIKElaNdf2eCvYvHBNY4B54PSzbhG+bv
vRf/VDeLGAQZ5DTNL5zycKPRqpOfIjph/6JBQ8gqhQcQ6b1tal2r5FVDixpsIdv1
0xJkCe+GwedI7a3/QATFBI32VyGyD7zxM5YF7wGQIXyEj6WQ+NAoRRF496ALKQLe
6+CD9fuCpnvBuvCuW1bKxr3cOXad0c96nGV9K6flCoFI7tBOiY+uxdPkZ+6zDMV7
wS3KKKYXOPXuULyisCSwTkOD5MaVdjnYa8W8MQPzvEG9wMzGSnSoGJhSGQQzHFb+
ex0xkTj/Ce7HaoHORCDi1BAWOqDzxku5exc88OVUxygyPLhZBWCOAH/ZO9cMwFYE
u+bHdyM+2lzs1WRLkyc9NHJi7T5aStiu0E5u+orygQTAvUKqmilvRsfJ+QV3lcgm
RAWO2ITH6cU/tXSmviE7WFvYXJtEmNkxmeWKte9omn05dGwE1izRbnfXWZljfF8r
eJcOKgwu0I5aaFjqyWPp6pFsBUe0mwOpDIdwh91zDupoSGlCit2n0LBt2zDNs6yD
9CUvAOZt+5tnrFTHymcpjf2XAI/AWrWtyhPbHpNduK06zNFYtUlzYXXm0jDmYUAp
i3juW7j4FY8lMATx7rocDBxfGMBOgit0nCPnvAnSE8r8G8zJxrZAsHoUx6eYkjZd
Fizg9bvK+KmRdusWCE8PGt3+Af9uWvCe6Qip054G9Q0/SWKf2WptxL0QrUOGfWAf
sUnf72mdLqeBp7Tf5k0dBKldaH41CGjcpW8SqOAa9z5pihDkEI/pSnJP60Fyehvd
pHU+cpJaJ0MVptBWLBb/BlqK8JnrCirG8MWZ3QgjUPo/wHguqqV/3Uv+pKeEGi5z
fNVOXj03H/VJCYRMUToxhDygvcYbO7xko/vSaVnTIvFg48ehOY/uLnylifW/TXNp
PkhXngJ1gZf2sdhwvANMj/uHGK60zjwWBj47TeFO5VK+jcBGu0RmYa9tm9WciFfy
TZL7Pwq3rf08OXEFjNokQDWlS8/98bvkfIWRZ7E3b4akifaGicfwm+lbAoikgWEt
GsqAoCMQEZF2xEB4XGYg7lfJpz50SJUhX/6VKS+Q1eeWL5yQ2HIcOco9+qK13vKV
AFRvRUErTXTLZjRM9cBXp+TyUkOMcuesdaHOTN7tn9q6jX2aRtspzDk0+vUoRQhU
Yn9idjR9wlJp4JKZ8h4nenSf6MpBNOt8nErbZ0km0VnHLoxCJOK+2kAeRtLZHRWt
nbOtKYKALSlDLp+fR87Q+B06Bf7gpB4j0BNLPOz1qMuRDsN9fU8WWkDY5wvoeONi
Sb0gT3Tnm3TgzLDFf3tKvg7LZDXthMl1LomCcqMRIRdXbggeDTERgGNt9aK7J9vL
sjyeYBT7oBcbbToP9vjtAhPHG4TtoWLBUNcvP8jG557r0hs4bxPgOqFrYAM+EkKj
bH394lVwF7K+x45r15rTYWwMLrODnnOKgapUPSjTKDbYJ/Nwaf2xla81AX6Gd45/
b0h93MrTNWYHhBMuioLUw+XlfWAFscLmjmAEQ5C4BCUuaFPM1iZiYLiJLG9K4EqV
lEhzUoGEo3CpDVTs8evN4Lqwkc/HUKF8IvffHsqTFSTm4ErGDowMmBoOlleXwmhH
pEGWEeXlvm4N9GgG40V4ZZWLS2GCIN5cWoC7CANC1HCMVtJtjRI+T0z//1xWoS3K
H692XSBC/SeVZkt+gos9CQOcowFkaaGgy8SIdq2+Aye+ifLSaZi8owpBvpQEtBZK
6SVoTkv77/Mo2fIYLvjFNB711fw877r9JfbO2/t3fPMMZ+W8dXBQwX1w0BFHdO6V
N5MmqrUMnTn5HPmKh9PvdS4uXQeybrJaXAdp6GP3Nzb17dQ7U2jPKrJjpijzuZr4
IMkp+ji4uGNcCBG48TDnrZBZ6iA8ukd5587M7UWpfHBXZj4XevIgJpbwpdXCfaGi
RfioFZ7Pn12zdaYDcIIvw5jKpMUgRgRMGiWtK+NpewDRefdtsr1O+kxyGKXXEKSR
OYMeE926XznFDdFViUUQ/f7s8hNsY/TV4nH5oPAtCXnyP2JLHm7yMxV4uYa9ytKt
Yfu2loDCi2nK/4QuqUZ8rDBkfRXW6cYx2xhcLNGIA37Fh1wA7kVTwb3/VGAG504B
XdwWAzVDsMsM3+VfPNnP9c22HD1RsxJ7XySQ9lD0cmxzl1xxO92IzuNgHEVU74b+
cUaOTHfZP4JpH10dYnIZLg7B/cCJAfjWdBVwEojfLcMv7Vtua2QesHHoBFRB4OfB
EBPJaBE02idY0ZEY/jk8viHY2x8CwDH1GRPEI4aM6yt3lRuY+AdIKYOPVCFWQIBq
l60mZJwp9mqWtkKNaX2ad1sdi7ntPC+Kn6FiEtU4NUKnrMed65DCvHJlxVfntRHW
opkHiHUQB5o+ejcDSQoezDoOzkMtGe17uiZ8PH5PKr4P467/Zsgm7Ok/IjrKVw/4
T1w6nKo6ZwPxTMOTSSbDO7f8C9rbPtQ1WOoW12MGTSqrxLBkT3XTOf/jEQblfnqh
wucnryz4L6MzjQ6x+g6KRJVhPjXcPnDX6JMepNJxijTokrxj221o6VCQk//D75Yq
gnrpVhpDafWCe75D4kwSlIpg3PiiBCSdo2Olxs0pb5AdXgwvgWC8Yta7fexsHHdb
XBKP/Q2KluMMJiQUq03zcKVIVUo0sOgfDZPf5VAg7LzErZax723J9pp/flTssNkk
9JGiQvaQ5f3W4qAoKOXHpeZmYqS1Q2dovnVNaQ0EFWMsloeBSmIdVYNYfSb7BCUd
zw5+YGIiIZ++mlt7pj8BgmTcdI6J5lUhv0YhDYI6Zz9l4qEXR792fVVeaPvQPeXB
LPwC36tkqWuYb+59ZcxU8pqTc7sd2/dhoseb7a7TcRL03syi3Fcg+/UaCbXG9Y+w
bj3LfFWNTY+C2TwUoxrkFAGe2k75208PA/eoHjKGCsIqrgBFuNU+syurEKrtSTYc
/ZSPn9o1XyZRGOJiKE7DXEKNtvKRGqo7aUEmvQx8Ngkr2nEEtme44L5tAjZrpwFE
1pA9s8KOLufApML4E59iVgyEI1KQP4ydKLoWLDgWd5pJAem95AVejSsN8p+wtUf4
galLOVpSZOz/7R5kqKdlYN471x3OQ6yT8+J7/hDuy3mucHpfAzCZ3QCDHMiqFz3d
bWaRgiU5sSKv65xEHCmEAM7HzDisbdDuGuqHnisCoURTkXVfnu4bIhDm4C+hAXQz
7K0zSMh+Z/W0FcQAwjv8RaNc5+jrUiPlx60MhRMnIPMAPftrDfBmwy5FjTWxwGeM
JwAoT2OMYYQqmwGl7oaHVclNO9ZI5wsXXXjIobxJSuEPzE1FGs4CwzjKHUihTtAA
A5p98BkIo+0ySg2ETdE9xZAA1/ALSvVmKKAJyCdj7Ieumz9xzvOmowLMMJ5hlFJO
44mub3Dlxe/+RPi03QbwLVvOZt4N0lvNouHt8iL3nijk7DYg9J2COMus7JsQnchf
DCthJv+dzz5aqnjrxBHJen13ZljDUBa3w6YeTSBkuEP/WDxu8bvcOwTPEyEw9WLs
63c35TkBKIw+1Q6za/KH2ZKw+iUwgmoEyOijDm8rM4DUlGnoSD7UQ26MhrKZMFJq
yN9N0+nhONQTGIbFeOE24NGtA43pQ2a1yMbSTVOLRIXTujSaKvW4qkxIpnk+kMjR
RWD5H7JG4d7NbzVfAWdr3BsVL6Kw1hxR+NuO4VhvVkNWWn/l3S7VP9+UdBN3u5dF
ifRcfDORWLnG2E2Y92af4zqknwLgGoPsNeg1VNvK+dvw/6WHsXjkzN03h+E0Wetr
lzPOY0Xgih2R1xq4Gn3/g4z4lbcpQ6cIS8Rqhe7wM6iM5nuxJqUxeDHbBk93U7qv
Yd24Ojc5p+7JOqu3rKvBBsZaRrl/gXVryHRc7aTvJdoZsCsVJnK851obJjM+snmM
Rf9bKgf1TStA28+3XHpG/N8jaeGyquPp3mpzYWpuuQaC3VkqC+NI4cVMX/J+DvF+
lwydlzqWPkV7lqk2tgs1Ryt8GRwMVjWq9l8JzIw+KSXq+8mUosoHGdMEZKfgThzM
/zU1mHnK+KHDH47ZuSQjAZPQbvAAQof66Mq+Mxcx44S/ov8Zle6L1YVuzYh08tEC
AufHlq3065BuPp8zZT9sPfekIQuhZERH889yaR0on3GW/G1eieLSrhQx9OBSPBrw
fF4Ds6yVE/w+BF3Q10p+moep/FolwTH3gJqpPGg97ywTHMyejNr9/fhJOOXk+LpB
cnrXq7bKNAnZCHeP5TeH8TBYHJCaXHe/cncZUA/XJ9YtLtiG4bq4yHAuXKIvOlCO
+wLJgquDx9Vot6yCKDCJI61S9x7d4PvefT0AcYOLHrfutzcOGNjRByIqpfQ9Cd+j
qfR+QPJs2SqU6tRALom/NIlZ9BQlGuopqDUQycimlfdCE3QAFuEBZW2y6jEa7Enr
4UxgQXY4h5CX6YlO7U9nJwqvC0TCkTPK2j0dkrYxdJMioiCR5viTD+paawCwjs9R
dU1J6TqWLlf5tLOiB7V/JgM5kiqOf33c/clZ12M5SnL+GOv4YUPLuFdbbECqjKcd
a8RpNTLLN0OIwT9v1hO6nVtPb11RPGIehX4jtTXOxmw+qTJ5MLBKXnSUU2MLtg07
lvjgjfkZ+1UQSfNQyO6QtJQA7Dc37q7cUyzDDt0G0kD9v9qzBtPYnt//MqF8ncjK
U1xmBQkPzItPCfB8jL5u05ygddLFkvHF9Fi7bqcUsGeN9czYF7nb0he6RvT8mpUF
8m1ZDFYBZ6Y/cOhgCMqABWadXbockVTBwJjzy+SIZ7RVyuhONmU8ozds8em2JvPS
KW0Rubl0j5O+/CrJP0BXAjvAGEsMPKwewECbHRs1CEXdJz+vKheTQwiYwFmVG5a1
ZGk7cgVQjPUXBGTDmllfBbacXrPmsx11VOQo3ydYhdIW6BOrfJtzq7/g2M2IVLVf
rdpZ1tT6VS0nW5EkfgORbVtzCt0hkS47aGL19uhbQJWIDVITPWeRK/8JSedR4bR+
o2PqleG4CvqxtFR7E7BHE3VHQ2qaG7Nyx15tMCfG2bFZDSG7Dr+TIEimwz3GSnGw
+pXjxZvs43w7w66mavBrltsoK4kMDbANZxlBg86HjjBPcoz6wPZNVY75dFWP2EtU
wSs3YJAnfIR8WmM5V+lQHP0LRvAl9uzeavP/rJro8BuZ7bSlB5F6/J5MRk7rH2dK
O5I34gtnkcC2c8A+LqcMZNn8C1qH2u3oM+UCBEjuiMUDwI113MxeVwwvYX1PlJEo
kHgPssQA3SfT2xgfKaQ49UFqE9VJiFdXrHPEeUjf2tmHu+Pu7fjdfSANrB04JbLo
LvwXvAvz1V/Iav0UQIRGDT10rxvqYA5VObpYD2ZgOP3u3ZXQ/62P2oNcwsDaj48+
LglwExPIkEiwUVUMae856vzTYwpMa/hp4D+1tuB1PGcewszK5xRnzngYYh5Vz9SQ
GCKhfZsFSpjXHQ7f16AGB8dhFNzkWBAnH1NeXUFrzJ3gn3I00dt4b0YXRz65Waoc
MiyCc3GeXE5qlHTdkV2Q8Nfz6NgtXX4hXEX/e6+8yB9/FPXNlOsvrcinFmHusxEU
wRW8aeD1dLf4TY4puI2DGZHPSaQy7BsT+ZJevMFfSmlq9Q3ILMTolptxetELDQR5
qmPIie8GzqRdEjBS1TD4ITfbbWY9vmq1WTG2KSBH+SP7Qfwfp34heE/bnmuh1uYA
ninYqdm0Vcw3cbiWeTkiR1LnDK4I+X5ZRBtutjMiarCZp5j99TnhRXYIVqvmjC5W
YhR4hx2mWjeA7eBEJYgAw3jEWkEF/WJOcwba+J/m63T5tpZh3MpcfmKonlRvGsKl
NEPlyOqL5CAQTIChskyS+d1JvUELko9b2yix7D4Ruyi9OeRb0DKqEhrO/UT6GE0i
3Lnj8OoRiijUFx+OZQgt2BsApOOLb1DOuYABuxyGMFlwhFHS8zP/VnuGI2IhX2Et
FsPkpTFHj3r++i1gpiOL7eRYao7DcY2WZSE7m9fd7qVatBsEzMIfnWXi3ZDQ8p6C
l1SiuxFufkDslt/ekM3WA9+OPO9nXFMOkODAKu/63HA/CfT9fC99sOCcxgo2hnUY
PvlcAGULQeMdvmoYdESJa4h1SAvJg+e04w7Hso+0c7RiSBb4wcnBqQkxlEill9O0
IaadrSzHEAiqwfm2dLp5SDxbZQRZk7j8w7FhsD8qGa+NF7gT+MD/UvvscSOvsEmp
LyYw7QhEtn90ucv6pyq5+Bw84vQb4UQ8Dhcpo0HsgpZbR0W7f+Cu0o2Cg9R2mXaz
HyaFpwaillj0brPcYghcNanzOMaRnamam1c9gn868n93m49K/LDQ40CFshcyZjQi
O3IGrHFH49Gq+yX5jVtkLYFl0U0fhIlc0Ka5LXZil7HnykvLmjY7mhPDQDMR8H75
Qt1lXTYP1llZFTocrWq+c/Yl8NA1ERRNORhcBQc/yMyigjpR1XzV2qLEA+aaYrnO
dbM+uRBmTlIWQwAFf7MJL19lXV4IV6MQV+FQJlCqctAvPrO8h0z4eGoYlsU4z8Vk
g3FRfYonKka3CRm5kTyqGrSfOBMlxzQwN849r0MCzVInOUsoVS0WTN2Ok3AENPs0
0gDVYX9nYbZ8E4BEmpgvniG/4n1AczgDgzNgfy10GaMt5LeH/+aZAYA/lWRwP4qv
SsX818XIOk5DDAQSSCcHIYy78y9S3xq2WwtlJ8DIW35IjwPGhpXti1/p+AIIRjFt
PyIHr8qHZbZGhokreYZGp5KElGxRkXdzkHF5CLddyEKtUFCeI2KzV33OUzlBPxvK
nclqQl9Gt6F2lxNiuLJfqzk4iLgKp6fsVrW6CTU8ebPwn8HdZD4xhhS6S0RJTUAC
/7inpB5odmUKh5qL2CXi9F/VEmqobYXxnAvu7rEWtDCKQwIrnbpyER7Ew+/6/RQm
WHPLGq1qDZNtO+WMnl8pMsx7Kzj1vmwnGGG64yJ8yUPpqH30Qb5L9VDWmRWVOuZ4
AGoCfQ8SilyFSN9yVSsshogx/kOnVr1kdr45oi/d8fU+VtRIg2/+vmvFwmuXsRDK
OhyWUml8hGP3+bugIispxVme6yXrosKlwe4UVymcvzkNy3E59GyDh3TeoxKeE1sj
uZLV/9cH1Ws9RKgFt37xnxpWvu9FNe0oHY+5JHGyZFZPrS0dJ/uE7vxSZ1/VMrmr
fwuep96VROe8uqh1DCag/Ud63oMOSGWCMUQsP0HWT+QTj1YSXXmM6jssa/Vgrdvl
N1Y8nGv5wJ+RtYSSEu87M1qCu0FAV07Dvh2C81gJmIz82KzItwETjPu/okAzqueG
qEjoLM0+/qFB08KOKF34A2H0USlqlPgzcCdY/2kFiq7DJ2pfDvbRHfAi2ThSt7AW
W6vESCmWswXId8xrMpk5gm/WzQWffmCk9HuM0UTbjIfINnRX1m31mRm/nRrob7uS
8WzaV3r1/PMID/gGDz9unqB95cw3lt17KR2RUgwLZVy5IA95PY+inrKF3RX+9oUw
BwW5zdT5Bqw+qb03tvep6Hh9eDYJC6dOACcwR4kzaahn57NxA9i3RLWsm07228UU
cTfaSUrU7FbIaY9d63OFWfE4WwcK+d/uWQlTtckQOPDbN1U9Xi7q/7kwMP4cE704
PpE91c3r6psyecP9X8Z8eaV4wgMzrA0ATJO+HLFEFbVxiWC8lDJH4KItzmZ8HaHa
hBzdPAbadW9i+vn2Ep6fTRymkpmEyi1I5YD6xDSjZntzSAJoEQ34MaWZHLt6rdKf
zyrjNAtpBDZOh+GFecMLmdXpogJUlzjCJKT0y8iA/yhrQ24yGKIcSigK29M4Ezyi
AA46czI07PliHPxP+/4Cy85AHUP/acJd0VA0wml0+rX3YDppqofRg4uI3PfzblrB
z7v9r6GFCe4P+scNOYMVwllNXWvbvWYBAY1rpKgAfBjN5PAVeqr0RVnz4b26wPOj
X4DYjruSB1v20HVpDNf2qH0i76Mw8r+MKW0zYT1uKwkOB1rg8o0Kp92gdmZVxjIj
qaId7LIpmZtujDpdVEqtNQ+ENvIPs6xD633zwXs2WBv9TNw11VGpQlLtNVSgcs6V
mNWw96LGrIohbWE6Os+MhTzpa2/SSaJSRdGu/Xi+Gux421Lh58NcUOYqnDodGUyC
QikcJa5VqaDNiO0rzjxxJ4/1B8GABGUTqDPYd4y9G7OkZ7y5cLdBWJimkszgErdo
EoOd/D4bSbplBTdFk/cuHxiQN5u4Qtw+B11k54oGgj/0TpWVpUaEWPZwU1IMYiNP
R8fOjmKTDaXOYhcf9FzDegAvv8PflBdqjLfJqEom/f/IudaIR6mOp4zpWpbgUJhS
/UkaEhIg0J6Otsb7cVPMWlOG3bBcBWyMPcTiBqIp1H82ypyvYax+FkfpLFkKMA98
1ZzfrHfRqDo6lU1JNml8bS4Mu1xByeGT9zdtvK1GC8lrMN9v19I7baAEq5SZPINk
CIgdf3/uhEAexuWjWxUQq9VXAUFZEPAU/GhQNxV4WuRwJ+NooI6ei4YA3TIeZJl+
k+FbjIVGEc36+jovlmOV+Ni4YEkKx6LNQROyZZ7hUA44hVXV0C0PWUMplY4+5LUp
7FCj5WmkRHG0DHQB4aZvfCqfo859O5eFTukHF07LxvAnOvrcGkiOvkoE5IXMLzNI
wCesrUcKf5tsA6WxSTpBRquA8fXpuKv55J8daVIascTfSDT164V07A0zDiFYPePx
bzn8WFtxZvW39eX3WJce8qO8QZjbHBFLJMamx/euCcyqGU04vcs7L19qZt7oxcav
cvZQ+/33XPo7DthdHgUFIacmB7C/dbx2x1VFGbVwfTQxgmuOMetEzMkjQYH2VA7Y
u+MHdPXpj6OQDSZDrwsbcKRs9Ytpvg37sgG0Yys0ISvQaAqpaf9q+ZQRSkJclfeB
On8HM8wTq6Nd0EYifWoFVQo92V7WG/X02JxRg+6SFGXPB6Uwdwp8Nr8T8xDhgUA2
LS6N33V188hbgaQOfQpx/qgPbY5VC1NlN2FkYMJVTufhsbi1RQvou0wYyyszaVjX
YUUlNZMnphrf0TNpITgyzthif/wZRmkQKpFruejc5KQxc3pzqZUalKOp3VEprK8O
Y39rQN+K1LjFwHOEFADFDq5tMG/cj4+qT8GwjGObsPEd5VbAM+PS3119KjdHyBrj
OeN8OMtSlqmsz8308Nh6LrGFyGP83apJ2lmAZ4VN8G8VHljSC0CJbRVhxlSHhMDT
aKCQ8l5vRp17tkj3fbR6CrOPFyi6h0o2tUyezYKvBe1tKRvfS8aEcth12X3NI6uG
vbAkHR4Q+50CKtU1NVKPIGpX4r2m/3f5O6fC2JBk3qwlrIcnM8rBqXSu3vjMOPPV
P0VcGUH0kItxC4orJ2clTquyqUuhqfx2Bsy6m5I82hhdV3ehayCNaQ3Qi7j9GExe
SvGpy5cfcFzPu2+wTCUTTlEgRFh+vSDZUtrl/0khsNJ5Q/1PyrzyxVpTa4TzC0Bo
DqsIFp/Rl0VkINuKeA90CI9Be1qpqMLoX4+y2Hf7idnQAh0MaA2RPa7YmpXKveOg
mUpCAu4Pmc7UJNu5LwnrLBtH2c//ZSEOtPETLHySdsG4sFFqWlyLMdOu8vJLzapu
X1m4/qjR3YxgNSlY9EwPw7oX7lrN3soXESySodxhJD7of+TVQcuYynWDl1SSwYls
ORx4bKaU4BEpos6/G0ozzqxVTLy9N6/Cxf5vcJOLit7sSBdzNRVAMDUTIZQ5+hy2
Kuj0d4S3icimNNKRQ5dzmlWTnwP58AiYGNmhsdKIrU9alXLA2fO04Pr4EtkzpQti
pHsDKzV+oMt+vbKqrM0+BAtOoogzhmm1wxs0qWqzqHLKegW42s9RVmp3mF64DCdG
fTD/CrXsWZorOBAn+2YZ0QsP4ATPMdnvyWz+0AwPamgCpRms+9HFAtLnTM8Gy3Fb
KM6IWJaH8eBrGNotbi3XJIMwObgIF3owOQ7ppxsAAaYa+CJQ0jTnUPGXB5xW35Ku
zPchJmQBOlj4nqY+pm+rhyAk9PTZamijZGXlNeiXEAmOSrZRh4eLL7j6rnaG4LYd
5RgaCu66m93hLilUMt/ZaccGHmOy+M/x9XsOZSvWSevMtZuxDNHwQt2ytqz6T8nC
Zu7Cb8KhmFYF+aUlw0RFeNqx3+auGYSK5x7o+O/1HzxNU88Fe1lyWq1+jkkL17xh
PLMcY2Ry2qrLS5VJJxjOf0rUyXNEU0yR08AO9W2zSEFsTahsU7UtP4V/zH8PlC4P
3puMoX9EabfnCYmYmVuIlpkFUzmS4YNYCIiTf+15IHmpfXIfL6td5H5l888X/apb
jV++sl4eLty6T6sUqLSGVwC4d674cEZPgHqe5c8eNlQ/R5KJT3+QUeo8Wa4atV1W
AZBDUBfC4QTXvN+aqTf/o/EG7QacUrFySqcKIEE1QjrdGge7PiB0iKC7BBqgPwY7
B6NKpMzc0R2mh2+sDnun843bIi8lFr84ElLDuLoXIB2dxbdcEIV2JlqOkOLSp9WJ
/eapwQYKte3jsOu4Fdr6RrOEthjIKIOhZ8YbPMgMiTrLTbQLN6d1udj9fr5oHQ4X
4C/0em4+a30k9abaOiDu1NNDuvqHU9GD+/EPwbW7G/x1Ru5OwsX7CsVcyFK+jb+F
ApV+7GRNBLZceZJdi4XFkCHMaJQoisbiy0x6BFIQDgG5SeDyr6/w/2Fr84N8BO4a
ms966D8idiIzJNIm6J/HjuOGdQzVrdRKdTO0SSN2qAwt6VIzaY4IiSJz+htsdt+9
PwHOxsGlY+BXF4IrsVM0EGKVTOvFqqXAOot0ic9fRJa8ClMihskcCvbWPJ/JHWTl
Z+rGx55CR/GJv7TRke4I98IOTnITATAK0b8IiTFy4qBv4i4nQN21Ynb2iuBk72nL
2AHPz1QZUQZJa+7/ZwtMuCNzugvtQMGx1tEx0rr3fNBB5c5UN6lZ4Q7o9u7ISbLT
aRqlSaRgLUkAvSCaJnB5pDupXxZzNBF8ZIz+dOF4ofiUZL72NgYWNZsKi18opIIv
4bwkYzwdrcYzVWZqnsf3o2g6CZBxm0g11b/rn1XpIsvq/w874CRpurRoUcnyvLB6
PcLMI6FqpfEK/5At4uSKrXFoWuRWOlmDOSvq83U36CfOu1HIH2trb9OGh7FlK594
Ucs1wmIO5VYEhl6PvQX6vD0yuJLUAJWCT6KC5wsGrgk2bdXsKAoDAmqHj6E4VpRZ
uJqsVDb8SE2px10MQsWJC8vEbXoC8qGULmCThvasiihtrIW2TgG9OQdXKJQu8sIh
Wb3pXZye+kbXLAZKwY3A9M6ibtms1Zblbk8G+hosUm3XApJCg8vk9QChU+7/m5uP
PR276kRhLaMcma+jfAbf+nEQTvmhAd6gXRH28jOrQC4baqVpV5RxJtsJ9fKKCsne
XPRsDbJ15QWL063D6kU3sDo9g/W9p4QH8OxdM5LS+p149VhSwWTLYYpOBN9OXtmq
c/tJnV/jHqvvGo4Ijq+VNGJJl+5+JzOKCzWmWRPh7kdF+avomjqOqMm3NdU8P7i+
v6uqb/UECZE+dG6OEpJnInZcGKx+Pw4Q+J9noKPBUvQ4m73mGZyjNoSsMqrJLj0v
K8Rw1sguxUra+CmF7bKO+4Tf4KbQrL1YW7UDmlJIo7pUls6ApIZwwKYT+2bjAvIA
6b/APdyyZ21/PAtqSFpGx5GYnUaiyzNBz9sg8NNd79MOf5Ct4Z8B4fPnZ5BxTdIj
VibxgOtsjzKk9EZMKqesgWEVTF9rxUaumRVeVXxeQMRFt3V7AgpQd/Zx9jyhZyMg
lG9+7tWcvywhb12zri5SPuOfT0f6DTUc4Fw4vcCFHUk/Kl3Eq98BhmM5dNjlmwUz
sLiFfbIEDuBUR6mMwENW+gKQp2iIhjiJhsbC2Da9AptBcFsc585sgs3+m8Cmloj2
TtsVp+UpNzQtbTMFo2SBF/p6gHN3kdi53DogofB/iHJEeX9Ddkn9R2AnPwtBscfo
c1Ph0wrzoMHzEEvFo/MlNsOZpa3AOBnuU0qilOxFZfmO1hdaUY6ttTRsm6PZCGMS
MqF9mey4UJmpzxLYbS9dc70f9WJDo/sZ14tGrmSFAgeNEA/0ixkNJ7aAKUwtzVTQ
sU7MQtiv/IOHAO1OV+XPLQ6lPh+F6DWtQjpH0rJNKptydcPX9Yhr9tZAblh2bS5k
P3pzveu/5B3Z09Otet4htF68KzlnHSq/Dm94TmuAYkpPmf/Jd4liX5pZJbPyVrDp
s8FnvUpRpveVXT4fGIW4o47WXHr4k2JSPH2jbvnOEitIRcEhL5kABI7smYujKxvX
Kfj8OFbg6232pZRT83KCSKz0CC/kjBTE71+nmvYfMR/6Cqt4WH9qLDbkWOfJmzkU
8BhQEWJPeHwjKD8vNmiTXBdln1wmj3MysvunXFVzaecrOxA68j9ZQ8bDSb/Qa+w7
vd7TIjJJ8jLojZFSFAT5Y6sFN/Qkb1MB8YQrEXmu/+7pePA/SpRTbwqmSfPvbDd9
EytBMZ6NWt2pBObl6RqaWXtNzWIZYEL+TOluHC4hu/WBLYbFuqTAEeJBjIKT9QUY
dfTcMtKzUrvvYDwomMGkDrsxQszbAxaaqewztH661oejC+Xb2E6bDh+byqh4X4J/
H5DdHuW/B73x4F49hCoif1xYiC+LPacOKk6d2g8zCDvVBDkHyUfrEy7h7JXr9Max
BS80S/ijVnFX6REtU+sH2J/kqdxyWUiJk9EXy40N8eiIgW87EJSgWAZeH4Vg+eED
H6WNhMfK2R+XCNqcCSHk/iMpXWglOUObEE1jWczg8Q+uaHlty0J6KJUuJRspLjmd
pQ2bqIeAhigsJBJ8+NUesRmgTKKuAjpxsMwHjizn6Dj2hPbPTOx6nPDE4VrVQb5Z
F0I/1ot5y4qAjMtBKhoNKyIJuOhNY+HaqaW8+L42d/eOJo3Jp37QX12ahOiiAApp
zSdx4JtJk/Gow9Nf3biLPS/1QvqaXk2ScW6SrwxQHoByr6e/uJD2yuFV6Dn6F9Ba
GaoT6sFjZeXu2G0xpBh13NVcKYCmtBwDKLu3Fg1yi9cFAIuRoFb6xRwzQJ8a4MgX
kN5znNmc6SJxZScoMDo7VlgZe8OE1IofNO/49IU6+0Ws8051C3P4UDyDVGnV6o+w
MgGoGBNyZxEVVCmmsANub9amDS3NMTnLKnZxnfe937FZZNuA/f4PQ3oAvOF2imdC
RmBI2SivhkKzgMixqQc4LWp6gCZvAlFhuhe2O9en8wGhN16c9OwB9+scnIkm9wMZ
tmpjUsnWqvwTPqFDNykNMblYVJNKAb94QRtj7lrJhYmbYaobEdvR2CyloO+Xb+OR
e6V7FsIUEGPUBHCtslGvludgF70ha0abqfW1BGRDbWTbR0ci+IjwotcNhcfPvJln
UMoU+c1H+99C3r8pGhWjE6mpwUzViJDItCuzu+Fra4r71rb+H3NkgEdsWbp20FOw
wf2svn07XdOIqMRoLwUiJKY7Jd5WWXQd5UMFBTCmAgwY1fLdeyPjhVqi4DOOc3qQ
l91rjoGQPEdo6gc7KWY26j9zB6BgZBII6YFQAvLZnH3R9YbKQZoi4zmv8w1tk9BP
oY1s5g4Q3sW200Lxs6XrR4sOS0JSXSotJQkhFFsyDu/u1kH2YGZK5gTt5KS09Px/
cJodIH8NZxK/qeam1t8opHTZiisWSxKM/EcFhu1ebuVUXGtZyZUz6njDubA0YC+D
SoE3HVfa525dWpqzWU0pnIStTqRb16LtJkcOiYbuxBIiZnX3Y3CAnb0J58+g4GrK
XTiJRqaaCQMuiSXLMBqwsniVS3YaPZgNsIAQFI9dzGmWzI2Df6lNSGYzhJQU3loE
AKoMs7fN2JfMB7C8N5GgBrgehBHiDS125QU4EYguzTphZgtE23RWx5JpoiXzD2km
tmiwnegmRvnteoWBYgTVe5tKSmZa7f8OaZC1Rv41/IeFx1Hl7aBcy5HcbeBiDu/k
t9iA/3s6QBQqQvbMWLNEqIs8rNK+T3Ut3xUUDTj6rTfaW++MzqALgjo+k+vANV9T
umAtwJw5Eng4NV+lJ8MG+iDUAxIAf2wxM9Y9DO024dAUKTFdD1Y9vz91WDrjTVP+
Gvi9kSo86oiCL6ygsNWrMd2wB4pQtFrPi49NZJCe4LXXYVw7rWFYlSvM9Z44mtLp
LzN7BMdKxVO8n8YvstOTTgqEWs5THZVAsw2811xRFh3Tf6GWNhjXayyy6UOVyA5P
TvhfQcdP5lP58S4Q6OHb1zbNhhcyU2KivmU3HJHOGlLsezRDu+QvrehVFyWabHG5
Pt/UhXoWgotdOforCOTTJ6Niyl4cMtbM6YB31bGzAT10lNl0TSn0rAEm6jvxj+N9
7DSucrzT/ZBzzS7gV2xpCZK1DqZpNpogpQh8l52xgkIVFbtBaa6Uuzdzpu3OLnWK
iEtTQ2uH2kM2dz2T218OXJKO5FYiOY9bghKDZOKd8AaLynshCN2K3Sx1LOIAe3cf
+VRHpLzaCVVzkxBwLZoJdt1+wbSpYVTmPddqHN7Mo/sWP4lWZ/EtKL6ZdGQ/YEZv
sIoXPXyI3z5q0Yr0hN0lx6MpedHfasD0LCs70d4C2YF261Cf5KZschW+E/v526DH
fofZs4ev4vicbUpPQDAekEdhVdQa+wsFF+5UyQT8OPFJattihQNUf3KtUbduSD8y
sUqUmjT1QGkMCBHv1h43DunqXXss144m7ASidaYFiJtgahRM48hI9Cc4znAAtAMl
UvhDgxKuYpWMdwBndVVL5UbD7IRGM2yheMIko5vkiUHFO41fRaHmbItYLf4v6Gi2
SL0D8tLnPTikBTvlcyJMfyBJdMisxUnssx/6tjnxlwsnpEm3LBpvGM83EYzBxOBT
3nqqntjxMvSv8DtIR7OdGoYzm4Xcewg4d1vlVzy3MI3bKB+0grLpkrR6uAzu0qTP
RiZxn+mp8GiLgccE6w9as+J2i8VcJPG49gx2eQpmzJQjYNvVmnAv3UQ8ExTmrH5x
liM+5IXztZU7+c8p4SchpYqhiFF1rXjc6EUWBwkjaxYGtuFr59w3zOahx6Ih6ZeP
wTG+NWbGSzWHUqzYCdkOAf7CrHvUJ8C1ErfIacRBFg49qLfDE2IdVDpsvagJCGNc
onfC6ZYs+VHBXkMB/CvA+6onoIn2mWaUx5UQnHNIkPKIU4RFSxv4MInntejDINWE
DwEkndYmbVLPVQ8B/k/cBSh6DCUdBaGq6Dz8gBumRyD16kpOIHGYxlhURR5nfdGs
DMVB4E4ka3mDEBmFu0eY2+vnkYeVxybageQmFkxyYjIG+hKaIJ67poX61GlYeozu
DSS+M3FSsnveRQJxTHsGilil5EzWT2bNv/Lxyz2AlZubxBPhEnX/T1zC1/+QWbl1
7hV3UrNPRVYRL6PQyTm35RmcB4/2FqWbkKYJ6WknWLrEKHZd7hi6W94ofDKSh1ZO
8Z4TVutMuPJCF6k9rLj2vqXuO3DEI+u2PqrBd1vtbAOK6JpTvo4L8+TxR69Mb2td
uARObBg9+PlIUI/okM+nAfccNnhOuB05Rj8KMkow6NY5+hHFmGOassIn/b3ioqwR
94/1EUj3m00Wj0uTbDL0jrIFwLRDeOocBnk9Y+Je1dV7TMOHO8wfATFZIFTZX9DO
Pi0jyy0dVE1hpOOP/X89VFdVEYoXgw9f29QO0RFF5Gx3u95SLTWWEmdSGP65jcQe
fcrDjXxN49Pm5LaMsbCJTQvwDEHh3Fii8VI3+KYlTqRaHqE8+n7vgoVRvHwEtfKA
KIGfFOFI5QFqX2h+f2siwkhdCKtbbPltj5mAvLajgvM4lKqbihxjocMzgdHHNZVR
2aS3X5lEv9tyEI3A4bn7NXoOo2cZZhpTKFbBDfUSw20ogCpo85RqaDi/PJzKbvwN
+Xeg+FclwVBVKJvmExd0AdtyS5nDsJC8+dFTRvDPeIxGew9znqS5rqgdZ83zbbqq
FaxOO3gJc7MmiGfEhwzwQSXoaRQ2bLmAug4fIVE0E10OkSYTjokRWIiclmWpKC3o
HuzRql+thAtJPH4SAW6ic57lHPtHyIp9YqTh8L1PI2XuUkBFK+45gq+xlGSMPc3r
EtYjut0qmd2flaKg7vBVBqxk3YIsD0+XfCBRjPXq0eHiJv8O/hy0JsyPOcKE2gL0
1trR3aAJLTmZQ5AW/W2XOc0qgs+PIpSbhUnF69lbPpBrAIxq1h5VoF0N8aSEnKHm
MMDJfkuWjBiSCLdY1X+W8A6PzjvNWfFoSD5kO3mc/50351psQ9Nx33Qar0fC30Er
2ySb+O+j5fZahGMcChtJic/085/yJTq4J312jalRYm2Os91vnEehvQWoBc29Ub1d
ovGyKHAcOrdGL8AXcyxqrvLRccG+MMwQVhEBSZvKk7HtznP0dKsULaMxq5VjgSit
Gw3X6IKR1XsBLb2wknC5a2vURGq4iFVcjTFjsv34xrY/6QHcjsYg65MCVUbl594B
Flo+v53XysA7h8U6HH50NZBzV+Im7uvmb+eFa+1lhvxLnXTQw85D72DdcqNWPsD2
ne9pcKIEajjFGi2QAlIjhr4F/z8/Cy/cm4n9G4K04QQAmu0GCh5rzkdCjut16jB1
QSNw63fVRvjtAyuiV9OUtPzd6fhNEpKNZ9BE8d+BjT6Q/PNImX5Lp/wA7hq3AR8x
sorO/LJFKLIx1kaFeWsjY+uf2O1O/NaP3qzxSSkouKLBljkCSRlYoeKSc+/2ZqnF
AkryhitRrV/zQOEyF+otIVtihUfdgzejSrcwdD/2CLk3uyvxwtbkZ7nFVxTSjXAa
gbF3wZOFxMs5Fd4Z0WpIm6c9hMrPx7qL91LB0ZwztaihF04OqfKoZW6zryCeM0Ue
gWQUU1PklD6hmmpulxq7UnkS7QufEDwOmcVyaA0i9DDPT2tCIKG1PsCzz3gtULzi
/nsiJHzvlpB0T60mSlNpkUzpUbw9JHDfdikG2fwyyRIPPZq3FuCxLsLScmsvFJlC
ehIhjuvcO4mGAudohEpP0234fRmI5CMHlzER+UsBx5+I2ok6ZGFb1Goc2+UGDdqr
ujq4D++iuBayI14/2AShXFE7O2WO8oLIyyrkDidl5Cv3CM5wuKoAQ70/0QHsugiu
rEj0fzw5DfmuE9diBAm7R9xgR+QWFpBxCKZ4DvaLsl2nrhIk2iURlunLaUNWg4n6
kQR7LjCliZSVxmMKUwS0VZqNl5qpxw5aNTm8GvfgoJJkvwnf/BUDyt3XEnL+oyBt
bJvwAHrSV6tFuH9mXjTOstBVnB5RUTCa8XzFJ2btWv1ADTod4eqq/tlmg0auB7Mh
sZVmWzLDatJ0b9e6N4JsDWtZ4d5Maw5X1XKZT1OO1OIKEl/6IP2vBz4pG7BQ4a/Z
jZCjgGUsrmhDXFngp/wz3x3UZoUl00a5+z7QKn0CaClQWthpDUcygluRlvM4YK3+
lhVZoggTU2eQK5fHKIypzbPK2C7O/MnDETCFWyRVjX2kDOF30z2ikhZrOYjGOKKd
tZZSnWDA5tUP7gGVHh59VUWLWaX7mqOjh1qJ8E/8jzkZ7qH4sTfwa9dmfxi7ZliF
1dCyoukggKFtaZRphA5/hyIyyVYDTIjjz9Dyr9+qMYIB3AM43BQNRwFXhCBXoBsk
hPJMsG+BhUsA8OGNjjuiN1Lu3MMNDQlWjvfZGCrpICggUdpxrM4q3I3qim6RqPJl
3YAvxia3CjH4HSiLmOX7eFusIKap7vPZ2ywFhB6am2dVDZCN8EpSHxFtCpWypgWj
fn95vbZP79NS4dBSYKyKRmBcMtTBtRu+Gjo94PLg1IjtSp4Zmkxjn9bIhjmvvTw8
87Et1ypyJ8AEKnNET4cf1N4BskqXTihoGrBL/f8kLYjccYs6lg6f6Y+Vg+zUrXXQ
jz2XSXYhll8o1m9uIXHH1LShI3J/wm+M1gMVc4QwyFqOYIb4/bfmGhC2Yt8XBOwx
rZgjcSpKpK+NXp2AQTM2IJlGYW5LuKeHO6RCvGdn9a+Z0aOWMnX55EOHE/LqAI/1
KNIsYaPtKV4hgBXYc2nFXpepcl4xB2Lw9JLTtE0DP4jO0mMVosehX0K3idoxNf9T
ei9sqsx9kezmqn758zCZfvjBG1qZM5Uuu+hJsNXLPO+tPa48lYQXaMI+68qtAisU
wzpT74dASBgUxkNhK1sRecSUIZyLSmkuuU1QlCLIAfKfIY12xRYdaCHiVK1HJeI5
g4aTAlMX557n9EQK99MjGahW5lE7GZdsC/JzrTaOvP5QB/wTHhFj3+l1bfqBmaHj
yJoQZxhEEQLEyLo9coQV2sAZsPn8DArtCzj1Ng4l59/AoS0SHeFon1/gzn/UnuLk
YmO9wyJHArgLvXjeeC/ZDDSnoxJzVETIfhdE1/U2RXjHEMMggfQ0GvJWMZWA9ISE
Gsc1NRfTmOuzQuBwiUS/1wHnBAALUUHOfUDn1J7Jv5Sa6ycPGohKNMCxx8Y1pMZD
5V2oZemzugXodD3wQsMB8EtmEHLy17SXal0UNzf0CtgNDuuy3NT3Qik3PDerFr3x
Bm1wOUm8Hf1kSq4rqKrCcOD7bKz/fvm8SjDxgnNv0TdVgD8H3Px9Npq7ctMVx1i0
BpcPTbVK7BU+f01CGdq3Il8mxEYbk8wy+w+zy18AQn/OXeRImqWuxPgwBzztRKoz
F/EtamzXrWNa5jygUDBJfOAidxhegoqsRVP4JmMwaFtuf03sBajGLzo+i5rEFmUx
u1S6ja6UsACnm7fM2uRDyorg/AsMTna+08Y4+fjh8+WhiKrjGLJjmiNCIm0xLPTt
oxtKOKMFHUIiy66tEYSF8i9k3OdlDbJJOBWdllBQA7fgtAy69gOR1pDggxZ6cqzV
7XEGOdcHNk+c+2iEZB816X+d3pOBg0wWhvNPqu9uQqch6h/K+qVUZu/2VCbSr0DM
N0dEjcyLgoRQgknBKIqVo+Lg+tnfz/U5As8LqO8JazMdvx+rlv21B3luzOQYsD37
Ww7pZgv6e1xbnssjataF9mN8Fp5AUFuCz2z2cZdIXdXRmktYk2ECNr3TAI7TMWGk
ltJQ8qVOUFzQJnWxDZgvwIejnJjDqI22N9ZeulTVHHR1JiaDAk7R7frM5N+lsHwe
Lf41hxuSDp2c+1VkjoW5V0pOC0wZ3CvMUoR790qsvA8l23+9hHCq+l9h0Krxn8L/
h4fIpEL2k8J61pM+TL4m5A3j4sGaai/Yq9Bf5MDtp6xmbsqGvI6gBWFnQAKIhpej
NohwegsWX60qqH/YkBKbfrfl8eHNmfjAlUzDUBPYUDTp5iIF6+wWyjs5eLYgTLPp
iES/ejpfE4MxC1jhHK2uoW+Z6+JaPXqj/hyHgqOs+V/+xHf8IX2FeBM357eZK7Y1
LDmKtMOEQj+zW0bIcPv9puX1/H8S9E0QM0Z7rnYOOaZYaYKUGqSp6b3/WXSkq6Ua
Ptf0boD501j8Rf9VRrzRJiT1YxFOAWXI8S06XY/4e1XCBIhfeMlI7ttWfcZ81qte
mM9yTo42mLk7KnRymUgEcDh2CDIyC/iqQhUvyYNWz8/z65GJfW5vPgqTj3Q1q1WQ
AjhAcUtdXhxCLwZgG+ttFon9dcYlPGa7uxRHhECFrFDTZJekp83J/WrVSh/PYsLZ
pDYQ+HyI2RVyvHN4ifoRzmy8PP2eP7LmQ2aDPSS2eTAVzbzdZ8d/2CGXRMiMMyHu
JvYlGQof8+sxlAWsleMJwInjMQLf9Q2GkTRRTPoOUqma/32fd9fw+omHsLyPUahH
q82L+Q30mfTrSJ8h1gp/gjh5xJsalshRCSB4nsf06sOXuaK9uRVR+VMC6tePYzoW
J52qpxZHM8rDUTGZ33miOnPbkWfls72kmEfezn8nOTsU1bEa1TPG0EQBR/rvtz4O
cNGWNgAEVxeAJMz8XOWuTwbIgrasNkMjVWKodaZy93BGTtxqzf/oJGvMJhtT3sc0
zoyBl1woey3wBJ7nebu/XJf+nsG5cJgeWH9DLYK1xYoj9KMMvmP6rgdOFeubg7nB
UroQu4gBcci6nBJAZD+lkmYu0h9eUBpfCDzlG8bugyMWfC9BqAfCxDFleC8MOfrF
GA5iLhY3QkHn+6e62omUvinF4j9BOLEfbuCTfdJ6wSXFIBS4PEk6WqTIn7gzQO4o
07uYMLzMnsaMhTldGEPazm4hcGH9kKbt8qQ7On2BZYVmlA90TGdT2gGrA5eqtw69
FBh3sKzv8CC/4O2rzIK0ZP2Sw+XTFdsBk1ItCTYsWaifFIMscKI7XDu5IDXHEVEc
X8fsa/zF7h4KShwHISsRhdvYmitt2eQawRqm7gEHQ1qoOtkYn3Tn/7xhtT+2OHd2
yWjGeAiSUNIFhCVmfFy3Jc5uW5MyaD1NJiL2dA61pLqgRnfReIMHCBbH48jTES8A
Kel3fr6dXZ2U1jw0cd/O4dD0188oet3SBGDcYOFrtaVToFOD6IMnAxHeHK+GJXIb
DHMonQG0jFAuCY1ZFUM3A47sF2CjNbG9l6lcU+y0aZhas+8ydeXG318MLknUYBmg
vx/sozHyZng8XifRduQ/nBiNLudDLRGNzE1U52GguWydXAVmT5AxvUfzUr2jg6nC
4MYddwFjRE9kyFAqAaMUibom5IFA2Z+cN1SD/RDhcuGlnkj4gKYdhH5/BGrUamig
CeXc3jHmfYedRiqgDJERI2+iGtLOOeul6F5Ucmf1YMPdNICMwvHbZZWxJ9eY0DZN
MzIb3nPSiM93mGbJXVSFamLTAezxK8htc1GLBd4IinOaA3L/kJVQbtHvE/XDsymK
rBbMhX95uz/NHt5/oI6AccxnG9kslztM1HxQHk2ZzcFV+ORBugQGJ6plEZjLoOUa
rtN4aaYt0dUq2TCvJwVQuc0sCiKKx4/Kx1yTz2VNC8tm24t/F8j/iZi3iLHydCKs
HY4G9p2tM74NsYb/SkCSOz1cQ7XarU1gctk8KyksZgWBAs8xCMGhH8QeAsY2VCGS
ZjMuhgwSOT06qXD69R/TWrE+WLf6o0tHgMP1U15Melir1DYfTtIQX5Mm22fb1CNH
ub1ac0zxnxZeefzjLBRVijsRhT7mRhEEjVYYg+71JSmSM1iUjiNKK9EK0o0vg4l+
9pJvSetDL6Bca8cv7T2HTonv22GS28GIw0oVOScZ0oICUN3t3n1EEc+WxHuhhOUL
SkaCmhWJ0Xh3z0DzP7QTck7/lrlQsb7O/RZxMO/U5i/NNZZxgDpLFfvsUPjHEGWz
hBUO3n85XJLVsx5ycr8ZtufsTu3bUz8EYcqCNZ+Q2ycukQxo/Fjs1U4tPYRf08RY
nNsNrcS56NatAzn1seqknAo8RrY4uhr+B0SMiW57seM85SBzQ/u7iVirVIDez9ui
0G2+MuVA2P6ylDix68/CJh1FDzxYQi3W3gMTBnncC/uGIVILyr1FzfX7thb42tUG
rpX10WIOlit11hZrdCsXJ/vJ3ELGqyPtaf6ZmjWjdfquiChhyQZJSfUOYBfwB3zh
DYfK0CGKpYarLNh2XeNF/oKVD86JIr4jdgWBDoILyJTTmSYkh+PcgAkLkKvYAqAW
3jHDN58vZEv4k54MEmQqmP64owfklJsUL+dQwHeGJokdHQX798KRgsGyljfPuX+E
0EG2LQAbx6AYwxEnpZYhlEGOpkaco1p2KYr6Nv5MBFCoL7HTq++dZMoRF1yD4QuE
aSsO+rwN2GZTM3iCuV5hpD8aHW28TtlZT+ba44EsSKvdUINt0giHsHYbxlSpbBBq
WRA71cBr9qCfVaik5+zHCG1359ZAh4m+onYv+h237AK8wXyTneKZ11ZQaJwfdFGe
EVQ1fREjAvem12uV4hSjBIQayWmE7yLCEH9t9Pai4szBKWNQhioeldq4bVrFMuvb
iCYK+/Zi7UTrmUPa7O2TGhHveBO+0xwHPR4z1KlcgBtDFL8gp+blTDO0VKxF24M8
ui1sxCsfbkuoqloIOqyf9BZWBJXojf1aNC6ei98gfgKrudLNYUgZZ/k0lM5vgRv+
hWd6PlwsLGcSBAqOlduNNM0nm+hJB9tPFPuFXshKKEqW3W06qLP3KVUMfkYHl9Wi
HvxA1fA6H5dNwujDiGDWVJ70t7ZxleC+fGS0naMz2GyGoD7xo2986GsZvZ5guntA
MN7ayzO1F4Mr0u0h7/9LbG4kKlagpUiWEhd0UYjGfONhJvTiwWzEs387bavPiIpr
C+HO3CubFIULW7jfkCBPUGfUf7aSOxM6TDUilvoQssNR0lgjLm2VEWYfl1AvCRa+
Q6zlffzxiWgAH3SZUa82HIn/YXzinNF3KwWGMJzyO09ugeZ9+YXRY59vNB2CRxCp
9IjjZt2yNKyVTnDsuRVEAi2ffQa0XO/7wHOSmlNyBI03BdBepfd0DCwP1BuDuvWb
mJBWRpdCPNBsi7wHqd6nYip2TC/SXEpGHCuhosKIn4SgiAa7ybjPEqDFR1afbbOB
6XtHR5VpPe7W6tPiP1ByGorBQcjqamTnvoBg191yetofjpNtiJp2tU4aqdHd9B8i
pgcwLVYsxLRpKOGt8+S9wi+BJ74knEivGCgUkS6y3eYFIGgUupXtI42qsXzbaqJU
Ba+nOej6br67JLB4Nvmn6kzmonDY6vFu0GS8Ki7HQl8EV/rZr8/4KJNjUqoG0SO0
kEYk5fMH5PuZ1DbbYLDp4q2q/R6+Lai/xQ6pGQNlwrhLsFoHRrG0J9JQboUvjQTn
6uFMXT5pJZjvB3RwsKLVrn+Zlf8j0VG6Gt5PVEP+EFS5SE3MkS8us8xua0VPoha3
9FXKqwHFVDqW4KeLd2AoEnAryY3JOVYCuLIBeAEt/OTwkjV1eoEBw6FFTN/fyOQz
P13YjOPBkddTw5BaL8JADH/3FE2yk0NoKAw3h0iA87rTDsTNreUXFE8edu81Nx7D
ELLAzhdCGvwGg33OH7UhQjxYPel5lQ69avGAF6Z32Dm/6x2fE4zezQ55HMjlkJyT
vknA0QEW5b+fS5QZu6v+xfEy8lCWv7A/g4pyRhJv/XsHP9DFOITXUr62z141I/M0
X/moGUEfL9IEFSORT+lsvMe4AQesTwUIxQ8aZOtQxQZAmZKPsSPzCqZo2VF7dXly
bl7YCj1Tjm/cHQxweTz+yotUObn+FwnNmo/M8xWYdLCrrdkNJw0454owsIc6Zm9K
chIba+c0Dqn6NRKJtJocVSuJuXgdBp50/u4hGwNbDPqEKMXmWP6J9MNQ5KJmcTmL
8SOkx+Gr6Ig8kmKWW9pMNJg6hd/+s9IK9vLGAuWjh3ax0Ncw/TmPmr9qVdpoXsk4
pGDhcbU2tmZtcGW9Zw8DwDqFH44axvO7yCY9YsnSJWCykzz/WOMy2ZKFsyMfnOJU
i0/LgDgl7BxHLYH7xppzPoeOCjigg+ehd46tBnIs+RtFkDBFOPpAorAc6ZZlR+s3
1O0z1iX8utKShY1HegS45fGMI+nSIEhqCtnGCbYMoPJZprLhUSEKSTRmap3CZPHJ
TGHOCTL0BV6F4Vq1xSa9/MGbkVbmN3c/CUMY6f5+QRKP+2QdPab1ikFYfYDRN1ji
Pu0yU7jbW9kKLNklPVL9BxT8Rq+4EwcKmffeXas1tH4Hcp1+NafVNc809g99b0m6
5LAIFGZ58Y9tpNkT6f+PCC/edPDn3JtiMp/xZPchiep29i8qzZVTuLvc48jBP1hQ
Dj+2qK+CzFg5DfJMHw2sCDRIc5QxmmIxJE5iWDZg1bpJpP6/2YQTrW+KdnELHHiK
9kxjZyOmyXqbVsefncD0ZOvIA38NXuKQAORpcNEGSch9//nBgtLMHTja3eAQV31W
kIWiiGaUa1quwi/pAsQjxKaFQhyv15o2tYRL81hLvg+eCDU+isN9ERYgko8msMVE
ZFGjbGbzsu2aIO4Jj9sd2nn2Mp3ANg29r22DQHlgu9eKLzf2Ywhp7etDz28TDjP0
dcScndFkGKkzkIwj26II6+AlTHhEfNSOhsrC4PC2nPs2cwTydVfLRSzAguLk6JnJ
IiXZFnLGimWcqQAgGPli5/4IdMUdPwj5ZE1QUEuUvxtdIJI9QreAXwSSSXPStqcH
ezrRjRwcsZgcD7yo+z6AGceSiL/+6VRB+7BNAbS2EaqNBESWr9l5bMVctB6nVRrE
e/h4QxFyphByWF36Wkd15umijhMgjjvlW8EpzJ1l40LwXKR21dVZx0FHJZ6AmdmU
0R/g+XJy9ydYCaUA0HWKQ2Zk/bZqh01KhNswSh/KHByNkmxm2PAsyMA6sJUxYlXT
W+a8Fub1TkufeTcHUORwkaWnlszdhDLBDju1GjTGd3Eg2XyMf45gXWbX9MjrmfMS
ywESq+zU2MxIPkYIzYvAh8miBDqM/gR8IDkxbrUi2XzszP6PGKomvl7SVPjewyt7
a1nwMkvGONgq5GOEcX6/9i0/81QZh377wf5QUYyOu9l9D/QSx1qLGxFDpgzSaAXS
dbdSCixpQffSJQCnK7XDRO1LY2ENe+hd5Uk17ZYZTIT5vunePjnBIr3zGo0OFZrU
/m40mLLjF/Nd1nEMYenirermNAIzOCpLf2Px/mwrRGraWT6UkT1uEUCpPIPKXZv0
8z2KTrgcIkjGNGD4qphekA95oY8qsLaP3HTK+EytlSIZgcFnLfdoaXXhdKBUuXB0
gNrwbvgMIbTjvWu++1l9cJ8GY8QtqSbNG1mZFQ7J/GoJgNslDy61FYJlOJhwJUlx
Gk4l9z3E2AtPzEx/KGkot4CWXsf5HfuqbnsBpwhtcpg0Wpmn67lMBJ4JaJM64rtq
7FEYslYBcOr1rNAXvIBUYGhyt1zIf2iEb/ZnUfWbgI4ncBPAZAFBnoFsgGubILG7
DLvDl0eOTaX2jjIXDR7zK6PinfqA6oQLvz9ZnZhCsRNFxEavLJz+G6Lfcy+NZKeB
mS3fHtLB71J83KGQAVcmD6dt+FEPlwBfhPJ1pGgsETw1zYqIBnJ6NESnz4v505i6
qxYZuHfbUGqEUq38QvGB84PqpJwZsqsvxPJVWccIQkZaa6JH9F62yBtyCLHsyTyA
cVJWvjWsunx7FAnY8TGd5s+gI8gWXThPJ4MRbNvbA+IES3IJ5nLSahKJvY7RzLZQ
OU5QmGOJVMIPJxWqN0Tv7jWO+HWRiLw4x1M82YrglQhJMbXWzGWXc6ZYc15iH86H
OK5W9qwA69mXyPkg/pJhTRmt1tpAtpk1yJLzjW+OhLHSPZ5ID+fAFGtdZGNc7BdF
zqTYhVJOOZF/46O72L72Lnuj1eNvH24i+czm6+HooeJ4KqOLtC0sespnFoCzfg9f
6o1tnicxdyz603JkcLSSjDySYAXkwbFjD3Fuvjx3JVNRMVSV7x2SXlaEwj+i68i4
m5r0vUT1yeYYfYNCDjsEhAGmwAFnZgTLD7+HMWrhHJDvVispxjo+LgSYyWERUcTG
NCd8PzOO3S7yIRfKsLPM4+Lq4wumqc0MvRnDb3YLbBH8idWDWa7oIxG11Q3l38//
gXl+pStzUtYiHsJprNsr9V6xFXO+Q3n/eMnlEmGZ0Zu0O89QZ06PgrL3iPORzT60
AeGBjhQEBaKGO2hKjLvOkUGiSsUKXk720eThoDWz+TObyaRNgDYpZ8crHhHhFIh6
twNIX5+VnUVQef5kI8QhiTPNEfqxbmwdQo4SwmOG+LGMtxg2HG1F4qyVt8lBj/4q
nsf59sRyKIz4gdmFGBgKOaigkmxrYUFzVaalGAG0fCEU2O8TFDli3SvDz4T++N7X
GTaB2Nk0DK9CObF9+4sBXK/hWMmdtxtWLSWF9ndP/V5CrdUqQgNcZCfS0BwcYnMy
GXOtv/ggoCA+34iWTpHfO19rre8byMaqxkBWAnQMnPgtckConQ3eRqv0YPill3fe
mTrW83MDbYl9W2dsXd87cmlZaxjWzdZewAaoLG4RS1EKdjGde0rbMPg0So96DxJ1
OszQwTBy+GazUnCK1vOZx4X5fukbbd3SxUN0aipH8J06oShCMbxtD33NWWFEli3G
hrTu2jHwfQsz3lBKPrE3bu/t/5H2rTZxCDWGJdHytEHXUCMg4oNdUx8xOs1Xn7Bq
IzdsH41rckKFTFxQqR2SA1mvA2FyGzKCi/a3cJL3MBBt2QaED1hCcEnVDrqorkP3
7bZXbaMBggqRQGTSUvr2mDaPawds++KkhY31ZERFV3cAx4Z7HKhfoLAuQMXMd7oo
ZgdfNvT+jKqkyAHnh4NrbEiBzz+hkeYsAMKdfGRLvoTaNq920PSDjwzVyP6SQenQ
GfW6jgHzdXQPhFBq6Pp72mZg78brWU+aXnl86UOX2n/oBVQewTfHR0q2ONICErKq
eARb5JMbXo8SYf/Mzn1CKpjvm6uV6tA3sbsoxp7MVlgw5aKQH164Ihu748uLGG87
7wvvxkYMD5g6cOInN7zw7e7KqC59it8p7bDqDtvyqS5F8t1xAJGjRZ5mztZh3M5i
ZJmsJaSOOtk4oia4QWs3G84owhqdqKofMq1D8qeAnMhiZIuKobZXiP5ERwG+f5lg
3tAPxew/Hs1wQY8yhtSxnmOCRttYIBlikHHpj6GWP2syjLSwPE+Rs1uSh5D7CDLN
p+TnCKbR0ibariRbvNgqKPtgNJd1r4C4qMedJvfSqsoejZl1b2UhCnZMk+Kyu7SM
NVfgTJVkcEjtC/P9kCgAQNx/w3sRVqQ5UCNHHZaS9n1JA2+bfMzqeTu+AlGwL6sS
Fa12yFg9IunwYByP5RTkVoR3wiy2ORK13+w9oALktNn46245Firyb0QRp/WsB6zg
YoYbg5yZPNtsOEiTT5RMX+bqMwdyvmFmfnOUBs4PPJZnRYWUPXzWZtMpV+syrpAA
8YKF59NA70C6XpvpSD/8sn8GGV6rB0Q6QP4CDIfXlw4+7azGWZU7ixckFl0bKdXN
ODE4tEUVeb2zwFrG5hxqGZJiOi5cY9si3xtm6O4ZZc9sO9ly8nzBHul9OSPBwb4x
L1BTPMFHR/H5/Fzh5T4w8M57MtsK0q+wllv6q1J4e+WQGsxE30gI1i37PTpEUfzj
W7iXyEMzgY9niQ3boPyeFa26P2BA0IYpdlfp5Pn34KBkAAZtl/v0fyxNiNwMh1ps
CL6gtA//jAEmzctEbicowfs/Q4cjTdKm1d7uCHLRiDyM+cbX3agab33tapiQEnaC
ayQdpIFbt8N9BJ8lPfY5aAN057PJZJsG9M+KVHh07Qw2VXvcm2jVtwhP3k5FSsSA
PuD2Kxd7M0bdDwfZQwUVHb3GYwqq6DzLB8FBVhgntH9Lj7Kh+H7knVEqF+JXnr+r
mJEQ1qOGjoyypldJTJGQzmVRGKMWLIIqJ6wz4nj18zkPxuLO57mWjNCRPrHJfJBi
dOEytjF9eqCyw/QVIHZtZl2cJy2l4wu8iw9JxfsPJb6XXqtmTtepFPRMk6vt6Zqd
vbQmtOcaFkWYVW+RsQRTOT0rIo5WN5ugDZU7Okdk9SUaBgdSZnbXRfRkkDpxlvgV
VuWwlQ6uFcjyx9Pnqjsjc0FdG1S0BjLgWo0ooAe/R0YKpX9T5Cj7jyA9KGrfuM5L
v/XhagOIO5InXB1ksBaZsr7KE5cKmyCPMPANCi9QA9ARd0DJrUIHoRPURkVbfJW/
j+Fu3oU4ctzS4Cu0yggIYQxXcfxHOi96MzRgpd6AAifHuyVLQtLfjyVi8r6mr1uc
ba2Vi6EunF920mnnhAWzrfsRsBidIr5mGEipuGKjXhD+ROasPx+b21Ba9L+ZXjYq
UPXr/P2VymjTHw4jgkMnZsBZ9+YCfom5Vt1yWvgIZbmTWjc5usTda7pqMIogZOBD
QXQZXfoEkN5KdjXlpuF1KlOry4Yv93NiErbPrfAcvJiKoQXNVemCpTPFI1jH21P3
GGW4YncBMuScLpYjuXPYxhvFzB9d+05duY7kY1Mc5mBNav6+DcPH5LajNWrSTWXG
TkN0ld4ykOt0Z1EIhv/SBQV2Ex9aoDjw7XT3wmCzVTBLWGFHieOnBB16rbUpwQWt
sYba8ObtZbTT1e8DodfMpg17vqxxu+Q2CmEdKfYs0GKxz6ESAJtvdswIfDd+vMCW
QcywTH0hIul+9KSxYwT94HuPWmhJ3/LUSeTz0j39XU8+X3OAUyncOzyiiV6NQjTh
w9YqkNt2nJKseHaefbqiD+THqycIKeDx1XR8s1/wTUVCj5iSnSO6Qxk1CAwa8vX8
Vj/V/YzXn+8JTZsfuo47/cptx5QQtSgPejeUkfI/rjY4PvPmRZRSZkCwXB8ue2Xy
K0D8YtjoYA1GRolO+oDGiqDbMHTVbxW5HPqIoGAZWafOQz1Xjtxdlw6mMQjVgyiu
JR2WtD0/4ohdqp4MQKUfgl0P2zYZsmq1OF1T/ajghqLqLPklh39Z2OgwHg1RySTc
UTrVtmp1FbAEOber9/cw28VjKoAl/6WBhTsNa16FkpAwjyjYEl1hwSfo7w3kzKFd
ean2z+v9eUWyYRvY1cdt1tY79fkiKGI/qoCqUYOcgQ4M0TU4wWQbTzX+PQWTyybn
E611t+RNYbiikV6go+qQIR86gtnYQiH8mTowM1/lpWcA+idkTPePoXFKAREEnO+u
G/Dm7XmlQpvvYYqlWPc8Ox4GtoFwpro39o2dGD3vUlxJej0PtC5qRR+Wg36QaKz3
dGhfFvPvk7w5o8NTSGcHatWzQll/62djmAj9GoHrtashPtKEx2C7RNpa8a0YbtFx
qsP07VUWUcZgy6zPW/zrpGtVsr+gnqfp9JKNuCCHOUkwMSR6F4eX3jr4to06HGFg
ZTqVza24NuPyARyyVffjhnzp1ukflNPQszMHjYniQMbXoeis67vy58u58LHaOs6v
8S1xx+uGf/AkMhxZjRg+iKyMyITLejIL/otSGBRPIA6gTiXRW5yBbrE/CW1s8vW/
Vb3VIeBa1EujAr+q3ZOFcciJdjZr0pQTgYz2YS3erLh9/jYD1pzqxFmJOUBxZo2l
Y9s8KtbmbJtB8TH6gtc24x+3zpmZFM3BOqoZ0+LqdWJtLPvRR8VIadgfs3+VmjFU
3Gp6GIXRxsmxQYAJAj6cE8lEVJqtvmGtq5JwLAEtWKpmb49kMXObArpH3qWlcCke
1NwPE2ICsTiNdzTKdDJ3/RSMf5fPjDR3GvRCt63+IXuuWeKWpSQsI2QaT4rygp/c
ZLoK2/oaFvIl3wmuX38knD7ULD8gQc7OT/3TJITJkILIb+fV3OTqVhK7K+f9Ywvl
bC/cdo8NevTOkhkhf69SZX00it/zL6rs8nw4j1nAS9ZghC1pu7KFRWXVNtTXaGGq
jDas4cTPvXOEQg0bJ/i/Ovr1Ryr/DHFeCOtIcZZTD3BkpSOjmkd752bzVHKpfpHh
kfoM0Q/E9lSPSBOBhtMf7t8RYnXiY7HNa3/mDZ92sfJfOMDPhCkRxTCAq5ocTcW7
Jpk/e4e1YkFFy0evn8j7lJLFJDiNiYnlZeuYR/IjKww0LsVAEWI3X3y8PhbTNaKt
tvc4L4NQwvyzr/2CuZjWzCwuJ9oj8qT2/4ANS6cZ08jZJqLTqLuSCTmF5OvOCJQ3
5P0jtAYqbEh6e7aijpteYVXEKGQvxk9zKACABG3i8H22SWi7nOI/Ee+8kTdVesic
4R6ThjyadRE9UKcUurI4Pymdizsdb7jx5SAImEXSHdoOSbV1aW3wCx43gWP7OEeN
zzGVow38GbMNHd/pIwMVN0FszTPaEL//5ZmzHFAV6uqROrFEGqV+yK40H81LfbW6
0bkVqSnqt4kbi4el+hzl5xLM3PZ7eLIXLFwVfQg7UvUTwxw4nK8DBL6rKoyXEzYe
R469kW2qqglt/Pcu/hyy3ONCMRlmhrPoDJqWAKcb1MbDNfEkriUyDssnqdVe4ipr
YNkY71yvFp8XgJq+uglm5PVUbLCuulnBoMMhb4CwWRs7kqhzVPyskUQEmwpwbImQ
R23CDhiP72V0pFGn3f0GUClYxOpKRGSYHALtzQh3u0j6K3pfiYC9Bh9wLaxBrKg/
bzrgoTvFNWxbbqcWEu5kW+3C4slsI9mgPKGFkl0rl9TPvsChYEbsO8p3Vp3/mZqU
fvTEpCDoWl3cRTV6WlZNUqiZB7iOXzg53uemT1ZQKep29sX1TVWdCw5zj94WsjO1
nvpYiGScmnHbTY2+6+oGQHb8J8Fk4HQ9QjIBW/YnoV5XUNv4vsOaqxOgJz6iJpug
ZredWDSPaIpc+XW9P5R+Amj2RLSTEqiFh0s5fss57Z6fOKbn1SXYqyVWygajlLCA
+CsGokGdCPSxyIb0ls8KpRvJrS0JAU9knl2kwSk1J3EIBlVafp8cDrUarNhTH7ci
U4nZ9P36Up74jM35bYlTGNeTy5/nYhX2XDPP1uosKT/ADionHuIwNcoWb/ytq8yR
IuGtRVEZRg0xvkTcyKv8wkRKLO2LTDritfmsny/WKq3uW3CbzYBXw1+OiPddzGkg
ygHlQfjgMk8EgtMw1bV00xGBYjZGVv9MNYsaWMWV926g9a4/x0Cyn3WVKQOxKtCf
2Gyn5HS22urRzrwZoaaPcZfWat0biIg1gQcuIkmogWh8M5PTCFEqqDAU1qP4qamk
1+EOSnES/KfZJRopGmn5pIMZ+ZQ7Wyr+w1xlmI/NdKPn6OG5yWDSlMTJctT43Tes
MG8hQU3JSVDzGqQ1o8qsgZtT044Y1aHc/yH0ynJEUA5kgTiAjTuTYRW7OD0N9iXH
c8urOfrsQTDZyG/cmCDQl/JJQWilD6w2QMTfvP1pcrZllxeABmZ4a3bEPRGbGxBj
leZXbz3A28AIDPC5bIyef9mZiXpwZ2qWHdnLV+timjjbUQzsv3+HiBcgvX+P75yN
vqgnlDCOiob8yfqJKoQOK7Ci2A7F1eyK48EMqjwKqqBRcXEPtZcbi802BzPxpvYB
/roJOKWVHqVSEzSw+G1Z28RSOiBGBjmuH09OCNFU6M4BF61xGUmx7/V4hVl4hFq2
JgrInt3YSL3VeBP+03XHQ9tXiDhWnm7nFsk6fTDVcTITRQ6PB3g9YVYBFxaJb63f
OVqCGbaEkD8jArfVXXFd1gGgUb97/C+i/+9+vXyTdNnOu+PWVsbHlZm2/gLKQAbt
OCOJq9/5iqrnZ4PoE8pzMIbBmzSAL8nxutZtmjtkd9gbkFoYA+gXWU2CD/jwVMVe
EMmAyUuy2nN8FuRgX3FXNyUZHV5IiuA1Rl6tk5lugYVvVlIKAXqeE9YGrV/aXiTp
UaWfelOPTA2XKw+fnP7Zb4heqwS8qaiLSxjpXcqORU71eZ59cjuUug98iV0VsmMX
e5YFE8kg63isS+3ea4kc+a122x8ZPil8E7rj0jkeM8CIDBW2w9KEp7ZLNHqoUjhp
GMDeKNKN1frZ4ME2vDETfyq7YTt0oK+dWazJD5PROzSruOYOkK1wYnXXUIFqRF3m
lly1dhIq4fxLH4dCOBSPD//2VO9Bao2C4I//pcYzqPx9KHcyePNDFx8LRLGxgeJc
PvYOSb/uAr8g9H2m7ps7HHlPPInP9ZEXrHH8rfQD+HDIzPCn1hCNUoyEbaGxi8pq
k9bgy6ohGUWtl3uXTe7pBc+25v7Bgv9CRXe9pq0gATlplEkZwfS4/lL90FraV4I7
mRF7xaQhNeinlwTKkldi3ryaiqvzp0bnJnSS9hgFjegdDw1z3bXuhZ7xUy6H2jhO
jpDOB9/8QaASm1sGJQr8uwtKqe48UJqPrnTAzqfmUMLkO6rk10d5JmCVXGo4/3/d
K637Op6ezN9/AbZ7CrpSNlQ6elZE/HA4vJp79h+0dPvuz2v3oQXTYYqx1cOHoV1a
i85uu/HLpUd3lPJzqeWYkMqj+bGKpBgYYzY2f/F1Ylmm0P0gP42cnrU4lmv+P3ys
tAfJhg0elRA5lG0TjmD0zwGzoG/AB3DwqBUefseA2GkDUW5s1Wf8+3V1T0uHot/S
cAapT59Wg7XHzpwOvhGHb9VnKEWupoPetFQIhxwLdiPiOBKj6kMyC/KppIy2N7Rz
Tfy/G3EWt0Uz1qQ1V7H1YlZsZOUJulpnNHNMtAVw05R2cYwFXte9WOy5V0sQzSsr
GS6i0GJc6pPGMuKIx4tqm430AGl/ol4xEbfumU2+TVoM7YnAf+ngwaf66Nzqy4OW
jiM37mDUpvtCFTCEVjS0cL1gl4TU7GbSU0oUS1ZC6OLGby12CVWGZrijpOHphSPw
tXvKGtux+KiLgGfjhs1SwnEch84QTukI4e4Pu5sDzaQW4Bz1gbN7jmJEFgLhZ6uQ
TWvCO7u20Sv2cYJUIaHurErpXWPB3eQ2JnsoLFIbvRR1M6zfi460m+NFDLL68NCe
xhf4UH/iq63DlwDyWFbP8lrxlxHFx8sDGocQBijGH9p7AJJf9iV1HiKYoA/KUX9E
lfABz11RHZ5xWzfmEVsl0J21//GFZ/2pK7p4DyeUa51P0nhZr5WnMtqBfPr+k8oe
boYqB334BuC+RueGOJNSKe5e1wVMz0qQAWmLPUU/AT/PEXdC+pnPsk0f6k466JgC
Em5uX1HpGmV9I6irsjvCk4+uvea8l2bEM3k8ZvAk8sOXIRURgcbyG0fbCToigJ9N
Cr2Sd6zw2SuWBHorkKyiK6ECpx5p/6k8ZAd+KmwkesRSr5NnYvw0K+zclAoAZGpy
WYGs4PXjx7HY5phqsp3nKgsir9SnuatDAd6m30+AJbAgwsBjIvcBOONohYabX0+H
chSsg4C7EayaNaCz+P6BdbfxuukElwaC6n+yY5oyXIrSTQCG4ELofpxI4AV2EDpz
5qtQRybFP0Lvc5TrOrO0SkyLB4h/dfTNDtwgmg8+J07XlIDUaHAPCazTVFWRDq31
RuJyqRPLnxpPFEI35+w92zMaOo74XEFMfr8FDwygxbJNAIPc46Fd9WboiEu0CrDN
cb72iQ1V85mX/adQTn0tefFBrtcB848oNXpLOOXdemYrUtr6QYOjChuHN4zuy8tf
dsrXpYl3wF0P8SMMidHJ1VDOUVY9maM7aEX65ub3GWj1ezIUvG0aTcpWQ9gIxg90
/kqG/j0JFWKcTwZXhxCH4ZEf3FmejbDcgjllSvrvJtpVvwSCc3lzJIUKmeOT7qmy
3cbun0jjVyEEId4dhk2sI/IyS3h/kceVvcLWWREJKMXK1wWHLSYPEbu6dJwdSr98
UowGs8+B8Zr1+ZDXtG8AlFaWdcHxPTb0WfdGiJbA6bADT9pI4TYBf7Q3hT0MN4Lu
fFoglePa1GtzMZ/G6PqXyEwGw0u/w7Uar9FPC8O8e9sTcG+kKpq+66Ye4ImaqDei
hxrvgeyz/Je9vkuM9a7mx9OZ14YW3bAqgLsY4iiqkR3Ot3WykLTDY47hLDT4kidl
xmm+j73NkIEUTXCa9lYAh2JG96rDKAoZeTszf53ehOO7awWTgyh3LbLSkwUuVFAl
HV3a+733p/L2bkz6i4B4uZwswMdcfsdt3nIePGVVvUM6XAvxkUxpbeuXFpBAjpFc
RU0o3TPY4C1M9B7OBaf6dlrsiJLSGnhXUJqEFIC+76Su8Xc4vcZ5z137KA9Pv08N
OtiOMHN9zbhUJRCC8JfMpnyq3RDwh8oxFARgQB6eoBxx2DnXBKqlWPVgFl89aisN
lsyyn+yF/HQvanSh5xhmhfRnZuQX9/lP2gneCnJdYGhaFR0CCkUV78VPNj3ZGWCp
j0psm5InImBAw/9jQ4FOW3qnd1wSCNna7jSVVemPnR5rl0ofHCLCxNWBvC2OrZoY
7+y7Bi3q8q3GuEz4HAHwKsL1Win2Bgg3mLirPQoBVtu8wgj5yfPgcB3DLRFN9qbz
/Gg5oeora1ONf2QtcDB84al3H2WUxzRKiaudtBzqBD23W4snUYX/WKm9f/DdaTRd
DLd+I8oeYIyHxT+F6PJ/RxF//FA2qjZKASJgLbiXu/QzZwaGlwq1GsgFHhxgWjtM
jlJVNv/zO0UV3e7GKAzqZ9GkV5Th4va0m+C/GR2vRmWd3RkdD257ZftA8FvfOInP
GHjZeLot50Yh0pWk5tZvtPX5ezn2RVTCkvRFrBehLc5+0hVZg7FxtTfXq1YkYvZZ
/W+6i4kUDOVAkPrEJT2zhOgNvnwXomwGtMuOvlte6aDSxSIJx1I0GL0GimDf3SdH
qICTMe7duDvL8AjM/g+3LupOA7eB8vaakHMt/wR5cNBY9my0JpOkZYp1bzsmrhmL
sGTWNHukak9bXFZq7pKJKTkVJpHO6uRDFIx2OVpCHOcX+v29ehYpiNrtwliA7Xux
btRnTrzZuGI+BXkM6CL0vdr1yiym3k8+IPBO6fy1jIItqNdTamenOMQw6KxCcsrv
0PO7Aw2VyskfdhA5Ws8rt9b/Kck/N4fmOLES/Ljio+8PNByxvxHE/Os8w06Afs/1
68jcrX93GcQEA7TQ4l5VTgQV02wEPJGgixNFBktWyYRZiUkyYQvzA1SoTKAx3RgL
CPQN4vL6zk0iIy7STXsRoXe7iM3QNScin9OeqOBQ5qbwsP+YjLqKR5nMKKXPAT/W
dtgrDX3kw7f+W7HP7NVD4EGIxDCU1Vv4lyq3aHonEOz6qSoYFA+Pf51Rq4ThpOoM
BDs5/0z9LRBTO9RNZwZ7XMd/sZy9G3kOD9pZAjkS9gnULd9SqlKQt60/DPj+10Nt
RrJR9KXECopECiHry79PPpWp37Ho+wYw9IY4K8wu8pS1sr+KFty5+LgR56R6tDUu
mrwD3aYBiSi6t3fSeX/KrDmldqGH9ugGa0fC+nfU5OZsJeOYhw0xswBZaLtzJ8pw
Dm+cndfqrnWhhFDZOZCJMc+aIMAghEGy98P3fS3hvrc+6K42f4Yoz1CW5pT0+cNY
IoE/KUSHJO3/RX0Q4eqjZvXenHcOTKYlzCeNJu0oRDm/fVR/4hdAuSoAiU5A0drq
ax6zX+GbkoXe6ocu6rJnErKvU1i9z2joGVEOjGBSSrkvoVg29vTC+QbevrrwIQcv
TI3gszNjz6WXSUj17UzgBVigoWNzQdAyz71sblzO0jwde5O2u4QB1cUOBbN3w7+P
80LVkSOH2HqT0ozwBqMgx4q8fUx+5ZILbVAmplhbhA4hUwOYMeLy+Qud3aGsGaUL
fnnaXIG8DlridAbLzO+UOQicC8NdbMZUhGjfbuefnyDBv8Ye1iti00qUt9Tge3CJ
sZ2QYDzSfeulkMDfkk4vkEYolDOmZkcjOXfwLDaMku4XLoZShT9TTWmk1cWl93qB
seKmYcgrgmiBCEwFQ3Bq6X27v95d8EaMFHRo8eXF+NVL0MZnZ61QD5bbu6v0ZwzC
4piWhp5Gb08gyvUejlmtArKtP4ttWkOmDVqdxhVCWxB5yS9MZuDNkiJ1vxJ+qOYd
cAX8RdC7V5braOKkpR8wjKabYucjKKgGtUS7XKvm+EhxWgJb5YBKIfpw0kCITlYq
y2SiloU4uRr+eMwCswwxWmCqHUZvKqfpsCAbXDX4CI4wLnVtVgmxEHFNC5Sd8HWo
+NFbE7IxDquf7UHEKX5Zd9IeQCKo4kosDWyPJ8IrSxX95Divo4ghAvyM9IB7ilz1
NrXICt5VT9g2SJbq2jvYXf42oNAaoI8zlUcQfLfVLAUe5D69b0WwCd4Wb4bHiNAd
xp0rraJnQ30A1QOYRQFG9ROjJELuAY03iL+qIv49VeRqCzKLHaMT8wp5arEI1jdt
e8ZdHNOl1abdC/y1oZXDine9fc2hK/UjwCpzSiwnckDe+itnW3PmVLdInlcS39dc
+WB7NEFJ5U2xemX1azYBh0naQg/plxA83+ZDWYv4qJSu0xELvY5c8od5d3eWnd7q
SES1aOSAqTGJQSTEgjXrRgQeiylrU0ujGr9ig2whn0MAj9YOP9ntZOmBevs/m8tl
wKqrqpv4QnlY/mjkx3vJwraQs5kvut5E/eWveblz6eJAO9FOq2fQiFbiEYEyrk+m
6BBZ24bUuMCy5cfZSiacy/RbfrR8cUFgj6MLmYXOPVA15ZbVbYyLSCK2IM80IsRo
+74GiboFAlIGcH3ZH+Fcet+X4e69KorxOMopIQ+fBdjGXCIrbx4W3hdIhpApXrBN
A5EcZaOFybzMTjB9wMCw4WXKOAg01MGt1fqUZ1k+sCHxb8WUcUry1qHL4OH7pfPh
OfWXtsXl8rTPEytRTz7QIe2pQt57qNqYuipYxuBr4R1WevB+PCKL3J1VVxkrpQR4
Fsnk6JvhQijBXl2gGT6yIA6n9EAsvchs1VhBU0Q/jman9d7B+6Ob616fW+nw6zWR
eyVdxG+jEO0/FHVi9MROCXr8JsUb88rKjbgRBFgo/PXxo3M3LhsC7oa+HTcT1tz+
w+3/UU8yEa1bxyPyhys+xJ8jlwQ84fP28jumSjJnri4+3KsCY562izXLViGSM0Su
+/qr9sYtRL3ysVIpornmauOH0gppaXEwA3N77BCYUFd+Ppu35PtxUyPLBI0RkNO9
5w8wgElchKVgshEzYre9p+bQESLWckdXe7vn2TfccElAl4/7lvOi3bHNZTNtzX+5
Y7O/+Yt0TLuN/dYnBeIysG/0hf6RFYsPsuWC3pxiouO6knE7TcHrBUeAzb56U3M4
YPwD2zvinKFzkFo60AVBEGQk5Q9gJK+GzK3rIdjVGJ3PnLx1gxMIbEcKmM2coEkG
ivVzlhX83hWBvNAk9Kgorb1bshH2kfmUgcRTl1qPY3yuAPdeSbccTKOlw9T2jAg8
DvX/mvpXrYV2m2ulrM6KpI9nImV/xlVeR7FIsHPa35Cm2tU+c8bqY3eepDbdGKAS
xP8zOLZB0lyojwZFHauQ0anTSBSs+QmYHtHS1wQRoiv0aHJwROfO/0b6IkYWseXb
WQJPtFC81BKYZPHtbprmhvhKTRk2e5dr7n22f5aK/LdpIeA4x9zHBhfB1oEHOGGm
/se5PnYuY8G/fELFF5gOuA5WvmFWo30UWqvKHMYbLwbWlzz01fcRau/VixEb+PBR
s6CsUaNR3af/zi7H36zS+qmLpI7ch1uKtp3loDUGJ42emRnjGV7Pch11GT4SMtcr
Bj96vxf+a8uGNCnqLSTOLbpnn/SzyujGIFJBfm+/+Lo3S8/dFBtvpWqHiKPCVxj7
S5Dq1cc9+ZRb1LdKP9AQrzpDec9cUirZfV+uw+Mjy0FE3fbbunAJYnm3l3FStmLS
pSyN0VgH8lyZmcaRwFsxe3aYRNbV5ZfAPpgUCGC+7GP9GLRQ5JSs03bQjMTttrJN
T+cSDtU8GLgtikDluTLOBPZYieREWTR2IVkIonyniQQZRocOC+y9KO58GLUCqReK
W64JPxSEUW15LNAaUXZVWFh4yqcUylw46Vtg4RWL8VO/qGy8xu/tpFabQ6SyJBAH
jzb900KikqfUnCYth8g9t+p2i/jPlOZldYUEMsvKZwj9AHgERggTq8JnqOWwg72l
Ex2keSgkli39RvlZKgL9I4z685gZmmzQinRbcAi1VDk12dP4YmEp6f0uefKbZpeo
ALrUJTWC5rGa6afbjetvulp9SVGTygiI/zpMmHfqG+x3Nkdr/i8QB17U9OV3bHdm
fKI7mGXT3jhCxsEKdRi+eSwJtdosQHspewJ4IFvEyAYzDLSptYvD7zmAMN5dOPel
uZX5sWe+QiqJ5EolEcIR87vLAUPx8GVvLuyIc78KQnmbkMtI3aUx7I7J+mvJbQul
PtU/JoMPnRetvq0/IEOXI5wlvL5bTkroasoA7pltuF3Ke6DA7vEgHygurhgUmk/c
RrFBWVO6LaXBox+kIdupH5LFqk3CzkAgyhozxJRbXpjgWeQoS1KAQkqkHrzKTYTR
gmizfLdPZXFXSY6Db4Y3k83MDNoPBouV23df8cf99f2TY2ZpsNCeMT1bYSx/2TYR
Lf6G187/D/5jjMH44i94tqGpwrqBuS7P53rz3uqLN80qSmnxIZ2NhN/2NEM0ctFK
O7D7svXTrinC7pXE6TNaGX7ZkIDEFSF/lnMPsCPyu+pWJOuecdUmRfUn2/CRD8dG
gBFvo23QwUR66m3BLtONYtZm2/FbiWlWLIru9cII5JIiQE4ylEkaN0uRcoq0cDAd
4PxgRGCa8DMKpQVMhGbZ8D78tSIKPEu1m7CCC6HbtTTnS5ihOZQWb0aPnK7Nf9VK
fr4r6j5UJniPjulqYTR4zjY9zfZDkiPScM2jJhZQgzV2sZQJqWvFuTVVSl9fyS7i
tR8Loji/F//TZVNyqOk23XyHroqJiy/QPTGuv7BYtipehe+B9i4yOooQUFQU0jTl
wVdhgPnrJUobJRvHMIGgWgWAzHVSPy+vE8DF6EPICUHDvKMl67S5w1Ee3TFDmmM0
DP5nu91d+zMW/yo3qKCFa11V+oer0ZSlduQAeCOR7Sfu44kuxztpFpGZj6rEwP7G
DqfCkdVMFhP+7XkKTR2gmWc0GEDVzF7e+mKyjlKub3b50DoMcpkxGacWiIa0DkkK
rfh+bHEpvLpMMFSzz9F8eurarsOnCZPKd0zXVtG2mUfFUiMFv2nz9v2o5NBNqSKM
SMhv1kJJiTT5zAvU2vDf7noJdPt6XUvgrmA66lNI83krAMR9+wC9bBbA4eYxqLng
MX+8BWi9CcLdegbD0rBerazihV1b4yM5M8IJooahEuveYgB7L3eBmXIdzDJR5FaG
YU0mpY5OpIzvLYYAGE9uIEfwiuvxgiD9V36hmi7+VdT/tPaeTjWdE0xbfcgP+fOZ
ouZsrAybwjrY16Ga5psmpStzMHVpax6+JmxnlP7OVw7TIbCwV0Neag8FGl4ilVFs
LEYlxocY6Y0B7ihG2B9ACCFxUVBseej9m6Mi/5ikkK8nAMVOP1rIlu18tut443fW
XGEKsS07BkVya5UI8eAVYDr2j4ZpFHi/pIeJArUS1KD/nVl45OeUX9AxPWzr0+Pb
KuU5MYj7pikvjPgvaDXocAc6bQxKLBQk3MfXYp1Bq/1G/GjDrila2Ia3Xynp7SXK
P4ZJMhqanUZvivIhhGE1Ix7sibYBhPHh7FVyfZeIZ+85UnduRk4S6MmrLn5yX4/q
1YYAt6PRTYHChmz+Omw/3VmH+nmCslmoBKl8dSW3mnk74bfFG1O784N2Va6qEprp
43Na12KRlEznW2PFGdRqB2pmlfLJcOHllin4ml2VRk0yQhPzJTYcEF31vXUOyXxu
7TiPggdVhG1v4K8Mz6sQssMG+PIx4s+CslpxEn4RuSt5XGTv2uyd+WYcUdDBRgE4
sxYhGE4wBm9T+tp/th/Qe+yoiGETzOzfD6mZwbn7IDYyhYfK6BsBsbTRVyUwdJpW
Dbs0yPozqH8U8aMlURl1jPMZWvEO4gt7uDCAfUWBphZKmszV171sRiRrD5RE8rzC
F7y/wj6vPmmGpqtMczSyuSL1WuowIvDyt99rNQ7zSmYpnK6pqsrZjXkEOV32uWud
nA+gEytsKmsY9tdFWedaihsyJFMJgUScyZroPH0yzIQKfD8uscVEVTVKb2hEJLLH
i+zps4AXLwq/GS08PA3kgSku2DZH6IU5Yxi9XXqGoOH0e2YdEuNJrDN2C4+0GyXc
oS3tAfA5ZX5u290boExAxK73tY20yR/4DYeQztF2XCO5bU9aBuH5hSiilYXdF1+Z
NbWvtXIcRlDf9mhVp3v00uJ69UfJBb9nls9DQUNy7ndfgodzM5Z1JgL7MsR4W8RA
e4kJUL9PuB1viANaaKlPAcVS4vDNNsC0lUBc+WS6wb/Htc3t9a5pCKIV8AsVdW4l
ud767PolXb811CwqK3wTKZ9e6PDWZYewebofijm3+W8c8cYHmaay3lHSjB04O4qk
0iqNuLIC38TL3HvachyRjU8yYr10M8/nJ7uRDNtc2LvnfxhUeuJCti+VuW45UEf/
158EnNVRp0dJjQCe/8akTuIPGij+kDG/ha5AsFMs2f32KMjhub9BI6RSKW6RRLnb
azSgFTW6DwtRju3E3M4J7gn0IKGAPQbKKVHMtFdutuUdfUS5xaDAmF2vYgVZnTQv
8EFEHjXG182OqBOPGHbSmrqIuhzXIk1IuD/JRM51eqyRqi+TLr3poj8ITDEWViOT
XFA4+xyL3TaQK33q9kV4QC8HlMOUuef563R4oqVohn/q7Wnh/TSFKMU+XIv/Qj53
zbXJkoOj6opokZiLItfj2WNR9oFQmdAIUqc7rfuSVlGQT/GMuo6gziJ0wivQQeD6
mQYBIhIG0PCnMqdg0/yMpzxWlTL1zyCsND5fn/1J8P1r0cqT/1LpjrK7gX36D9EY
AeBeVdTPP+q7QFmMDkJR76CjORq1hDBzqDQVj26iN0dO38Dvt6PZnPpRzVrxSoZ2
dJF04I1p71Y4TAC86xsFW/BVI5tYPWjVWgNbV4RK+DtUPborj2KW8EScPczSyOFm
IzrFIa804bgLU0BmOrHZ/lwIuBxFpL0elezuEimenxRiRv1uv5rtBsGyV+EXULDC
XbR1WVphY8w+aTzH15lyl5RJCicDWP5j8EUsE6/oTOR1cNnnOFQp84rlu6Qruo3/
IUVQXfGOL6eJmb6/s3vZBAu9dTTqVcbagBy0h6g0SQT4K5h4OmpFZXn3Qra8/2hR
YM6fphVdPlnR3PTII40j1z8QEscQc8UQSvHrlwk9puF4lLrUQYKPadUomwP77gnA
WxQKLZAeSmtZESuclIn0c9ljf4s5gmYymUYmk28hrbmZFkYa8hf2GAlUshhGEqNF
NDLr748OUgeaqvDArP34iFNtPhM7jW3RzFFASHL57Y+Av+3uD2RVV1NudsjY/n4O
ew2aHth3+YbyOSn9ExFhlHAgKfK0MgT6AYxN10u2/yxGMshhJX5PC6z7xpqx3F98
Lxis7gO+xBT7Rsn3kRPkyLeA5ai+AMlsKyQnWyEsA5ToJ0ewtmozF7CvC0dMfa8S
46GgdQiaxutVhwJwbYMAZANqP6bJneHbD2XFW6bl34Kd6jpOajEtwhf8fZAlqx+g
ssVO0SWIgfKo2fcxRcL7ydPv6oCxb9NsT740Htxoeve7VbiOqCC0U8yFbBgfn2Cz
jhT5d5sbi+TG8OxBDZZzHTwDnNbWT7rQ6qp0PRgnrAXKt9d1SsGVmRODvSDFzfP8
Bz37T+HbgCtyOEL/N9p/rc3ICsVR239GZyKXtjmXeHsOwJ4DIXR56TkatbBNFHGe
fAafaPmRwOPRV3fkeRMI0FIQka5ktx6ZKzFM3Orv6roJSi+lJLe3MjpWBZeXkeGc
y4LlopQCKFrZPsWgvcnDQBo5XuqpM8E3DV8+17pDGE7jJi5gXilEFWZJXYSSsUTF
ikylir94iwP5u6HXxmC7KJBP5fYplG3dh9fp3uS/aPorf0oyrK4gAqhXaP5WJWrc
kpl3+0L/UN67/beNp1otk6jPNfjGsavK36YNcg1xmqDTRx7jCgWmrCMvDf2dmD4T
SBbLr9DkWNSPkXSGC9Ndv06wtveCozpioJxk++b6UTN777AGUrEmLKj5T67iVjP7
NtekgJFk15EG+YH2ReIL1nt6ieM0UdQuDRNf4bSgU8pukXxdraRgvg9ELFZKQk2R
NToVAceSfYwrkU3QIg+woTkvPRVCPwg0Vk+5qnUyVsBsw0jgW38dIx4YjKGKr3G2
R0mokOk9ZPm8yHzedf0VBEarbWsyYQ4RedjAIpGQN+PcTgqZDf6a/MUZYuglqfZ7
xowuD1GsBI1upCbENlkniSIuYX0hPB/MmCFNh+oe5L5Oj1gsgjJmxXeKQzZXJ5i9
Wj7k4wahD5WmrbQr+qxvJHCfuXZwCIhnAGhB6d9QYF+ZXPeUYF03WmO6j5ftDSz0
4z4epsc2AV6bWx+sgpY6z3B+YPOQncyx0D4A26F4mKsr7uYlxOWs7fGvi9iv35cP
cV/LtOYJQboAbS73dbBjShex4aJvxS5NziUDa9UtqLg51S406tKkZpGg2JtQR4VA
O6ev95SQjUN4WOWuo+YU/67qbiJgn5iyPKw27D+o67YFNCF4U/SUlfpJuUifphcg
ZGMtfQbDAVZlhhCc+VoLf1qSYByhcdq71EFZpORmxF2LOq2PaTu/VyCyYGl0YbNN
9PhpEYwzrxtjmYctDM0GlF8n6MeSYTSl4YfPj7LG4IM3NpOLFsvBmbtdGekDifVb
AKcQU4wLlspPsSRF3N/324OkCM77lBzmyVIfjs/WRKCmub/wo3pvELJNmK/ShDGo
UcBu8cWz0/c7R7bYr2KyPLdeu6JeICqjaqfiYOoDPLxLe6zblWnRhzpxVnPA5RrO
++GRLKQ13nYx3d7L9Ia+v7HV7pS88CtIkC1HFEzyzpQ9H0Zrn8qdKJACvQ9CJi7w
Bh4EofnQpGQWdiDw2rJFY3wBgHt9I8ZBekTZyZaAr+oPeCiPcntACDYllqkD3Tt+
flBDJfGqHGjGHgJ+6wzZ5aVnxO7SE+xuKl/ceQ4sQPX4u9mg8OumxznjhbJysPkw
n8IeNB+e09Rmqhvk4VlngA27hFpKJwMX0LE4gPg6UbVM1eNDZt2BNC6W9WGp5img
G8IqRP6xWAvT0FSPvxrQKsaX2gSw7j2HsmGaMP1UkmNB+oaMRpBooXWV7GF6uIog
kqeQx41cw3UMJI5coR2ken/A2ffo874hrdNICk9ynKChV9Msxcp3oCd6TXosoPsK
mqLX2UkKM2ajRj4skNJZ13t/coEwZ2tk0lhJMRXeP2J2g+LYsAIscnOQOFzhHOEg
N+m/SfLU3sfW7TPFe169sNhyHc9/L5JfDGctsyRzC9i8vS7VNK6lDyi0AdPDNtvC
cDMcczYoiKGfmRxLJ0vwHVoUKGem4cDbkYYSS0FukW+e9LOG6krU4PhXA1SM4MZY
5vbSTZ98F2I84CsNjN/02JEBRMmlkxR5rSRB+R8ojq5ukgHvybT6gyIyfoOPKCm2
MUq1D1zLmJL7iwyufrloYGwbda+NShDuLMzxsnaO8J1BuN/m/o1zZIFxRtzmrFcz
8lTBu5mBYmkkGnZqqlbVXwvaWlDnzpb9mwHd/nBwJguE7mb5r0n89jJrZ6lkdNrK
aVsfkmP86hq+FLL+znQQxlIH9gOp/3cioKgxFKGRdFzq+ajdC7Kye8i4bPMrgm0c
BcrXtVI8QnKsXZ2qB4GULrTsU8Mcilpd+rNykZ7MYNsNE/Yyp4JkTYEBelwoyk6G
e414EqSYXIBQ6nxde6qbBTpjLBN0Sn4LCCl7djVm8OXm65m9Kr+2YrJJQHkFgi/j
o3vSM6E4hruSyqpokHX4TCuZYixYboxcEstJakHwdI80UM27olXInih/Y4zjVwV9
M7qVjAX2fNd7vwxDrn5TMzcTCxbPa2GtK7V9XgSuTM7BqGGGNMNiR/Acrdh4fXHI
7UjB8MU5zQZv0a6E0qqHh6JRQmShQ+F5CkTDyvFZWrALK/k5yU8uGPNxYlnieOM3
h0OyDs8M0AcqHIrPHHZ4aHrx4XS5qKMY9uy3DIJ17nkuQYcs0ddJD97kBtmYDIq/
JWpy3nVsrnxUZFZ+DW3+qBRzoFvOD+SrrZDkK0IqTLiXo4J6OIzO6+00Ek4X4G9A
HP2GFBoGUu5Xsx2pQEUb9btTTNEwH3Pi1uQvnTJFLrAm0O4IukdxtLVaRYh1lKXr
PRf1g8Wz00JzwAqRH8ZaJoguPUbWP/4vO2x1K7Ej55LbgsIFJodefApQMsP6gmCs
IV6qobsUOHpUEsIgz6haEsHUnBhijLWqx0bVdepe7YGCozzxLdeAooelbsS4a0Gc
PQbc0bZ0UVIn0QIjYD2jOxxzK7WpO/4quFKs5eIc1xD5bS1kbsEZMuZh0gLK8r5q
KsEv/2+esiKyAMUqXoxXtWWX2p5J6gUUFQBjevgD5z55ktRvoVhM1sXYeHWafSAe
RqXo23MOs3q6SqWmCXt9Ta4TUhDHUPYx68WC30ZjqZ2G9svRNyNBSZ2ZsANDm0cW
n52S0A+sVQGIK5LTT901ZMJRHXc8fzfTjsIt3UZE8SDyMcycvmFwxsmdJyXBkwSV
/0dnI/VAalnDXYu28nq4Wzq6jyZWBxlsO+Pqp0+HOkuVphTxEE+UWhcG6v7VOuE/
/L7We3D7Mk7+z3qnetkbxJaYcW2afpExSylRTe3WDxESTU4J47OEVtZvmc+4aQfU
NvvFOAfC1N2JEFNTaQTC6dt4e9YIxmr0Wr9wrkPI54Itdn1DVh8xRguVhkfxB6sK
UB9ESXwKO9qr5tkFTYo4fep5dJ/d9p+3mIfHccQWsr9Cl5RJTpp8k7jFfLS7qnMv
LhIIMf5u8PndCzIVcays72VTrh1egmT823+qAR2S8+OJM0IcUOHQMtWytxeYmeDJ
4bUIzRQK9aLDBHKOrBMy6C8MWvmQUTu9KUZL8DuhDTAUgmPDB3gRCbLOdHinQtR/
50dnWRVRKJFQVLN2A/9hDGC8zIPwcgx6/GA0spVESZhnQiIOXykTQZuXZI83k2OS
+h1dvDomDIqJ9zgYUrSP1kuPpAePJpmTEk/ROg8J4ja+vDwTVAPW0TQM1uOUKsyd
+8P54TMUU61UnTg32xdJ0fqeHEv8noP3Slpj+5BpoCfv4drmXDZx2ya922AXU50a
LvIi0Q4RQyqGDASnaiSpwHKKy0KmVLpVgZhA9bbJBhMFfjBtcxrhNQmZkgBkhm6J
6i4pLpfasX1yF2bdq68Tm7YTQV/dn0RCJjvCpAhOACx0zXRutnuCszjS+HYuwHu/
NsqMDAagUHx8uNEek5e1XvOFKlWRXrnT56kGbu/J2fitVCDfIIoKhzlvbKaALA3m
W7uwcFFoK2PMsbvb9b4hex8ESfv7e8LjOxbUgXxnBiAGBeNk+E3KbWlOwwEjQbC/
5NLYgrqnOTeQkim0EgUHHT9hORLFYhgFUlbxF+4C82xHGbwEYcbnEQwpM/wKJjld
JKdAN67STnNNU2oD0ZJ1Z0X4ai5QweHev4oFMlZpcbODdvqRZ4cwj+8CjEx2sCM3
CgO6TUWCHCMMHQT1m4ojgSiBCXZGYMPIhFnp9vYaKduY8EXBlISJzf4q2Vu6aEat
HYCaUSxvo5nYX81REPCykVH0sYwPQrBXrhUHABlDfGFdLaCrdPDDhQJmh83LVsaI
UNqMxeL26QjaThg5waSHahMs2jC/9OegB1exXTtVXC4trGd/WUuCcinyG2Wvd8KN
G3q9tuG27mKVot0SXurygmJ+4ookU1KTQ385ufAwqKU8OrU2BQobXP+ond94UcCI
WDzCew7epHw23Kpw8avVp9YYefKJZUHnXnTmzMcp1w7cnuOLjh4Iek7zLArrbtoI
Wy4z7iZRL+kEGBuB/b/KnV55EWKb2XDa/tmPN8rXqKmsZ1NDUoOaSRahVeyY4ArV
gVnehpiR6Ln7wRyU62t1xmKrZwB7SZwnmwMUS/VgJG/ZCguGpt+UA/MPsU/zyAba
77ENDYHUAvrwcUfWdQKLdIG3N2m1Dz0jq76eovXlXuzcRebQoVVwyUrAfnfkdjT6
mvOYYkR96oZL0dEoxygfV1zWnAadxh8b+nGxFzePPPVnCaoMKESX6zta4v/xnV/R
tDps0Tf3qPCVKk5J6xdU2RdintLZvRQr8cKz0nWiSiE92aUWsUqCFffARCn7/m8O
6UzMfsmpKckQNnZQ/rSu6Pd3EtWxrnawEZnoY+oNnggDzyA3HbSYh7WKkttmnUmE
gH6vrbUwYhLC5LeMzIidcKcQugr1RejUSF6L7cjUe0uQSoDFcsfWK32C9LevK3+f
9pmBPfUl1RwJyiWWYZVJHdAvsplDrcqJOJUFBQKNosTnIXvAuba7nBHc6ZWFVoLt
DQu39d42NEU4KdWGbv6HLyVFWaHxjZV2p6DY/1Htw9DQ6eu8xiCMBdz4e8GthKV8
iXc2pkgCSLJDlSXwJkh/OFoKA089+dQyg8ck979jOvjQedE4OJslVcAeJefi1UzN
0HaNiicCZmxTzQjEFoLM2jjZAuZSqJ38w+Uh4pzWihtGQJ/p1Zg8+MpjCWMBRNlO
EGK5BPKK+N/TxihF31ySrwq5JI1FA9/6KoylgswKE07p+Qtu01MXDe4SVFD5W5us
Pti2xFXSGwSO922Yh6mEFvVGMIJMZLGQ4Q+MKc6Fi9MAKVbtb6jU6xBv7Tw6HxyH
1OHhYKr9fbRvwqvciVp/Cs+nks1w63vkrizHElqVRfwnkI9EmFV0pohODqmPi1h9
QbNy4oLJR4l2kAhZfBzIyoIy063B+SZjPXJw/u9C/7Z7LN0rB+C4BE19EnLuBYdr
y793K6B+vBBBLm1bS9X46SqwHUi3Yvq3sFWN6CNJ6R+o/3z/dt5m8PHQelW1d0IO
WGwz+Qo/L8CK5HASO4HMf/2WHPDvdDaGHlPQAYDQ7AnCcDrGpc1sCxskSEkC80NN
3ILb5amH4fJejG0FpBD44ueSXxEhS150NggPeS/MiBp8lxNwRI8E3is3Sb4YMth9
TZwOd0/kKdDsU61btEV8u5Pz8HzwM71vwEtEiLQiQZo4CJgbaTSQ+S5cc5OehyYv
OwBC5eT9B33KYKWxhlRMvMZQt3gd8TTXdweOrx4F7i86eyq0+2FdO/CkPpPdvsRK
5i4Clh6dyzO7/0moi1Pgo6VdL+WASHEH7/yVP/DLIAy/I5ZUV3Z0oVzwOEcizaG+
/VJDs6oyg+Y9gqgbEI4a5pyFL3AnSLiXDlBROLvX9fCbmY7AIesP/mwV+cNSBGoC
18LjVz9kA7H3UFyn8w6Vro2qJ6SVcok4l0czLAttGaJC+ViXDh2iA1OTf02JpPc4
J3hhTcJRYtMjFNeb1zQndK1lKnEyodMiCWp+Afo37Up0nmoEvW0WVDhblSB8RQqZ
DE3oe/PwKKpTlafR5fKRtldR1MjXIdnGPG/WmO02pWgQUsvgzAsSuXRz4FvXCeVt
yzsBW9JjdkrspqDijJAi+UNEtGw1YUdLkk55VaLa7UDAezzdAzmz6hPde5wVB0K6
Csz2kFRty1dHZoCFKv60a3kif9jItUa4E3ZaGqcDaBrNqb6ni7Wg4Ile8SRuGCYD
g0LhVb4eGUklgHlO8AbECLkTHf+tYYvcnwnuBRwM26IeuwBcdjKlGxQzGBvHFdPj
V9mj0JQdgYfpoyrCxVdRoMaBOi1mqV5aBur3ADnHWqlZRR+nTKk4MEKF+fdkFhO/
8dvezOUQEVh33EUl6OSwPJpf8ArE3yxbXYqMc1g3UQlbuxsTADwywz08aAMUpeRf
4cffxf4lJUJ0OPeBUtOr5QtQkjGk9+vEtxTRMurICH0Nubnn6ymsnj4m+Dwpi3C3
n/93HzN70REHYuAw934XyEvzXF7f3u70mPhnt7Gds3xRcC3B9xyubSfL8W6OKW1j
q6ClQ62pl9XThH4Tfb/LonC26cpBPUNmAAzt+tI1F4zg0fc0gMuVrxP1IYBlaxFF
wImhFMh0eDLAd4IIYJ7y7Os2G4sJgVs3k7jpfqOKu14wVOOzo6OSaX4ipFTVlIHK
qr2XT/APoDkDQZzQuehEXu19NX7Y/TP9ksYYhxGtbD3cjlhXcbG0sdZupeWagUAl
No1DWindtU55QDAJDftcPPNL86l1EJhOKZUF3iVt3Bg1fd3m8SWNnkmaal8m6PaU
Hqolyr0AjJLan7lnDDAXL8RPymhORgKSjI730b/GcAyNytv+Jpkj/fnKrwkP8eyb
w8ER41cyIArKxKFc6eomsnTXNsd5qEuegqxUciYblz5UoFDoidEDVEJMChyrv0DF
wJW/Gcb8jMVas4JaEpcuto9z7U2odsohSLqq8s1NN++SOhAfhVOU1VG3Y/5usqCN
Dswe/Ad37cp6jFOcvwcJ1xQ9gVN/TfQeThE4qEKq/iX+5foPmqc8sEo2ynuLl9WA
4rulXvsTCATMn/qIBcHuRMv9KktwGHGzXeCUNdMnE/ZbKaL8a+6TstzD4/KvB8UC
D5onx+n/DKixABoPkJBTzBqxvbjnnS+1EjGBpIkKmr7u5Kopcz8ODsmU3G+dZNjv
4h0RUB8eZqMNqZucAzIULeUSd8nk6GQtA0Rp/Kj+jw5UKxf/tz9nyzsOUdei2Kit
3edgX+Xdl86kYDZiGBnDTAEPaEY2TxLJ53bXiulVVo+hMwIvoDL4uFxd9Oagsxq5
W26U+ScUQdNzLx4JAnn8q9qn74Y2/YiSeg7WOIyg8BATLnu+DyUhAGb2ehww79yj
P3PntNx3QPMX1yoiU4NfF2nz+l2tAijMucAeQkDwXgvFyZWPvwVn1pHvAKQU8Cdp
8+7cOtI/0/dlT28rBkFNqsV04iL8C8aCy+rv/YeDKp3TfrUT7R/ahLpgRCKdHgVp
edMKJmbPI7aM0L60Y8sQYTR+0GHwgkWQfGL2XWQh2JsKNIwFYuAtbCuf/rD5736p
qQwWWkkf4uc2AF0PCHlvPHpCQ4Dy2Mpq6/WjH1ykLILwLGG+AKG81FE6d1mSCaIE
3qc9V5XH4x+fwDY6eT4uEr2GUo871EUA+TEFCJ1SOogA2a5LHd8P/hFfa7n1X6TL
vKJfx5i2kgCkizPYZlOtRnyBb4Gg+SubOdOHPK5Ybtmo5mZSAN/Bik7M2079hXmQ
2VVFEe9m634ZooxMrxlNqEmAM9IhaVTO+p0GpV8E46XSc7HZSXiKsaJr41cpRlHg
IFQiJAoV90sHvqNpVEwYaB9CCA2l0iKELBmFjIrU4jp8H1UtCctZLOmd5dSwz21l
630a/ZlLmhTVr+WYw12SnDuuo4ETigT7ObiQTE8yYxclL//59FnG3Zg3Tbm82k77
RoEt1m+scHwWZ+LkXq3WJiVXGFXwadj94pzIZYACb5yaAJIsAwdEkgdlB9EDttcR
VAMP/qBRZj9uyNa695Ra+OaWozgKWox+pT4CqmDxxMix/tkPKu46cX3kTxreWiEH
+M9WkobaInR095a0mMfN7Ltc6M/ZK6VfdcJvP79FnVZk+i83Gm0OaEqU5pGEE+Uw
1fxBHlgbJ/tOB/0JjdUwlSYV6+FW8TD9AtcuvJMZA9KaBMtCSdGz+IcGbG4CCt+G
ZzPRrmMNUptBvUl8As3GD3spSd2cpBzEGkdMakNwVnZYmKx230uYLetxLsL84A1E
IwBqQp6rDmBYGVQ9nd+baMSSlHnB38PG/wpgyXOX/3VPbhLzB75jxSTQ8bGOIbCm
yzSagmlJQ277C8hk0860mh/L9y4MwuHugeKCoPS8dROZjpgf1fhMywX/KP12kZmv
8XAMXSLcjkpgf5B7RKnI4+j7ztczy+gQQPHyQ158qK5JfXZP/TP3tcunkOOLWXQ8
+4I4D6K10mi8cKM1oI2X9QF8aOWszsUy2kv0QtPYoTfDoSdah01sBUo+hWwrjN7M
nq/jY8gp3r3rbjYFuV+gxtYfQJ6cOThmYp5REFAjM/pFE/lTTa1JwDp0uRF83oeG
pee9f8FmA9gJwRG4CFYZ+Uij4Xdarhv48XQ72YjhQTiq84FwZa5zaqB7N/QdTH3m
lxnGnxfXgjs3Lt0xA9sRwb8w7y5WutyjFJ2Rj1k1jv3WqIMZOrJm1Fx//2EJqLjv
QX/DsO9O9BJ3FDvuEm7t8C/QqiLY56S4c5W/p5/lGS4enZjdDkNP+bHaZTQV8SoR
fr3QZwzYoqsj4kYN0NPOtuz/cl8yw9MLZkcSQ3nEKFewgXjEKyvD56UtjNWgaRKE
LVS3+CMXWCcmXcf61F5C4CBpw2HNrooucjSrV3YpddleiAgkrKcsZcFGgW2Lp/qS
xrrBX0g8Bsc8BWleqXxl/wkb1b6nQXyzTssy2x7d+D44LddsPsKw8XcPP7Bh6KTs
PRWE4/WBYehrwb5zaS9EJek57sAJO8M28pC5ByscK58rtch73MsXrx62BRJMrR9G
w43QjdVnUZAgbTlNG9WX+Bnyx3kSjiLsgW6MIGlfYdR05PtZ9HHKUt0wWjs6vDMe
x3O0PkA+HfEdskRBccUSpTkUvRtVrR+5Cb96YyJs65BFzXV5JGNUx59ir8XRQ5Au
0Jt2pPgo6ZDVM0s8F3RjcFtH8ngRNNU5rR2VqEIhzk5+BpWEiUIeqRiOIw9C5Rpz
grdSesfRxzMlTQOQV8G0W3FrjHL2uamQjvscDrhbsL9iR0VDNqXnKRj1WivVOPdW
TF8Ypy0gzlLn6G2jzFNXrXvKEcoawySXdG/0z7lAxcZgOciSHXl2JDA8Bt1IBA/R
23NhXvYOEM6Ivzf4PeIat6iCFqX7bck+z4yepjd/SlIUoWcOrsmA13DeEuyKkgB9
0B2BBQ9O9Vo7MI9wJfiej+vdPz3T6fkC7C11f06XOy0wxrl30JmyINePHofGBW2i
WiJ5enyBBt7OwCmJeLUUHKqLDcjqv5gfJczO0loB4CaVap8TGDhUIkKxAi9SsAGN
J8KzutIWvKSUtj/HuwUfta4G6+1mLW6N935OEveE05wqFNjUmGdju/kdo4z8iw40
rt3eIM2XRqQJpuNc+5rxGEFG0GptSOy9b+tgpm4uVJyQvt8Y2LbX17rSkn7W6Ft7
9qdu+XBcSgmMRDmTWtsmEOGN1JJyTl2vO2dEkS3Um74RMQ0Kf7vWymoqD7LvJ5iO
jzEYCxeC+ynoDX+2QbKd7jFoO9ZVa0UIwHkiyue1FEVftDi8uw9PzUY03qsBgkrU
eV7qLkx4hfgEWp3TKBQzC8kb9p2/HdAgfutzXa+9fGyg3hJ9Pha/cniCGK0/6Tud
w18IWUYY9bKVVnZ7ix/HE6uN+pmGX0DWNhZWZ5xx2xshyXwzhRL1zMYaLhNJWVKS
E+kaxQSWXIBnSwuOWZhO8N9H2PqpdfcwikioB9flq8c3H3MVdDkruhfwmyk5zEPN
hTqyMGakD4MJsl6XjtpaEwBmpa1xUnoBtEJQw1HiiyYMC4nSxv8Wx0pPfEmUCqlJ
s+mi2g3nTdLnHgFI7lEuE82Qh+camNiZOY66LMkKogGwS46XQVWkQBL41eHggP7S
jIeQ7S/uvxQDmCJAR+5GPUkTZ3TR1w9zvG9aR3gEHDvB5APnsn0qzbEgtHuc0de7
/r/tbHFxnPrnqoMgIT8ekHge1OltF/r7VjWgQNnaxDxqhW/1v2n3rDTguNtDp8AO
RgSKYhuWRMrs1KwXr9QGnzm6qQ39s3X1TIbjZXKBLd9kweKKg/iIJ6nB0DHlWCxc
9r9I4QBQpvk/iqbYMXXyEMm58+iRhxyfILKLCfyJeUa8UuY3+40As7Zc9yq6uKtC
Hbs1ExLthQ6rFt/fYjJyxyu7yiXqMgnGdZ5pyjdmIRRaCxU79UMs1cV9QN5jbiXD
FWnF6Rd2nY7zGT/fPYcitOFeYH0YgdOgByeFhbXUcd6C0l7b/G1LkFc7Zt6XJkBp
ZikgIgkY7ApZxlE3IkVBcxyQlVot2ojf7GCd2Q62gibh7MBmLNs0GYmJmawdvvCG
/oVwfka/P2nZCy8RxLhC3oMQ6HiKefe/VltahqfjagJAJ8X0+4HAqEQQvwLFgAbM
i0hqkjIeD6KO9WNcCqDVDWfdtbush7LR6fwKgHepr73NWIV4hs3NGWR2D/Ru9BZc
CL6HKcp9QvNrNNlZYqxHGTAimaUeKaeclOzf3D5df5X2xr/EFRfZe2L7ASYTKJdN
x91Y9iDSmQckAqjwyV2HLmZEFDAZf+2zkztNaGDbz7taIDKhu1oHQmySB0et1qop
ljbF6OJmmYDn7RVd1XtxqQIeVrIqThnTJMAlx0rwsPkorqLR4239U8w39RNXwcuB
x3mZBL97wshugVnSziYwCasAQJwez78qWfXpitjcmhn26P1uAnLOTuyI62A/+acP
bbJM5VGeHtN6Iu3wgc2N1nBZPhue9wwvH2xt+ZPVmrXuEiHCxg5QrWSr3F87gPeK
Yb52LlGMnn2dfDO2Komykl+5gokGd1zR+FGDmKbcLYNnExLqFW2Q6+aJv4JFthn7
ySZk+cB93cKn8knPg7jBNOu/TtIMq8ZUKNrFR71KTJgIFAIfWX43g+rJo4pWBaL8
UTFseRFG289okolzJdSJbrMfczuJ/swUGaM55dJV34U7qQcWBhOH3DnveEU37sSq
8HHiWoTJqUKCzgGrkIf2ERlxq9bRhuOGWaDwnjZDzdF4bEzaMukEltLIgNKE6WGS
vmJMVPnF5UjwpEGIqFcm5twJzDlBKSmne4K+X+ooRlWhnhKkF1gau/xoaLzGr12h
aM1s6IcsiP8DYkp4BQgHBqiFG8w1BI49jgtcQxQYvMRffNfbINDytnwwJ5hISPQw
l3kog7PzlU0/3ignZjignd9AvomVjQfLMKIW4JUn3C+MhjJmqRgU19pzh4zyPtyM
mN7na7WXeA15BWvny9jxgSK55BwVPqhcesz4lYSEAwx+yUtT7pNbKhfB9mZxu/Xn
eSC7n9PLpVZpNw0E1gyezPiwhTfFOUpHXPfQDFhHcIeb10jqe31pZ6RgHvnbZukp
LIIq10rovGCw5pBkZ9e4r+Z7ZURtnXBaMqZbdGf3MLD7b6AhtKr97PnsQpLDn0Ex
LthnqGsbVS/sKZwrMDFqkoWaONUQP6XpkApSGsMiHF39mUnY/o+xFjd2y4UMdIEK
44uFVjhlowiitHPA0VbK16OAB/74X+duBcxhKshxZusdBwk7+pIxtvCHkkYGUx5k
krJk7MtCeBgYUhETJuu3B5wW8wRAxqE2deXXDw1MuWIEFk1LHA9ussNlHp9rHXLh
0orZPSnEhKETaFvhUMIDpeTyP6/zCKu3jDYg9IFbr8dWWRU5FvCA/QovHKxkr1zp
8GOjY5zokB7JBng/JaoejuaTyxKN63TdzbCEfhJVag0utNz1qDHqojuT7MXxzEgO
IEYTHJfndfK+4Bu5u9f9v7G9ztrbHoeJSemTgMhjoGq0ozzWxiZW9d06PJ+zL0Xb
1NJY9+MwQ6N09c5gYh6eCfakcaA491OQErL4sQA9OKDz7ZwQGEmANw9heRcShNcq
WxuuBYpxfooPNAvXjNG4nD3oWmePwPrULTr534jC+A+aK1LjJBKfE49hQhLT/m7c
qY/M5SsqHrH8H7eAgXn8g9vsjnZqIxuwwp04cjnum0y0t0HNtPaivJC7BsRGf2FL
XCZp2upO6CpyNjrZdyPgZfFMdrobOMwoDaJu4WB3HFBrMwHekRS6FLZ22QXlZwyP
knTvRUyLXNaBOd38xmfZw0yjgP+88S6G2zxdn8ChUx89R2qavk5FylKFHk3F8SCC
TmewkdmTDWM0T9EZyyrSh99MjY9cxiMZGWvc2ZyPFxSuA/gPwMiJu5iDHAaBmYzz
LPDZB4/DsEiXvcwzVzoW1dU6ZgUfjTEr7cMKJnjlC0GzEtpZDrQJYG4HfhoY4Zy4
p74ONCbaJO7YTldvCt7oWNfNZwK9MjwtivszWMCtULj8tHDYN+XkmQ8w1gMB3bnS
o8+hYKuFie5ZHqKlIPRD75IlxuwDGCbGHSgjhRbglfuL7nPNe+geGE9wP96P/+NZ
0bzkbPx5tUBBJFYxOFhTb+qFSOrFHEzSJ+DVyS4TxsIGMP50WBBVH79bRlgvEaeS
y0zM0AUkkhxU2fAyApMBOTTdEPBtHq8g1CFGl1BYKIT68Kk6vt+GMPveZzdODkTE
sLvsckXz5IWzoj7qiWlcZOipz6AMViDfdx70vjzOFycyndHYj6Fod9bKe0WZdIwl
JddkAwIMDUlHCJlZwbeeOW6r9iQKepY1l6wZM/vhRGUsGzSlCrcd/S+VjrFW7a+1
EH5SCMA+qEwCkrcxGM3HWajzqXLt9/7cKnyZyb/0slGA5jQDUa391OVTuyg21PvO
Y7QzSyLdGqRfLlj46NmAA9BbGzubIvWlKkUFo1FiZ9eajdVjcOKBU7xbF0lkSgL3
yRelLhnE7QP91r+yVkW50SYHPERyACdR5VfuSKvpEQkRFlB8vg92BN2u/ikZ9Syg
dOAwqMp3KyeQtW8ONtr9Eix8nZ+wieZLKIEeEzuAxfSFX5yaU4n4uGNjTvGRd6T5
vT0qhpL1ySAMGJ4X9DlqNb8pKSytohxBoySXgRPiPG2tUR7CzOja9fBjHEulIFPK
1ShpdoHgIIU0/+yI248JSjUa5/HyVjI/LBIlsHoICGiLaZ+pr0Ar2uZf5MJ7/Fy3
rCejZy74SgdbdGdFcUU3AZLR5+L3r4JsnVEnedDkBd4VIK73D3dCG2qMEJrRA4UW
5sFv8P2NamCCIxEGvwMYXqFHb/r0O0+mczqUgsLS45EkRpHcbwxxk600d1kyae5q
+m3ZpqDKC2RYYbu1OkLJINz7fR0ZrSwkJAkseva3jAajbnmzibL/DoApUXdpq9sl
7q6iH0coyYEumFddy+v0QANiYfyQVGhc0fXCe+vcG9Mqr+yzS26yplqcEpavT+Gg
ldpTkWKpliuPy/Q8/EquptEg2V9Rv6sqBwD0G8d/r1Z1vcf0YsBfJ2VFrb4sD2pB
8nK1QKL3DtysDWMsZdLQohFvrwh/bQsRUlmiQgDqTtMPMGO4MEPelXtJpNs1P101
7+U3VsU+yihHjtCUtMAvnNjr8ueJZrDABNyyh6imeOL/55DOQQz2pJPVkUCicSG1
PwVqDenCHqe8sIT8QwfDoI66JMBHFuX3kceZRWPgVuIrgf2S0+0iVYdDhnCSydAH
CUo3o75NYLBbKiXc78kh62BGl9uCPyLn4pH1DuOqxU8BafHNeGv6Z4Q7Fbo8+4wc
GtJxi1QGkHpn5gjOaoVR3ku1E+J5HFUb1AvmN12rHYvfQqodP1QIKEoInWLdroU8
DvZs+VmlPjFrgwXkYo8BA7DhZRSrLwUrOBTqg4xdF4NjQNyxQxfoetjuu7nn+3zF
XeQqSXC83LDlFOeLGqLtn4hQVQJS/c+vyFKdxuAxiuDbI8MDvhgAbbT9Z8XR3eJ6
mu/sZxosYaTNNEE+9Mq+7jmokFDLHi4FO/3afwxQ7/4GcwYGgZRfY6l8XuIlUu7s
YClGIIfQPSWA3iS8jtATQP8ePppwrgj/Wt14tiwq+SKR6XFTaCAqyrot0/uUP4dm
D9cLMI52vjWNzLGWH042/EOPekxqgG3gPmweWognCsgvqtNAfHa42ZH61luGowHE
p5xwuFw1wcs8TnZgy7ScIS1xc7i1ZWaj+7LF+Hmxz3aEEiD6cmWh9ooMZ+LPLI0s
6lEtlJEAGFtSLLXZUGO6JoDjMXCH7r3vpCLgfJpqBRTetLrki0dCOB3MnMmlZCzW
IXSaEY0drDD+dmIEJGO75NftCrwmz/3cnyNNUIIdZypfIcXZvUVCLwMEG45FFLIN
UBB90UXc9eeBJTm9Ccav6zxFLjBi9X0+g42Ncr1y5PaYKhK3Mr7ivAeGI5tVkR16
bfI/GojTmFyvtq8Ba9+sDKY7WpA/B9sommrzAR8Q2H/YDmVW+74Oz+Na/bkurWJw
UG+DMfZD2tSjx3Dg9si2U+DXo3YRhvM3IirIb2a0TaX4b217ZEDJvMFhEgm8izWB
YNBGlACp1XQ7nv2GgizMvWC+As0QVPLdOTASLma4KXd+A/3ebSirj19caQOwiMFB
aSaTC6dx/rxr6SkcKRGMlvQwdKMzDAHbmOCX20otnh1V+oNrPb15SBA/smSF/oHr
56+ft/kFoKSI08UyeAFvIeZEU76BVtM7OELyUQBGPpErxqjOMDv9p8Bu0iGlZ6yz
8Dl6LbKIU7ZZNEFF1hov7gq/URohomaFHsE+7b9jA853HYp+B7/dyGr2cniJN6hl
dAnu34cFp0JzyXZ9HlAKmt9ZOiFXHZqQgE4U40+Xmm73LW/35G3ejT4zPdXJi2ns
6qKKR8CeYaIW/qqZQQxIaSNFMBUJowpYadZZSrSDYFDkIS6++NTkBxBUpqOCQSCs
7rstNqWkKzPcXHX3RqD1/uUEOrtI2MZvRSgJ+VNTOtmJfuuU1SWnkJf8D7rj3G0U
Qoytz7XpGDPmUMIrGg5y/LYWHc7Ou1OwM5dxFLmWps5dbySSZdECGdjfGMtIN7P8
MQJNcrIZ24zB4g4a3AswX2muPEZwCWILluQq4oceBe6SsZ/74qUV3yCtJTo594IJ
bwua8JiykgoyLlAP/RWKrDQVxqVwIQRiJO/6/vSY41CkS7SkoYcq+Ltb4FhhaCUe
lVU7oED56QeSp2VgZPcVZezEkveAoYijseMnb+eWnw+VyTAO9aE0TMXJ7IjodCbe
KZsn+/f+DbVMr85ffmyG/U0bfbkbwXVXOnlFwq7eIiMG3hvGThNQBmmssXbsqOkc
s4NtxlRJ4KZ2rE5/OGRGb90LN3FwPb/PPgqkD2reWvNuXv0AxjjeGL5/9Hjdsq/U
nI8bfbJItYE2n5VfGveCkKa/jXlvoOj2wXSUO/YEvcim92+QagKiqDB5Exsshty6
pzw1/GNcp0DHUrHW2zafOLO5E/yZSBZMZiNxHS09/hgvo3yKROHD8vpBLOrpVO2W
KpH56/mJZnwV1ZFolc04xvk0u0ixDS66N9MTmBhB6VvuGfYl80/Y1lN5jImgHR/K
ePGxpmOMH8IpbUyz578Cm7M6G4MLL/hbUocxKWQjuW3tdNIIu7IBGj/EXNT/4tgP
LEE9qAcr4UVbiCsFArP+VNGtb4oRnf8hFOUOmWTNmK8pIQBuwLXc5ZWosPS7cZal
o+qacwEb4lfinwOLXJtXt5UlVwo2kmLc8GoAl0dsZal1REkl3dCTWR3ysDU0yRVq
4EMX+e1S9yWGmVecFTpgZU5fW9z2DYBY8EV3ekdlyxEf9W9U5mjaeg34IkHPQHa8
SFpQFngZuYMP1T+KZfXzhWTh9KPVZpEJXH2/aiePXyHP0gxOzBWC2B8smsmwFPCB
Ar/ou+6U4YJ2D9OfP8TQjMKFzVK4SjtAHnnOfWcxvhGoe7owvTeCYedz44WBhyER
A5hYWe1Dt/Gy8JFjVkpOx9JQseecKePsJjFnSaU/xLk9L0hUdnua9SIT4iGQ1QsP
lt8Lu880nVfgjh5eRVDJwaAR7l2Jsx2uFqxy905R7c0fAq13JclbZwkP6BVY8eIe
p4yPHiOp+WtX09rr+wuEuFYGf1IeyjOLL26LRrGplOwWLEEeXDZvnWNUfEd4UOHg
XfcTyX8NaIVee8xhCcVqLODYvEUtpqg03ST01HOAb25YpXWIve1ZQkTzLyXQ+9gI
LW8Z2D9nM5LZ/lMA8ZNg6mYcfpsMAgElitCrDivjf4a3TQ3wqQuchlmXLJH53Aqu
dLGARVzUMhwNfRyruSMb844yPpLnNGODIYPBMjCdXLItHd7R+eFQlQeFdZ6nY3uc
QpdX6vKpuz/yIShn6TnpZSxBkSqal7xqMaL3N9zHZvaZogaxrB4ATghfz0GmF+Cc
qU7DeJp5zSq9mmAlzq1bamAQyvmmG/g0oVO92E8Mh68BR4rHCxZ7DV/VGd2LzX+N
hPrxQQjF50syJ84ZyiYnXTPvugCl0XL2SqEXRoQwRqTN+rhQO/L0LhVj4UpPQ5zp
FjN08vtM26dYhVtb46acXGjcpC9jzZEqbq1fsxm7V2mfNnfzFxqWvDyvYbowYLAs
ImX2V38hZNWG12mz/6/HJJt8j1jQjzsyXj11sddoKrNX9O0v4LvHZqDziCKrWzRr
BwynvvVAfntLTCQh+uDoChx89WDSRHYm7NYfaDHTVEsFzhC9DaUWHpoS6yyEYkwx
/67BicSmYkfNG5J4nblwzcxGrzRFsxQrM4bhlNhAN21464cwzmWxT7Bgpe1a4u0M
Sn9/tve+jp6EzS8DCApEHOS20OpIaHRb/14hgikcPiHDNWh98DHUoGb3jYqEjnxG
tIrdax/1eAzU4kapBc7lf+Ca2ef9yNWFudFU0oEgiKvUats7mhqaUPGS5BtIQNSt
o281xdzbM73z+tMUjoF6aBhoRjX9//zsAHBZH21hAmx4x3VaYUP8sz/1zIPoPaar
ABCgCM+8aYEsDwJ79ARa556dsIV5DxCRTcEeyC+njF4w4rh0flXZU+UPah33i/c9
PhNIdlFP9OGHcAGUezfGb7l3BFX+E92P7wbxgduBFdEHa6x1CK8wI4Jfu4Wf+8wj
4cNjtnp9MxuRK6zKTyn/NEXVnvZQD81P7KMkZNaQp7k4HEsSuFcSiEm3Cp0E1GkN
gGOqq5P14qD2M6TM6PF+o8SGou/Z0ppwZyVZrgYktF/aQbdrt7w9HcwqYLpz141N
YTvDXtt1ZJpgcz9SddFL3B0bZ0XbdVzcS8vjqX0ig+KNl5mwKBXu3e+tQVEhDMz6
0ozlp1T6V2t3Kk5cpRvPijni3Dvz9dVMowp10y90d1W/bnLqfl+tKkGZf32zMZRt
7niCHv7BkozfC0yXtoOXi6LbCR/bs1hqZgKeDnqExSY7lXU5E6PHeq2Ho1wDWJOo
zBAuzy3U00QnmdEyY5ya8Nxg5cdKI+qrBMJfs/FpcqpJA/saRMJDW8h8hUmAC7zI
ny21kOJM78Blrs1nbHbTyh54vuqtBzB8vUI4cbjOSgr1T1TOyjEkZHcEAW1qSlCT
kelM2fv44NpKMXQfgq74ArY3mhIIhJ9ngvp4g3FeXKsR3UTgLgD5hatEzHXya/+l
xAsFtFEuDuad0PdeYmN9lRAdctSfre1Hwx4+Y8m2iVOHHj2XGtiPPK06AYsxbjXl
oJ4iscSnFETeh5krhnHETln2nxUj3JhJFFv4Ri3g5wQfCQe5szWzJpHjyFQGwa/b
iHW4F9cbykDFey8zlnqST2ePIH1dyXcC7Yl5agXNe+Hmr9N5L02ECeePINhfIQnO
4PUySjEnEWFH+78Agv2SeaNi+QnX/ovxnIEEaDaEWIJUfXgMd9IXwWV1rNII9QGr
T3yA/mkYGzPTnUCiTbsXMSxmK9+OTZtZAEwvkI5a8P6x5J7c34q/zeGaJ0naBDZC
3tjzUQa3nj26/O/EY1Pgr/WBMjlDTjUYuoGVK3DtySkr8YFA3XSbwJzImsDFtXcw
XPmTATxllVUUsChyCxCYhI/ry82gblKLEBzprL7MhsbxET3m7cwvjZr0drhSxzAG
eUSH63zmcojmi3DBLA5ZSAr/YprbBlQwZFCwOE+jwISgJQK3nhkZftgBSg7YgpjA
jERafja7UTsBVb7rmwXp/xdYVJZkvbpqnq+BIiYiwhfoRLCVv36DocbvNjie5btm
4bDrb9fP16PY4n0AFUWh0odjthmbgJa0QlC3Jdt28dj707lvGlyQihmO8KnAYtOf
rnBJP8qczqFmcxwJbRa7eX8QsK5nme2y0uE+vtb8AmEuuEcxuU5Xsy7/pGXf/XbC
kbFrY8sI/IX0RUx70IzfKnNhueYjlTgNhYGC2q3VnLRYI7JEMcPiDULskXSHH/xl
O4bPZxjAUDxy3f7BFlSaIOW/HJBsnQldJ6iIfiTSZAE0y3+ggGvePr2H146+xoFr
mZAo9r9RXJKnpJtRp8/xF8V+sAov8q1KdwX9L4dK+uICIPgEZH5DW7+eESAN9z/k
5KxCWalpmB3Catjn16nudwBwwOdjq984lPQ4pCLaN6575VTN2RoH4gep+EyW8kHp
FKV5zHM/Ofu3tiS1eEooEpxXdDF5dExlY6llLTH87lQA5nCXWauqH2jxRuRbXs2r
sTl4Ki64XnEShW59bZikbKc4oTcfWzWEPT3F2KemFaWjY+Bf4mgjJKUutsESI7eT
hhCc1BcpALwlAUsZB8pO5HfHW81rN4cJ3ukALAwb7v0PauWqaoe6PmbDY5BzpJ+p
Q/caqijkub6k4eSCItvtqn6sDTHFMc7w8WSGlNV23GB0xRga1LpISbYDAKvFnf/T
JPLt9guWkREaw5xxZ7k/1W+5HHQsfVn6sq3Bm0e4kTrPWz3ePmbdK6C5QEFFdsPS
y5vGfVVlVl6UCSx0BKSjO9gOJYEk6EjJFAQjr/7kyOJOuTJ5cTGwWgTzWR0CYzyY
rCFJ5iVTkyC0z8sBkcjqTPw5E9QjHqrbnLb45qY3TujZ2tlDL9SVNxl5JR3HCFCw
6lNDTnVl6tZ8hCrIuAxHDzclbt/DQpAVw+brmat3v/b6M/RACh5CaX5omm1urC19
tK3I3zfohiU7OgXl/v4gPLKNYwrMOLQNQOt5jHAJxhuHaV2IsvO6xeYfDQCRgYWv
F3fd9ga/V5/q55pfw14mvFKMkiAA3t5BPYUWVFLe7hdDN+HDj/sganqY7HMrraY7
a6Vd0/hpZrDyu/vID1K7GJBOyynLGL8c+P5WU95WJhqb0DX9wMXJdjo03WJ8Ooli
0RhhPrGMwzUKbXHrXnY39ryYHiH1AltbUihznCbunjYbmnBOkx1CZr65j3q/mfCf
opbSb8cLhlmd0wfXbgV4cmOEQexKUCcg75yGXQDCzzgbgseuIoBRSIzEs8Aq0JEW
frBOwvCJ3VeQ/doccBDriyVbNljrYaqIdPs3053pXrEletJ5zCg4SbW1CwKRGi3I
SeOKxWjaJ5v88UdVzgEQ0vAh8m5/jdm3gqmRGLVHzjABaxy7j439LuAeMLg9o7zc
/cT/KhPGqoa5qr4VwmMLsDMaw05aDzzOTjG5dHLgPqsCH5mMKdCP4dhXz3oEu3KB
z6IsmEbczHzGQKe89e8rTBpKBVMJe/1YwuUok2Fp9QY9XY9nN8XSCGEmtJKNYPON
YIHnvJgNQAYsRIhzkkqO1nQLjh4WBqh3RAvfUeWu+NG477rKIt6GrasIyNXtQA8j
O6PO9qxuxrju/zdCvV2LzIHAQU7r7TFG2Z1dWNJ4NyiZefW1ghW3eHLwFwIPVi7x
pP9acLRI5BkbYFE/vJsBhQG4P8OqX1bk8lwb87kpVMl4rExyqPK+gNaF7vCKO9Q4
2MUSo7ZW3DSXr6PDBHUsFUV6WmvyE3nmY1eHu0Zl5Yw7n0xikqoh2fa9Zayk7nJq
JYPwm/ETlEO21h0XSicz4seQn6RpuI096iIycF0imvMmfRTqwjrYA/uKkt3674oH
+yrSYOnT5Ll9suTj5UFV4Yla5JPHBipu3V/k448ahthmme9flnZW2tR8GGkdsqCI
9xzFFBntJV5lNSdAMjAAw360adtAzQEX+YrcjlIbjGNtpC6dv9xcodY+r4Poaquy
SLQsDc70KoUnFhjf9+oOKiHtIHdyRJfBbyTB84PPp2bwp/fOn1wn7gQKmC8/mIYR
xwdHvoITvViZqdwgu+AbRNQEHcLdPZzQnrraQ9cvWh74jJLghkyofI3TUI4wCI3F
K2WmDY/PQ6Jj/BKQIUt0jy0axdYQRJxBxAPyU/vFh+aQm7C48+GAbMYoaiccH33b
RCyWDBh0BYwtDGWQRwFHyc/kEyywyNJmTAMfQZKWuKtoc49kze6n/yV5B1C2qDz/
SRZoDDSgChOktSwm9IfefKorFGp1CeE9HlEIqQAVof47JYRI5tbOab4xrDOF3gvk
v+lNFVnDPmqnAWm+lyIigw+UpGUPaPAyux0UVI/Pif/Zi+75IDks3EeTMZYmr5P3
mfpvCUyf4R5dFWMdWsV3ImVvlKPRT9Qn80rzAMvmFkURgG5FN5ISXz5KHflpHKNV
EuS8BOh4AQySh+fZ+oRvICDMHFm61nQbAeaXestA6fIhks2NAM6fpMWcDvFuIk8n
sAGySj95N2C3imylUkTahTjuqgVXG/xbQiRIYa2WKruAVKO9tW6NksxLmOLbRY0y
P8+DNerFdGUdRHqjCmlK4mDIluVodsgB8U8LqihHZ6Y77iZd62DbzaRwBzNHtU/o
YyzMUTcRugYouQ5TO4Io2/oPUdpQWYToIWanfiB/eU1o6GG9JOqncfOYlbbdUc9L
DCNSYBlCbeiMZGM+on5BB+cj7JZeYeUkxcMGpmCorfRSSyQloDmsdyOhpwjkvM84
sBBE8RWBJSx/YltF1SiT04/ElOUhBFg9zZYJLSPT6YafCUIQH5++h/gns6BGFrVv
XYwepiWm/sepUwlFJdy6OatPJMguXYgmm5mfZOoAkVlchIqH3PYJCAVV5M4VsS7Z
gN8tS4UKcH46CCFiS/Bmc67f9oBQA0/Eo498mhhISh4bSouDJGXCZl6kzB1fvtXE
Qi3mc9F+9k05Yja5ODwVZzE9Nt6aj0vgzwpXUbT3LK7J0/KRuR4db5l9q9YC4s13
QysjqXSAMnKWdd+cN7lVVoj2Od8tkyMr8DDyt/tJzMzn9CJXNbpcl1Bcme6sbwkO
sZhJK0gr7qL9atM6R7k8boZWlfhKaHPiHol/oDh7ujsMO9F+7vXr32gnRa24fuEp
TA73ulM5vTEqjiw1ODUYbQoy5lZiz7BEXVQ0l+AbOtKmj9Tas8mDRk+JZWDLqCk8
lLQrAkMFWtIr6YwElJd9yR+JdW16zuRCC8pNaT5WjeQ41eaJGSrh0ZPN5guNEhnc
7jfFDAGkU33T/9ZAWrwoFMP26RMTmOXof7orn9RFp95HKLzHtF8qYp7q1HTNG5Z/
Rgs3soVkPtSNuO2iRmTDOwZxKzGfvfh5AqcquVa3DqbFyhF9mzGqqPf4quujFkvp
euuXlFeDnRG3BC1DK6e7rLycjs9rugRH8Tu1BAXkLDdkILypyO2fmm23ji1+fnET
QeZO/+otm6puStbKs8/9HpB7Shj03HR3bs1AVOhy7Ko5hJN+E1dtYBFDzZZtMmFy
5YbQ8ozwT1de9XELcJvPcTSYPk716KwYQxh94rdFY7D5MB9rF0qs4NefLHUGUk4O
yGILXqyfl5bOYAwTypN/2HDhz79QpRQd6f4AZ9CQYvrOvt75PtPogUNEyMQ5+Bjl
f2/HXmEuFz5mTLCvEy8nxzFjO9XTU2vF8se/fQ1YOEpxnMPx+z+3HT3i0EKe0fkP
MU0yxgZ0knlFKFDCAc0I+ys47fyGQKAyjqUTZRBM3dbKies3KMSra7AiFFTVmsuW
ovCW1o7ukGYadBevhgv3ZwSFz3aq2FoSMOVi7zp1l0ZT97kTcjyk+WCKeLhSYz+W
4NJaSV1psyhLN+p76WE5Jq0emsZG2bXNBJWlUYWFcKxoDj7qh1eFqcotVJAoCXI+
imRu/Ljh1X6ydx6A/xb0cfnjb0C2pxwSULrnSGQQIGyjCD+cuhbE0eruDsYmW9iW
wGnrjIiOGFlsK6FNQOm0ogd6d5kxNhjydprKmisXook3YXXReLxnPWxW5CYtS4od
O+EPYEqOE15fZG1dqS7QCmvOECuOZp9biwFNUWCytuMWhnj7hk4q0WeXbASY3EoX
B1i2iGZFsA0hzeau/Krt1n+HL2I0liKUNRHCEyDmDjkxIwOq0HmWGzsSXtjPg1uO
OzovzymGDgp0WXsqkMmPDPblViczJjODbpedHIKmiiasG7pKPsPi8R5PQV1ThjUO
hI0jXkZe8RceycepD8iH0OynpkTwUt6n40fsZXxIDwEZgYgEfBPEq0GkjoqIgMM4
YL+0LlSlqnK4fjmT39W6Eek8/N3pBseH2H0YVhFV/hXcYNLsAA4PO4/dB7aXl+X/
OZSv2OXLJDlYerIo6uHBfkqB6MSnAraswWtVnJHkeE6G44o0tp18hRfocBdsDV20
azKAf0AqeKyeLMLoDC28x+Lyt9/XftcdipO0InC8tIV2ZNHuoh6wpg8DWWsJa7wn
bq9JLX6n0q9HGUzw+a0Z01tfwFOT+JPZAgxoOxxe3zsUOvIZ3m9xgD31+6PP7b8m
esklPvM19ETtqnaTMoIma7wNOEOb3MPGrkaZkXyrl+5688BXcEOmlwziDDRz+yUE
jHwpQa/1ex0ZVyZQLyFWD/EsjuxqmOFhGByOe3QOgdXkeOoQG/xEVW4x7H4mSc1g
qh+6feM+a1YsD3B7/5LzgcBgjZgjWyiGfvLmgE1Ms0Jfc2CRrLKvnlqa9ZRPrfnA
+X9yOGqkTcTahMF8KDyUf234yjmh+Nm9jAyWzjMs/j4FynaJ7o1CDvjWx4JtOq4N
LJz7tai5+hEArdUjgcY21n0vPxrH1avmv/v6GNv9cB+dWVH0GurrycA952jECAXJ
UIBWD01gakItPogU6iqPgYKgDEmiB4TNIadkzGYtasVqZWLjHb9ZJTf24ITm4teu
PORrunBdNkrlbHfVusHb7wuOzsRc9O22sLXEH7OsgEJ6RNStV0WkZ1qfsw9yqJ2Y
VSbJMAFTYG9BgEXvzLaCIyh5+WjEbnRxRU8DaWHRbWoEXIeOGTkHq65loCZ+1ioX
NLY6bSI8Toi1Ig1YSMBBmaH1KWYCEPyaZ/9QqchqpNMM+uvNHhdIw2862Vdgz4vt
Nb3rFGEcMCGS+weBA3MOyXTOb9yusMf6r5Y3XrT0XnQc6QiyPeq+h2SN/lrqgMEg
0MvAYqVndXNRrbCwixxgVjbkKNp4sK+DmCotgrtnu3F9oLrK9OfSqywlvIK5qm3s
Hmsb2n7g74pmNGoddD3mICiaILxIrVGdo0qlVcn/R0UeK48Qet7t3d/MKLFCNG4E
TojJmJNGenyE51QGqjW6pHOoPVbFeMlo6mDgVjsOh2ay6R1FkFlhLHKOEZnkDuxe
xFiVymos7kNsOspUKAp7c/g+MDhNhNoCX29TuYlmgvZ7sZvWwRqdyXU10TiYT+x9
4jY8CxNcYgBDWnXl8HzTKJVn0USs3U5vTW7TsgUI3vEbjGn/oJ+dWtP1RZn9AF1M
PPm3CEs3c0IupMoWGgk/Y7AQUoWOsmXSaHAemvLCMZFFvhIuIOv+WKauBokF6Y43
ZL4ZyFefsR6uWbMN46zcXqCHc/qvqOcwhhlxX+Y95WC5posuJ0TaDWAftn8wpHQK
QUoHtuP3fKguvdlzinlaQ8qDmSnpzavhUSO65lyBu04JY+91N7yG6oUp48oo49Ow
XD3uCYw2kbgcNywdm1189DO2jd0XHgKlI5ko2jIhwYrydBUxVYmqSL8YUEwM7TGY
Z2B9XtxAvx3hco5g2WcDZQ68vRkuhOyLE1sEF3Ye8/HQgXySzs5T3QbhLFYyNqf3
ZvcsawtZlVNxG5FZ6VWdTzHwyhTHR55L/W75RhhoCDZGnc56MJJ1Rf0YNXsCe8sW
mrrsHUy9t+9KDivfZ5MuZ/016bERYS8oQOwH76p5uAVD16HjITKxaB7w0RwyiCk3
A470hw4yasCMpf+HJWcjfW2+zzSa7Ws5N+eaYAOWOQ72TisyCUdWWxfV6SjEl37f
isZCvR1VAgZqWcnB/oW+E1sgvXqyyU7Y+66pdbi1etc+rVr24svm+4Fx7JDH2Lqg
M+TWmHtQ+HIfgDSQUU4aVyjsZyyOtRqLorBCM7zQQ423fk0+5qEeU9J3cb2a+71k
NqJtNz8hVI3WD7P9b+4u4ACdXVmTdBF8/Sm77pInXNpn49mgEJzNN45hnEGGzkUD
ebBwKSRSNg/FP5Nz+FeQlmI9WLMKis36RfIqCSC1nphnSIDPckSBbTw/tzhmfDhi
ES4vZvsFKVNVCm/3Hs5jgHffOMi3zxkF/UDRYO7LQyJOdmFJbt2/3NgMKFyd3GMn
w0UOh1s1f7ENZQNfrjfFTi/ti5GGyVjnGoKJ1nOjmx0+c4nFThB1ckE3iA3Hdkji
ptgLsODx7IeBMak+RXeZkc2dDDNiTsEFL4OaepXZzyviuYiY8cKBLtfWUTKBBYxs
YC0ROmn32fCPZzBTGbXrHUEGVOthTs0oWbXuTkKBxD95Y6Bcy1r+evoDsmYtAG8+
Po5hACyokEnK2mKS3EiTWtm2mkTXTkg/anoVsjDISz7xezc4ztr8Rv7n0V2Lmdhe
+1ywsayKdN9Ld+voNeyhuAejXIXlwDZErDsGIrvWBE5ydtWht+7HRoO3XaWQH8EE
x/s1TUI6/cN6yvvenoleryG8dTqJVkZLTgghtkDtrip21YPwRg0VOeHixIGHcW5T
HZWgFTLkJfGFCAtlR4YdCv97DKDv5ra2NN2iEBTlWeaXcMryNcXYnsW4AANap3yt
UOaLzduMHlsHQd83dRD4CCvaN2402EBDz2IXcD6RLshZMfqKgCGIRTFIBc5mWi88
zLUU17OIca4J5tKnflHuMjZQBHmwJ3dTMNizqJ5hmvoPuOjOFEfXgC9EH/ser2zS
6T6ASLTN+26SDJs51lTjS/c1W8NJZPr28v3Ifhb6zwNLt5e7nooGSKt6EY/Yod8N
fxdCOc9n4ds3L4U7F3UEud3n4BIQTKaMBudK89cwGmqoo9x3nVYmhs6uRlVZAbTS
p0594fWZjpQy/3TEjOVPuNzNRASoYbakDnMqqnxqcrPsQw0wIdGYWdwtcZSVkiRb
FbfLVqSrj141kvN+3jeeHyHoRIWK/ddr3g5q8Gifuj58z7Lo+Tf5AtfLM9DmicIw
1rD2DQxrGSp5qSSjbzV9sGQzHFcRRPZqj2facaz3gpKJoSy41dG7Gmzsp8ZYazjd
hu0zVzNa/GUArSNUFPyQOXcodOybYJsqj9py5vmHL/hRIPcTC3lHqOuNRR376T0y
rWW+DXuaNgAPaiX5sqykmxqZd+WEv+Y7JMUA8Bcba7vvGTJQEKuydO/MGkHD3hon
YayrnI2BuIi2+NprTk4KEqlrAgMHUPdkH/MqYxEIpcwHgmlpaY7/DNXamAgzkpsS
hSTrFTfiaVUfgtAuDhI5xw/oUL6w0j5Il9eNgF/IzxLSJ5X0toJy7JYsINKZjxh8
sjxZnvyXo+hU2vGwQw86YGKdt5OANoAh2pVAhCfk2iQTIGTHihLdpFSCDMbHGJTB
6RMWLALkUBDWy4kuc+8+n2FbZBchgLcCnPMZxiSONzqqwY9DvNCEKGqpstHMkHeE
BRVfUX94zhx6jykPxLFQDJQd1A/Lmpq3mHZCAhCtBb4RzjuSnMQ18STKwQkBo0f2
zgAGMy/vjjnWLAbd/cKNBK4V9N2gILo9xDAQ/Xja31/Ken405DzbTdMKfLN1+98Q
bXzBqwyWS8BD708pfxJQHRIq32GF3GAQsZUY3+iXiwMyAiunn6j5qjfUGAKCRgXc
dyYDnwLu85LkmPikRGgzxv6QPGjz49gB0qy7u72s0xsYxK2kpnr5a8N6lYwHd6Os
/3da4su3s/5Mryy+gq/4NqCcrmmF8TSzfPAVnCx8YrCB0dlnYOhsKC+U9qCTOHUb
9dAxRR1mhzxN13YopBFtxY162omUpZexGfCZg+JXp4zbwM8GBxSyEf7kG9Z+mgEF
hbnGdj0ute04gObog8hm5STAZHCw67oSXvTsuIDgdGFGw+O+QcC1SOU0ESIgX/SC
voef9Dv28xL+TNjzxtbR35cgzpK6OhGC2EGAp3UaO5nC9+6xpjMe9xheLcIw2Q+A
HM5bdXU2x+NhyenbiRY6+y5ERctPj0b1zbr6GHKos0J+3iVh5In8fg5Ee8tEhEXo
r4E4p/HfeQllV4IinehIKK1V7FRkUaHPKDozsDfY0bI7oqAlUvybOJEES7CrolXQ
U6csKYREj6h0VbMZ1hd9/aCpzx6Zq87LL+TT9gBzaTKglwOdLnin1sKG1AiblhBF
QyXrkL7sMdDKe5Ig4fwNUqyjhTF5/ypnFm229lSW9B19eXhqB2iKOFlt2fj4+9Tl
0/S2PNPf17zm01VLZU8V6qo8VQTzHYmeDLK8BJ57Taoiko7WGoZ8WGNKdFVbUCTP
JEA5jUuuMBJ0aDNls6rUW/rFfDRJ7VAJF5at9WYiuC2xB11Efppq03XDZY/gFrK7
2xfcwxk47ObyvltnWSRWcvt3gGy3XwBGHTKyfsmprtMl2FzKBvWpXPJErYeO5QZk
YlJYgb2c5p+L36v8Sawhg5zzxZLpsctDIbaLmaJu/F+8U9uBxBH5iDkLtLLXFDY3
jKKLVZ/okkSGtEmzFJ398DmIo9De0XEbA9POpMp18jCYVv4bExvsq0ys2wX0cRi+
5gti2hhGajjFHSRS+wbz23YzZnwMPAPoeyMPErKyQOPUiscCQTfhlpuMDFxnZMaO
zrCWW/4JnHJPgGFqRyI/TDpjbtQumao1ki6r9I3rXnv9aQkhlkuXrAfJrvrWRFpL
M8++OD6ibBsbS24yfkjkUukiSUSlo0SisdZdf/6nAsOZkTC3sGz61uY8Gz3b4DOT
eUjBoRaTBJSHrgLkRMbu5KIL+YVuBalCu/8u8LUJZnz3For+CFzACjEb6w02r8PQ
1xlVkr7NFWN9VrSR36At++OU14b65rFkCZSLCWGtI065XC/zMU1JEw2h3KF7lMLE
5pr1D13qA1zN6RMnIhjofYA00639PJl4Ea3BmdJrC47p3nSvx/KiDeBDKDurlH9R
UlST6Vb41BUHjtPuVrjO6wrDW/mtotVvBKbZxTOzhhskf+IvQkrBhiQwqLkCzmAB
EAOtQ6+8hK88dHdwe5L4XwxIU7FsL0KF+EbsLFtmpwB8UFRpws2z13yIijuqVo3m
KzdVhfLnWbwleEaXxbzD6mEmedqynH76PpT2sN8kuRyYzP3TFsZEptCre7gbC1u7
HrMI34jzOQ3Zd/H9PjsLcfSLSpuwfKq/rJhubztmvUMFK+hMRhkgP0x+2R2Q63Li
fFy0b/quoa28Kb5JeIZhhEcNjC/NErnpUloKamLldzj1eE94wyJ0v4ugQH7o8cdf
uHNbia0Q36pHjWrEpHRm01STO0HPGN2WTWZjohkIkovqVoLWL1d8IAZAzpZ3lRgY
Qls+vFr3DuKtsnzzd3ls7zyY6A9fwtAg0td09KLK4nOQkHAqadi/mzFvcF1mO++G
tpG2CZdr7T+jC499rNKZ5g7xbUvT0R4LQXKbjV/pSgl86833E6L/jgTC2DR+RsjO
uluUCKnAcZFEUxeGJxxaMe8Om7MJEaiSZgRS8cRwglRVq3yiQyo0z2fEdLaFkBVb
DmRVKQUWpDmI6X6VUBDKDVEUV/OU8A5ij4vsu2UMv8TACIg6pk3zFJj5NtwTyv+K
4UxwDC8ngZrgCBbJx0KCVIg9R+narIINczpRsHDGq/B3xW2K5Fl2q8w8mATW2Nj2
apYrNvIZl2a7vIi0p/fzkVi1HSm7Pav0nHK/GMR2ciBctVQ9b/bFTe3AI2hhuPLb
PNuka2XGtpaTEIdekgwsvIY8vCgLHxpdLplKBcWd+nhLhq3OQKUKbr2bGAPLWu9M
OJ7l9OZHEdQaVQ7NNINC/wo2XCzIUUMlmlIH0F+MUKVjCjT61yxHnnomUaD8YHIA
idtsPGQjYykNT/DEeIXqZSNDMJ6zD8EV9snyuIdRnZAwzGqTRxJyiQTW6dQRP5Xu
ShFOM8fqPbFiA1Kxg7wv6OwAu23MzgCtMCJtBB8nVQIxLCnWEhAUTklzqKRWyF8U
hkDXMBZaus8rmMVfQtucPoUBnJWDkOjBwhT59c8d5r41Jv9DOICFm+v65pNrLcNE
qXFK4ww4LSJCz3aHWG8guAn6kUS/horINBM2svEdxg88lLokeqlknFMBH5Iasy73
WEU0ni/iEGE44Vq8WtmuoBhiV/PJmBUZdv+VKdwQKC54rx+D/o+vKX+VdUm7FbUv
hpTnoVpqDKCWutC8MpemuJogCWZqCqjnZHxT9Kg21/PZXBwOlkOF9Rn1Yfkgp1fR
pSVvFba6bGH60CY//2LS7wJeKwFWJbww2WPl4zNB+bgkSEPJ7Fibn1x2h5r7Jjdl
4E5A5m1CW91LNxja5MT/EdNtrvqxfKtkwYRQsGkoH99Hq+Ww0mSIDRt95UQOo3Aj
m123gfkMj/7PnCpdBdZDFHXtuxDGyHBu/F9itK6P4dRBvTzLZRNkWu0ENrwTa1xF
USCJ8i3YflqWSzjK/pxizc+XLEESAJuIGnF17yhPmlJEZHR9XNQeBetb/99I3TYU
Fs2dKa8pVB4opEKCSAIwHVdqnrTGCXPcaSwWB74wSGK95PggmBBhLucrU4pNq1YH
EvDGVUsXkqx/BdjbQyJToC0cFttn5ZXuQtWxcqVGjMysYJmqIMEPlPy2hpYGhfAk
j88lthhSNQFwCGP8pP72SMu5zMYC1CpUtflhj3V2QFgPe4czOzsSieg0tHiWg4Cd
9ya9LKROsYepTwVYKGjxZ2H0aH/usYYH8ve5YSkjFSdrsowR8pJoV09rYM97pvfe
YTVRxMYOqjzrQzun5dvU0Oj7q6WRDF9euZcnc2arkEIK2FyiMURX/bZBYEvxOWXN
IVfNIY/GODwkouzna1AfOCjPOMF8EbP25anzAHPtRF/EMATIZBCEBqlns+tIJv2i
MkBaS9NikzFIE73HoZMW8Pxl3KJo6GdiSoIElZ8JD31VMnnj8VnyJeq5eLRKG37t
TKAB3Y/aKSjq76lyFrKXnLlltvFvdXiDSONo5OUi9BTDtjAyJTwA810W+/ucj0dk
/mS3irmuBmCjIReo+ndi6w96YHXWnKhMoc2k8wSzOnqqs1sQwsxwJMGC3IRqKhFS
CyFNKGIJYc05GiAbtACOjDhJKw9x8nDxdrapy8gNFOyNORZxYYFRIZsWw4pl30pb
3zrlCyVg1OUqW7On1tvOmISPK/Jusco0K65UFv3cVt135VxHmBna0Ed0GcgT81e7
NadNYQgtw7H8xeHWufHTvv6K6oUOWB0scVbtpj/ikt9F8hQ76TH8qRZsM5jwl364
pIXfF40waTpNKeijlKaGF/dZ+hIkrLKcGadAqDea5FBf204REKOar0ocu4yBN6X+
7/qVS0Q1+jyFRlKNX3UB8dWMVF34uSRT1EMqYhy8ggO5lCN+upEbYq/JlM5s7qpX
XE3QC2l52qAKhuuPM/nwByL5Ja1eurjI9Fq5PlcSoVWBmTE+yi/GWyIS2JPhziCz
P3VoPLMgakDBtb1FBxPwKCZsRMvEyPvkvY+H96ZpYlZLPs0036fQS84YDJPglLq7
wnfA8HONrOL6SitfnLb7Z7+ZwxNqiUQ4Otk04n3xz9s3j1ib417Jtm2PC1FKY5y/
XKD7vZ+yFfwfRbVmO+ZH02dgOHfnHiLqfLheC/9Q6fFP5o+Jma9P3bxLTHbCFvBb
SpwjNO0a5JSCFjCSBtbuOB2NIvjf3hS6JryG6Edn5E+T6OW3jRUOGty45mbLyIyK
EF6XEDx9fe6+LKZtMJoNZnHnP6KrVRUdn8FmB1sQXiv9aO/HHMnNvjbiJqUCgq1V
zQ/+2YyLGfW7BIoMa28zIpNe7fgZyu2ub30i18cMrSK9uDUajk9xLCx1Rw+ZAYyk
S+zJjkLPagEEmofkd1spFGYHQUfKrmADr0AYiHs9NQH+FAk3zuTgL37buoIPlo21
5uFCq+tdW3vtdAn5tLgD0GxSBrejW2qrhohDkdv5epB6SnwM+IuRtFD0UM/dA+2u
yEPXzWmnBtJXCtGB9GXD/+X24Q8wVi9nOKnsPzH6Ra039x7ceC+RuDbaalZfkXKA
6S5OmJrhYg8Eihtda9kkzShB1la5yUdlmh5WBmVNEX2jvOZj3RFZYUNA6nKM73WK
gVAcm1WQeV3P/c/h6OCCyTWQDyq6Skn2xQBLyI/0qMBfXFql+rSGl7Bh7O2J0cIL
dAXqSoor/Fu8j8OIRTN9dIcGb8GO3eo1Rm4xO6AXbA6vYHJMdtYs3FP6RVogMfbV
QGWrtDOPT+HdCrfC1Eip7HQchZS4abPOh5MKJdKcpRk1t8hO0nhR2jvUUZ1KZcvR
ZKHKGd5er7DFKCNEUTTxw+0+F4XxpMK4BKIF/dCVuPnKYX/wb2mOdocW80To/KRQ
3Dj95tayvJLlhRymZB08RrsvOlJoB0JMzml4WHu3pVbcxWUe5JOkmsgAjCttNeSl
yrSXBa6QsD+yVlx8+YsV5Xpf4aLY1eEZY5MjEsTifVm8fV6Wj/wpZuG5BY9wgFHp
UFKHxXy9YN2YJLuB+5BUZeRnjFFTrqG/1ZCS6Jb9MbSlwp9hoyh1gfx184G+ivdn
oqH40CKKkcNfHrEjf2KKxuxkq0QeG28NJdLK1R+cO8Pw7PsyqLoVJHlP/7lfVwgJ
kSr7/TgYYU++J9cUvWj8+Ag8PoP43gUVWbcIPQNJ8MiZnwy5UPZrQ6zQdzeSfRtm
7M43Bx4VkHjCa27TlGlgXssBxnjT85r0n5ZSewjhxY0dqIb6KvllfnZQvflPSEHd
mHLub5gBOOwfE/yN/P0oAvwVVCMrY8JcLpTVOPFq94sGVhGEpeJdz92IK4j8r7sl
Tuw8IwQcHYgygyUwjtSHDnlwBt8fVdVY/O+GTh0vWV0o0/0XMxcSxpl8jRFNDXuK
l2R2OAS65jZEYsZ4EZ0JiUtMqjSkOn3Utk1mL+EF6bAsu3BAvSpPsdTyxAH0p8Q7
mrjc0wSTNUbOZ2A/hmDuNlzOr/GpIUmgQmg40NoCJWADnsIw9WlmAMsh0XeEQXM1
Hx9W3Hed9a3lqXgKam35RcfhHuIo2MKIr7B7z9yhF4PQT5RhwDwoNACSFRuAf+IB
BEJDq2Qekp50whiKjledWflp8mgFyd6ZmVjjTyk0HtBba+x5+814EyhkuLzPyEYS
lU72U9ONUsT1y1FAmpvoLhVKUpbkrhEeD8n4EouCjJm3Q+dFC3pVCojqIP1jtsGR
GjL91JQm4+WryTX6qVTGzFyWWoN53z7nNqr6MciZ5RRUbqQ3Xk0IuwGm9T/9vUz1
UNYqP4tIY2AxRmvzbsXBhx2SqlcuLd1dQ2PTg24T3wS9FNP0LKm7TH7k7CD0e3RY
+xbnbfDih2W85JChNox9zDTOafa7CV7JpSxVSfOwN4MhKUZAoZlHxtwgOhzqf+fU
v7Fafx8rMyFRV9HLcCmiowjuJcY2OVTc1CBNLn5XD2wSDe2J/1dxN40NfbrmPJyp
8+ZJHX2tnAOy96LrgzeezAphh5yyeSZPJ4b7ggoZwwr1A1mZxMekvA5jXIRhItkl
bYHN7HYC24/b1tuMkfvlkMtJMYCTEeqtjSrZb7BxTKZ3STYf2zKTZafuL8LqJFV3
8gxPHrWKGadqkTbvIfTw1ZnPbZFIg5AO65XBW3UuNNgOJXZtS6SrH/jAR6KrjotP
5Y88E6fIavfHtNs44PogkVXuJMVp886TMIMUPH/oYB7N2a90VV1/D3J25BloUGJa
1FYUjOvvT3mgBh91/CeB4Vob+Ta94hKd8J4ZWDmby74fn7z/9IAc9S6kLgPNXQZE
TgO0pzYV/0ufzHZzv3VTIHsMaEOpfUcMY1QFC2n8EtCOT64zYZxYu8mfkl0nQaPj
0I562hqwb7KOE57KvleODT+sD5vTufaBWQYD1tpVy0PZ9P2+sVAQD2cSS/Dhwrjb
Rl8kmHgfr1y/97v835D54A/VQ8krxtjm9tgM1crb8U/b2r3MzTMb/wREN3HrnASA
LJTgtYxnzoxoy7CMWqlHzhqY7WsaSWLJ5YELOxWLFXj/oESyN7tHwM5DyBU4kUec
7isCsnQ5VPseR4kwWLrhZ4K9XWVB5Hl5/RzWzbFA3lXcLSg/nbrUyu0zcaC4sDwD
AOSLTEqEG9MKeTq5mxQeEFyn/HdFLhyf8k7u+mwL2j2epIktksDSZnqCPLcU5BJi
sA1d+75uC6KoyNqTj8+df6ijdqTghHtzvzqQS6mGJ1fLIbsO6Jm4zt1KtF7dMMbj
ZnAZcOViDubsOEJOWjEd9LlWpbvP7xEAlz4GcZyW550vt2hZSjZDOj8d9ThgXRkx
F6GsnvFZYcSZ6WuwYppBkAwNp3f+BImEpQ42PJC8SlAXsJADzFYgdW8r91iCZ3CU
N4kuSwaCj2tuAAuK6y09wBbuXlrPxeHGpjzbqdo0n2mTVnjil7CRkLitfAiC+xET
hUeiys+NTfjFqdUoe8ViVBfVPE7QaqXH777ZFcRrbzDt5um6h6aJQPdk0egmIynx
UYV1iyZnfGMPhq0/u/qHUTRJi+agsZcllbTqmliD1ajzc0YDsa3gvfOmoNbTaqml
LTJTy9NQ07RjJor9eLaJIj0IMNztP0Nxt76HghkICwE8QE57p18NWfIdSqRnlzpN
GfTwESqrJ/wK2Lmkn+XhUd0t12bB0aK+8RXqpuBTQOvnlQGf42bYhts2J75wzvN6
/QoCdQGNU15eYP8Dd0zKEI1Upo8UMJ4oz7AOapOpvvRsgi6JlaDaxRLZ2arezTmI
m+ky6kkxlSBMcPkV5ET1KIkNygczpOJf/8zuHJA3vNcfE+wF7bIalKG6RULMLYwi
lQnGK6/Dz0etPVfdKy705Ke4Hh8xZje7eNmxPABryEP2hIqHXcQMiv1BVQHjJQ2z
Qt0Im22RimcWgh9IOYvC8N+IsmJ2HWAMpCkDM16wBbBMCYNLX9xIz2zSZRP3n0DS
eDSqZ4Kd4gje6xMl+80LV10NDcgWwUW5cR2LA+TX+MisYp2PsNVJQcgvWcXd26vK
PRMWqiMWaZS18ElgVpw4VzohtJ28Y8jTlgUziWksK2WNPJ/eTENAsbxaeWLfhFx8
BFPN8mgTsC0Dmdw+s+72sc5ETn0SXnnFHHr1Qx4bBrEK2IoFhvvvc00jc7u53Ouo
/z4zXMW33xpZmBX33sN5OGHeKF6AhianVOuXD7SUFBLn4HcbFePRb/92sCppx5a0
I9iqD0TwbxqGnNm9sVZ7afZ+vxXclCaFybrn4WIINb/D8nHZ8JNc5oxPZ3qJwS1L
zfM82kg/ZqPS3s09dcRkf/wJsHHoypt5ueBCBzLWIJFShYcyFN2pUCCMLAGb+9Kg
MtIxIIB+/WkRVuDH9aFkIWFyhC3HZ1TUV0b35gEmqd+vJMrPXZYQtV02TcnzOPro
ql8I4ixbEGfq7bl/pcvVyIWJxxwqbej0ApSsMz2jNoPUfvxjBH5d6BEyFxL47Tyg
BmzdqjX0gxieIwI2EmQg35Vuy9JuJnxm2HYVNMyagRpjePOThRzefECtD3Nr5wI3
JFEhFMTqxXYQhHANOlYN8LLvLRE6NYMiMINY4DwE7tKS0hn99CFbdLZjBuPyypGI
WR+KXNoih/LgYY/pzU9eUknqorwSGddNd7+tqWQhKQW+4eMOFACc8S6tcISA1gW2
oMxkMInuBVP5IjFuCm7EDCrf4HTEasQJathLcVUZMt04gbQhXg0A+wRnfwo2+Zn4
sFSRycdoX0p5rli4m6K6R24Xnx501r8ypbYCuDzBzifkqkgBm7CagmaWJSpZIrxC
jmyFiA5pHwEhK34LJ1ECnKoHq4JbTamdafiVe8OnqsR0oXzxcA8PYVX8frt2gyub
O68iDoyLLOepOtrI9HlEwE0GlhpqLIPCPocW4dIdKSMhEP+T7sQVXI6Z6eCs2ZxR
Str6jWeZofmcoOQhPjpbJhnc2O+D7zIZlP2gVdaQxKnMFDwCA4YIY0feVxhCpYLy
oSGqAXGD+kEh9S52+r/ci1UqtTdDVtda0MaQnl1onfbXLwKf5XYeV9/GDBbYA2YY
7o4TE3mHnkozGuIJeMPz9G5f8+BhofxdhLx7JavKhBvkejTkiG7TjQSQuz7gnfS/
zDsYwk6RJk5fZpjDKpg2X2MT4lkX7eLq0tZj3PvkCjLLQ7cnWqNAigNAakilCYdQ
OpsE62nal10jxAsW/172FLWxxY3F02Gv/kpzjupgn0tK1gBW/1TA1M0YmWE8vDt3
NfaBQYopsBvUZc0THkRvYKx2JaYsZUoRzSLvbNPQiR8nBYsR/zlSrFfE8LA8/DKs
0uptpZnKotNJOVZ2lxfZx3bLOseRoFWogHBc0Bs1GLc+KIKF2nAG8NJ13dkYqw6b
MI7QHCblNmMe7XAIdHADVuEgV92gL4TjZ5lTsjgG/Fodccm7r7ncadqdgxtb0ycE
1T6ccMVE3on5GSKeiasXZMImk2iiwZWvKuxkWtYSW4NOY/HsmxSpyo5vCXeDTND8
f4ztCSCs/9JSc/mey2xVNMo+RA80zp2ZlL6gGU2ZH7AZB9CgLQ6e9GsDGys5IiSt
EyoYCU6RuUWiKusoDhTfcpffHfF7aLZaPsBh9ZnKPJQmAfIc6doNwhVMh2RSuED8
uliXgwhnpx3MQ+tdrXRzteD/gC7t3mY+dgib1c9ReiWz/eDf6DlKz8+dXCEZoR1U
WEB98eFlKCPljZoUNXcW+tCQEokgbclzQQ1UE5iJq3EGtt++qBl0tIinaxNpCJDT
UG3xG2caQmW3Rye5+BvZQE4CaLPWV/JcwRaQ9t1mDXe3vyNy2bB9Y+dwlV4Ya81y
tQydReelwdw4/2UUcCW+xnFVNkx8NFfpnasUFktqEm2vFGWG+dT28wbwZs+HFzLf
apmpdnQjT/V/XofPfKtBAxZTsabOyqcjC4xsI3c2TRcvYVmnBn23idAxN6gnLGKh
8GOGCxMmwD0VTcgPuCWOXdxSfZw0eErsOpVcqqbEEyzdOFezXBwDcbRgXrV1rVV/
qlDBG7xrDbqxWYpze9sMVtjhozgPD8uw/m4zlOYD1Z2RxNCz7lsKrPmQkzWGF/W4
EHyLFZZ1xFijUI4iOyqIXBhdP+mqsW5CknLTU4gf5XaRFq79WKJLtIQf86l9nJ5F
3NzmCT84NRdW9S16aPVDg1O57vOsIryPoc74ilfQWhhBaf9ZRe0ywdqsYbD5Df+P
u0gdGK3+X75avDaSSxZKsitdwqwQYq5N2BGxrfDP6yKL6F3IzKNixtxc8ZFWv66p
f2N3p7XU9pufVjA4rZBw+Lq5RiatCZML2mf92Q8OVzYxDndaCDPDb5ZtmytfPIHC
N3JcvJQ6p5HdfWvSrIGZbVM7tFjE+CTfZvPwGJRODm9iPsSfXTMaA+n6fneD/xBc
5JJYlGSkJXFBVwsNc0pbLtxEQC59SiXcGJonm5td4iLGbhf1g8LIDtr5I5c4qUMB
JVDyQvhbEkrDIjbz9bdQHvZcweDP0kH2RbDu17oRcP0g/2SOJMw2nHrFqQ9iz9bW
EeemvGFZ45jha4/3iWqx0cLhQ+elI7mROTvphXsppFcKDhmJamoH1fvtU0A2vjSZ
jQEXMiCz9Kf3mKPGXPrIxMgEQOt3eqaB8wKcHQBXlIDCyySRmJVbyaCIhHxRRCcz
Begu0zSBYYUwiuGLLsgY2KlKwXXzdSgEvrlWSYYtVqlJ8iRTZy/LwA33Ux2aSthJ
6r4Mw1Y+zH16Z+oSfYLXPgu58/NbWDGI6q+q1DgWhRQD/eL+78S4vgusVFDq1krs
WKgEz/m+/kZDy5dQgXBrFcQTUuCBkaChAlHXopqEb7iIlQiq7mntn8D7O6RPvpJk
yL1ZO5ZBPJT9ESacPnby3iCl4MqbE8+kzOzG1RNZGHfRlq6i4AERjcBGfqdiI91Z
W+KB+Jb2ABAKu7DD+K5lEjwymK+Xh6rruKE+mlwQ3JDIrvOgfS8bL7wYNdr8s/DT
bJrJ4ScQ3ZrVLrxyyLR7jXRQgaVGBt0NfmGlgCJMXfwmozvXrtF8Ly/2Oiv4fv2T
AtzQWCYBv43VXdGXloZ49Py/qzDgnaWw7nb1wkw9QIv21qdBKCxTL2yQhFXzNRJq
ZhBQH7bYh5dwITYtYEW6X7ZvMab/nOIIUKSukm9C2kAd5VyqPUS4kbE8kRuowcda
K1BGossSONFhhSybqavWF+v4n+rDNSJsrPR4q+kvYTMYrA5Q9TKgE0psqvdFJwQB
LlqploUo+0mHvvsPweJDlSZuNEfrH9iNmyCY856kgHUJQ6PY0jMrdiSaNmD2cxBj
UnlFzMgKlfP1QSN03kfkF3qOTKg0vmwj6T8koR5y3CtOzwtlLmVf+GsdmMSHfbo6
JBCI1dGHkOeZfKPsimhNhWoBlcUoQTJhqj1MLxg5KDqd4JDUMslbb1+kTjm+X0DK
UBvxkFR5u1H4y35XMaoOpggRKjGrOXXDdGSE0/6qxKS7iKpxx+ZIwqYZeFSQoJCi
cNh3JZaGfluX6+HsW6CvhCmzNFY7+Q3P1ekAPKZzJbE+xpnozHxDE3c2OPYXPSoG
1PCb8aq5ojX5q6yAUcHFv51ElLIP26yFtc70Lbf/zEr97Ves6kTFzH0rPQ3AsUe0
rQwaXHyDUn9s8CLjPHDes4lBeG6kQU0CqRdxyRXc0U6MxRam6m9ycvPdSoU44wHN
fmnCzvrKL6JJ2WnMs8DMsttF1IRPu1zDGIWPzFekuJHnS6W9zf6uqrcuNw+Ho+nI
lv7SmFGkhDuW0bpGqU7W2h7F6BMIM3ZO/DtExaEXYxrOqfM6KHHBujT+p9YZnt0l
zhU5J7Wu473/m1Xg1hl8P5+ym2ptpZceT5r45qL4spv24bcZdfZL0LZhzcyRQlxi
/aJvsPrhf498NKyheZ3wXVWusaHIcsTO4+2FvuXppDYndXMsIa88g1LkPtuU49Pj
fEmhhIBrWSGlNN0y78eIH61jVVYiSSk2+bL6TETBtiRt8BXpS7ouEw/Lm/+eh6DH
Q+zCS+Ar/BEZX0Inw/aS0fV2aVcnF9KbCBrWaN0gI1Z/9Q+hhKSI+H+OxwNJgYCQ
jr0zA5BTphZ3Zo/nuuEX5UPRTRrDudyTFt8/RfHK2Xm/nGDUIjb2f0rqXWVjQwPS
1EbUlSvDl+cw3xeInMXXFI4wE0mxdMvIB6K39LUn7AJeWSg2rmofbIYc9Vnn44Ni
CMGL91sqKOymG8xilB+gjcL3ygxMfMKZ1Zk795kLuAZTYn0h3FlhBo8jf+uLh5YU
8nbHjDISat6sOjgoJ7plTbSEUqs4VDwexngOmEtl/nSstIwbxk9nJ8AW1BQvajAK
sadb/ZmNN4et7BjXy8lS5SI1TErTQ1ZnvqqEw355h3X14nV/8w+ytXhv/EkpSG4B
n6NFMcQF31fwY4gFw1kCGXeQVwkWmXeFEF3bWQTu7q0fSs/6X0qd7Ln2I5ys05dQ
kGSPUYPDXTwPRLRMG6BC/BqS96Sd4jU/kwk/q+ZSzRLgrcCLkqW/NgvOn7lPcPZb
6u8rYrYRydr+QjJDo7vsKAgKs86mq1F5tcjW1WZzc98d43B4wzoI0CtNwP/YWi1M
rC40e2qnUgU/uw4jMUb7csm+jr8IPt9CrkMvfFBDoN/8M1asWFWKIjgOh48eL10X
Sxc/BPMAYDOsoXSRa2pEjQ6GQzNitkyOegb7qoPr5sGeeFlG1zv9PMOwqq40tAl8
DXn6HH/dqfgpVvTIu9+tQ0mbngrOJY5IkjNNksgxd3k9GKjCCIKQSojeEOcDDb63
CrJMxQFaUoeB7JJ6mgK6qtD1PvuNGx8OhTpbYyRYeTJvMVb97dwAu6nhRRutmIeo
7IdILwjH0Viex/KRpAY6fnqiJWz92n4iBB1b8D673ZZWOzkL25sdmD5Ll1hQXPbU
2k+UdJ5M5rh2i3HxHExaifg/auxyJDyNG95HjDUoc+wETZ3bV027wyLdJTUCD79M
03ag06iRk5GDOL5RtDvoBdDXIOC9LPMgYBufNfvLIGQDkTl5jr408XEptThiFGB/
nlbAz/rMLCEA+NnFDVwZ96nj02Ub4q8PM5Z+KdA7euwG09ubEWyBets4YANU+Lr0
ameJR8lKMWv6zYDldE9Qh/byBeVMlz7XqoYdUbTlU4CVvJaA4cbcNOnm4Zz1xE/1
t/SmOxC4qIh4aJyFvJhW7t3QfsjQxSITmV3/bTdxAN2uSKlZ5xAoKdoFGVbmYjgq
Rfx6UeDPQkzaSzfvemegLK39x//jKzhBiv2QhBD5VYT+cpLOVHO8U5B54Z/A6Xdc
0FgMhmRf9auaJH72Ho8uB3OV/h/N/oZHX4C159vEy+4aN3WuNFp0FJ5Kgpy1di56
jdPYMisNmGcCXM7sLRrG0ay1YAP6e7kWEDMHb7luz+rS+MbJzJezBN1SprHh2sXh
v9/dYom4WUC338KWmlXuIyg96Z8y3rdlXn0546AoVLoeDnnCiLhFD9Dnc4gi00oC
IgfEdBqA2qIGK5ddMl/wQGBTIaNomi5tohZdWosICHNrxtUUlQSS0yAp8qSpK0FF
GyNJrXY+KoCnzSqa9u9nIId9IPdRNZZSqw7LtvQiYSV9NnMfrH6qRleicOHEHyOI
wpHl7WcgCrZ4C0nJa6M0NMrO/MHBrk0PjrC0eVD8AK6eh+g/pG3/PtRHnD7W5AqI
CxQ8pygjEvXdR9z7rFIvCMZkNA/m6HeBTR/mthmFmdSPJgMlkau5qEdTVp1kSfJ2
jQ6vVoAgM3i4wmyih77XtR5I6PO7YKC26jznzLYthFVZ3rnL69SpEvY5EV9kbk7D
mBMIFanwQ8KEGyFK1JxYs933EsV8E7OrMsaYlmKG2WDA2KrPtxCLmSv/8tZdv79m
oBYbAgKRx+BDEuIMXzLLinEmIR5Aiy2pXnsn0//j+cglRbgoKhTQ6HJ+sRePUF9S
mJr1M7nfknJmjDfYQcYPdLfDqnZDoofJ3TxBNl7wpZ5wHeCD6h52+DDJ5vto27Er
yVoHht5WDZi9NhOvM4rb7lCq/7qs13YZI8oNQPqsyzmBBedWR3KYOVEtOk8tm3h8
2L1LmfcMuIamjP4OSYW39gTufUaSkBNsvM0LnN3QsG2G9uenwxfv0bShsWlbb74t
cfG8ktzLxFyek5mGtGawKb9WCGbg+Oct52nG1hD+TbTAJrn2Ny/Og0Mgkj5y+lK7
bpc2D5cKTlIxZNdhK0vyIzVWKWna42G6yrjbe9ZilyyzOAuSGiIYQWmPeDc5fI3Y
6GKamqBAFkt4hI7XplPSPOYbOyWRC9JXxo8kKvn7ek3y1AkSeAJXok8rizs2+6Vy
f6sDC8d4y8KLOlzKqtwzrIZkNylcInP6X5kltzkyCRbD5iTqSqNIZeLrztJqd+Z8
wSija54AgdcUDj0U/qr1a9NjfaV8vD6JKG1YnM4jexdvmTIdZEe90J2nt0cxDDdP
WJKNTX/k9LRpUUnhVoqsqR3EdDAUh2ulTyFK14k1VATriamAJyCtzt8KvNlGUkNf
KFHPWc6rE0HiVgASNGJiVKNuZT3e2QWyz8Md1y7va3XiiROuSBVXYuPUpuGewL/e
Qaeg3XuEAU1vt4shEaSVLRJdtXjUcaZVN8/h/SfZIybu2y3VSa/hA7xuUU2RER3W
ozawudIFjyQwPDGsZVlyVlqZGn7+KtJ6dSTMyDJzwIk5i4MId4/0vZ4XfxTkEIpU
bkHkQ4+QqcdytPb8Z8g/wzKG3EbwBabN/7UCuXZTP89Edzse1/9dhlfT68OMl+FF
06UeL6WcVn/o9bOum/rB7BTuOmZ+fyFxo2clzFJXtT2079E05S5yLRV6kEHh05Pi
Eo7hA8doMwHMbmg79aZRzZe2Ry2pvVutp8DX0/JKqqHd0X5OTexgtU5zqdmr/bnO
s+dfBw2Tzx+m0xvoJIzgmAhaYZLK/buzInVur+RMEQcJRkHCudHWVZx9hYBTr6Rd
wXew0ew5eH367YQWuA6aEHywDd2DGIDcSoCZHRqXnsKL71BW5w2gybnJKZ1HGW6I
nDsBt1QH+q3Ufan/5tr6wRFO3dxdGok1FJkycpTgEdQxZLr0ue6Dg9i7fUletvVB
2BVwK/EH7Qjvi2UTogEqxI9BgRFhGh71zq1RSGSPvthmlvFs+MGFEV55oS/EPLSk
L8sHfsEyZZdDi8srVeN2NbxwJfoHjjCNOZeIchpRzy1grgeg0kRHAvKoKb3Fwe9Z
0/Weyd+VtcVk+AwbCtRHNMfi5cB/Wa9xqUtCKDRcjnGOy4rVyqQyQKAlbcq5L+nX
KgjTbEKkwo7ZJf7D0fVxKS4dVHhJqOpLsw4z7l+wtT+Fcic75m54N297SrEbS8Ei
OFaBE7pRBihuugtvADGDyNm6y8AcRkt42GnScPN6XQsJZGtkAvx/4KPQtWuhrWeE
hz57hWVJz0b3b9Seot3nFSZGS+eBieMp1ziHarSL1e7hP8EDpCLnK5RQjvo0Hq7y
tySjDka7B545UMB0sW/hoAXXt57sHsECRKKzYO7jJFYBc99tIMys/mvp93raBLw+
UGVvJMajDWv1BxWUaDrgbhdtmetqbrVOPJS7w51on+2P3h9H28eP3/Hd9WhRhpnf
SGlT+ld75UZq0SXmOVQKMBFbZ16WEjQDOcqmU+F6BpdIR9sIPQ2r5A1k7pm/N1b0
HL134VMQhkpZfu9BvXN3r9WQWsT9H4XKjh1CoOSNSR9AV4SWbd1pCTSei/iVcfmz
/lBSoV9WIZIAQpf7tGHObxvi43NW43mq7gwW9vwWfWK5Id2Q2QbnFK+72RKtfXLl
Pp/Qyf0ask2YgWjdmVWpH40fqkxipH+4REp+4+BKWbVxGCDLiA04lLNmW32LR638
R/69+PxKkz1pcf2zLwY8R2Q9eT+j+YOWrNtDPxmQJhvzlzAYqilnD0OPqS+Q6jNH
Ru63zEfNmJo6Jq8Ey32oRgHl48A21s4ABqhLODeGF4uzcAhVACx0LZ11H6luJoAW
I5U/B8oeXnivVxTltYcehA4wYeuRFFRpa4aS91n/WbEdApoM3FU/OwfJe3h/t2JA
+nLirNJdJTFHKCCNgNwnxbHUBx2aD8651souk4tjxmufBwMWkGqBU/5wsBukjLAy
f+dprS667ErWeNLACGVOSm09o9aI3Gn73YbxiXIFwQF3D2zpdLDQeCmaR6PmwP2p
RC+LGxKj28IJdXVbmLSCO0Q3nJSkwbpj6+uaaqb2AQ/2Lka5cvRIaWlxRLSR2dOX
G/BQKrg3/HqSfZV62S5qbRuz1GIw/UuEh3AS+BLBZbs70sCQkB7CSOraNgLyFV9E
UV+kcgHGoxERFkz3RldjfVD9GpPJW39HRCdvANRaZJZp/WIlLVKEEyw3kYZJp7V6
nizLWtAg1Oz96XHaNP6ZpzeKLImkND44GRT+YsO2gP/BsSkOUmiTuWDgIbeEbSWj
UtCpi07OBRzXaXe0T+neSr+4KEQiiPYUhD6JTMFz7T9EXUmIDKXlOhdi8du9/cSx
tv78Q/lcX2PkoTbHlLH4BLAauLNZmU0KWS8kikJelyUkBcDzNvkwQibOnzDDVHhg
yZEnpPO+AfLGRvfcED0DJuHHBflIaAQFnBZjSMs13N1osCoIH5z3upeGFQJxzHs6
Tov/RBmvJ47/i9Fzs0WY16UYSNiQMNL3KWDyWHyiivt7eixaa9IYOYXqAsIetm84
DX9qZwEoUkT08wCw5WsnFbQFWbeL1+q3s18LFWxH4/tQt6zZFSSEQswaU+6C8RqT
su66Xu+8UaB9r/qy/ev3Lj5dftqVoV4wUGDB/H0UhYTCw0+FfvJVYA0LJP8pdf+B
NOHG1cnMLhLkcWvttMdBuOcHEkZfrYUXhNK1XTFrHaUqcAuaPo+hxN+YVpNHNdOC
xJ4feMSk+y9/HI1k8vyuQBqmtQSGnXJHf3aT7zrVmB7506FxU9+mtt6RhryKkzzP
g/Q7Z6vgNDcHIEViJE60mK1Upmoez4RxaX05MD4CKcAMJtkl9BORbtTq6TmZpGEy
dzShAFv8y4LlTxtTuJVMpfIKipQQirhLy8WHikNJICSEMUQ9C0yv8he+zS1QuBUz
/Lma6Zp0S+XdGqVpOmS7du9+eDyHIry58jhLjmrOLdhXLSgzQsQ7YgD0NTDMZqOj
jRkQbZSzQWYH6RnsWO58lCj1OJXxPbKMLWXsTOahCy3L3q518oYtZ36IrQJo2GXq
otT5pi3SyjmLlJgdw2mLzz7+pI86H+kf3QOQgqQKunMHJuIFxRxstqc5E2pkubEA
hfGataZiAGRsAoH7yLLO2IkRUPWWqBF5R6TckUDzpLkz/hHA5QXeqwscEfJLxJz6
BM29hMjtPOUv6iKqEj2nLWoO/fRaJ2fAW0KB6J+3C9D7asPaUbnA5EKD8YxVh/1V
yWPMHkc1M2s+Z3h7YzcAFfCqwiuf+8jxuwsIT8mnMfZXGmAAcoeuNxbFX+HBP9Fj
LQhfL1TnDuK/3QXy6AxrWOvMOWRdczuqr4GA92JmJOhcBO6C/JaXbfLdKXWD6Yx9
McaQDMLXdyZD/vporaa+mBm7UmhYzj7UIfcibelJRbYEG0X8SybdyyUqwwshRz6c
APbTbptT8kBwl2PYNkKf2b4LqGQ4YcqDPKkHm6W8ISJcaU2Or3lhcq9ojwa1/FN9
JeJRdXMrlm+QluI14rK3++AuAxh8mxGfbl6h14J2EdwdyIu4GHkV3kTjfaYZhdhG
jFG4xYOD6PRSOcON2EzDeUlILuaQ/B80H9e6vRvvBjsAa6c3kV52MPXpegmOG3Wl
qRaoMOnnxrNraPRKfm0KaOf7O70ZaNeiHSKbYgFul/F7q7HzmbD+P2FCwT/V/fGS
xY/BED0G7YYx1PN0eEI3LKDs3B6QtEvGOOVvhw5dheQFaggdgUhStXBANm1yI1Ip
vyvvwvBag0U+LTHZrnymoroqxHs6E2Fm6aN3f1RukJnra9CEXvt5AzQ3IXj4vQ7L
ehCLWXmCRym6YGLKy2HQmaxisufBSAW5URIL/NbeSD6o9OD9ppGkVnymeGG4C5F5
kR6gbkYY+d2+5HjesSm1sOR4Pwo+UUIGqOuKZLVI8LhS2QeP/mVsNbcwOwWXPMx8
MUduiBO8U8WqB7WA3air2qGYoB7HdhCtdLECj+41R1N2Ifl0q/ivZr0a2sDOCphA
+TN2QN1RFYH4X0Srpjb1xdMsTid5zaYKV25fErO6ODLGxxlEaunxxz9xCR/7Ozqe
yy2+Rg5JzjmaDHHRxLCTBpRGfD2R4qQdGaAg9Q2SYwIcYmhHEdLoIaiGl2OvtVY+
5SQYPNMZWfx3DNykxph9LuFzT78are7ASRMzSgL6IZ57BRXI4CYjb+fvMDDAAsas
RWab6U+Y594GrSF8Afnm/AK7kVBpWubqi/QEAddSyoJclSjbNP3xVZ3fcKaJGAoO
Zj7gny8fKX7SmRkipNOOYhaamBxe7YqVxuLnm8RBvmA0DC/jbkXd+F6daWd4c5Dc
WAd6Do+f1ysIo7lIB/NlOtBb40MGegS30O+FsvxLI/GGwqFM2K51I+BIgVzLQMR+
HF1N9t5CdQ0/m0Z1u1X+nKp8+GAC1Be85sZTbc8KHxsPiO6KfOkfweS6ii7HplJQ
YYW5dIv1OF1A6F/nghhHKKVixLTGtCEY2GiYrc/CC4L1nb7B1382kz/FySCpMwFv
CH7c8f4hYFd28vmkrOlATRA/EgE2YV16j+4UNgcdvk0g1vLJXB3yYaKZb4S9Zsli
m5eBGxl8pxG0HS+tl6q93x5z+Xdu0yYzeFscMshTbp+V0MSJqiyXQLc8iCrDdGkI
AAFSUnkB3kxJAEDsojrAsQVCeFoPNYIMboCCt7mRuhYQnDMI/Gv4FERXo+I4f+dX
OumvwjgC2Su+G+I+mvrsdeQGKMClXbBPMwn3JrTQNFutvfYHUHiT/0ZCASbJ1WWT
68hnM/KmvRu9n+XwS74EFo0W6AX1dTovXtRIa+F9i0SqJX2DaYKUeZRDIgM8jULc
gVsby8UnohklwP1OUNovk8q7yO47UhTkOV48UYjEPxlB/6azn9Fx3edagXW7OcD+
VVyjueDs8zFbR3AaaqHxqGVhZqG+MFSVhKlulu8mxCeJXiekZHYXDiBLo1S1ZWlA
6Swnu8SJRwZGODs7Zp+PN05P+x26T66aMWboTIcBE52hgdsT/Cxco7y45tps7tdt
g9qtOe0kI4DFzDBEA7zMHRQyFkyX8CJaK7icTwmMo+D7UReLwM3Sa4uXc6KVCVWX
n1klwso2N4LYXeghhpTMnTYm+fEHc/gwdCyY/wJ7gH0nf07Gdp9RArYf1mmytdgc
2BLI75mf7U4Grr2k6KWkDfa04UGOfZpEOaiqFI7jyhbFo3hb9X6dbh4g0yju9bLE
5qFUwDB+XpCQiKe+ZuDvgEEI/vZ4IqUUNBDbePU/FR0j+9FlkItaUd52DhrmV9ji
MBP17JLiGO22yupib8jTWj/+o24D0AIDD9yYqSGYvyAyYhpEnDazUUoJpA2/+Tab
57J4AiZtUYXY0onFtXEDxV9f6N1oVjIg8G99VJn/DYBvyqD6V+D8lM0Xrb0w5vnl
3BmK+wt4Zt+0GCB9VAnJAR4a0ZAI7NCS8VjHpo3QFxCoVvVds9kgysDf7k4w3g1r
I1gLk3kL/SlilA3VRdZJJMgYWSEqdsFQFG6KrieKzzRq7ZwtXj9610oboTYX6/Yj
BY3vDc0mWR2qWVGu/T9Ofhp2uKQAXn8KXFE+z5lS4vcU7zjJU5NGZ3XlcNQpn7DH
js4lcF1u0iExa+TtQcasgGkqne4V6ynem7qC0JoD/AepHb1jP+Rz4P1pAV2oZw8h
eqX5T2W6e53ucBd6OlqNcm5mn9hupai5/lUxNOxOZygWMOvj2B83wBfJfUtPIWur
0pHO23K6l+gDbqA3eaoRevD5D5ipesO7M1qHXaeF8KzaJSlyUGLcpoDILOX8yTM4
eTNptRn8mZssmfKPa2EzL/LP47vc8zvYmuaf9eS9P3uTLIWNls00y7Lotpsn2Bf9
yprSjgOmYw4bz5nGv085SPXvpJ9zuvM7nOnThZBKAZW7jtPBeY4DGJ4z+gg/3p4r
zzwVTb66avM0jz6RzYOV5vx6dOzMoRejEzhgoml00J1DRRsaQFmo3NCtTtF9OI6S
4yonYH24U8BP+TrBTMKjx9aYq921TpMysX29mgsR7xhTOX1RDl35eN4j2SiZvIOR
M00de/tqXe6dl4OVmr4iCKN5c/vNtmBu27nvY1/jl0cuPyHod0S3foK4nC0wQcAK
skKR5YvkYADqKgiVFX/7x4RNDfP+adll0oJGaM/lJpm7YDxIGn7wUt71xZkEwRA4
OehYy1XXg0ThpVpaWEKHWPDo+EeqD50p99X1qfFIUwccbk3DsvsMC4j9fc6nJq7i
KeIqVbetb+WWH6thuwIaltq0pnFYZDtaMaujeO6k78sNZS/imzWs/BcB5q1DhAmD
9kXGmFKTbXqp1/+i8ATd7cH9xEZdLgtB/K+pL5mk7bdlWLCdMskOZuxi0DNN9ie/
ym1c0LKIOyouFBwvt/OlZj6NNbohmBUpM/QfXFkmKfUXcIB7SuEXcXWmagJhjbjA
WqgPNAoMvA5icP9zwjXYwgqGlBkCkeulpkit3vy1+R6heKcGIGh3wOtwJKHEym+3
RTz0L9T0bPUrqoj46zrfg1JPcmu+6IhSEXfznW5skXWvDCVNxwphEqwMTmak8dF2
7XdYd1dQhiQdG1+VrtpZtG6EvjOc4HlnDc0dT4M1vaXb7UbT05+X4flBvv8B48uw
PTIgxqZA8CeuMfI79rg5hf6UtsjoCiTGe7GP1zotCWFyQoBm2U/7gXksCaBpCz6P
lb/zOO5QUNtGO8NCCveASO5twW36YKNP4eZytzTt9lkhrvW9qokvc2TbSUvusZwU
gfK7OGX+0LKxtLSOgIVbAmRMUwXnIPRE3DMNQSp0a1etfR8t3cMuba7tlfBWnWai
QtvFP8g6notknFQFqXvnnQwhxwT8LxlrLCWJPss4GhDU3K01sull5Uix8uV8ErSl
n2Pr2wYIhBbUXmRiePt7F/XmQQIfUl05/RRjuR58hRxB0kb8NUyDg33TJh/XXUYn
sKDztwMZuKLlCiKRA+wNP5DtjBqx3A3GhEAl4TaRokPI6M+UPLioVWeCOtHZjg78
jhlllR5fzjax2RXcYwM1uNbFx7vP1nspRlDocZ9Tkqin3t/oFUkXksbNvuuBfEJW
1K0/XWhvxoP5iN3vwwhn18Z7fRw1un5t1NdQq2ZB2BOraP30Y44zsRoJK7IUA21l
7PM8hBKmUmNWKimNpUtJnPK+EY1OhfoVPhdT9haXIaiMaaSg/icI9HxL2cqB5uUe
8YsqVBEju9QzopDl24Cr2t2+HYK6ssUnYyH4pJHgEjyTPcvtSLlpBIz5wjKnVBnJ
GH/iadX0Pw53kdnuT2UWsV/sf7OYe9yDvpIm2pX779v4jVazToHFWEFfqnDSMXdn
supSdscDZmWaSPK9fJZ6b6FBPDyZqYvUyobz5Vw5i3QX2A4iPp6FsAWKwVf2reyM
nlFbFcdw8x67KBXoE8eeLnrgNE95wGmYI5HNhnAwiUzK4dna8NhOebIv+VEV0Ixn
m6318npOspyifueEqfH9HzSL8uzsmhqNE7A9fyap7p5hxvGyzhRg7p+KgNmJkkPF
q2LUNcUWq0NRQRchjmoUup+WdcCO5sPWoHBqPNtJciDju6cRT7AR4SVkdyPf6Mt0
Q3XBzHqLwfeziP4B6Vr7j/6qiz2FEAr0Dm3i9qRvdFev9LO0nc9+bNAb1OfPwG6F
N/jUlc+RvDC5L6ll8bLW1xQerkrNoGsf0BmWd3icRVwgzmk1u4ll4Ig+xSXCIrr7
d/mUyyGz/gQiJhKygXrlMACWQCW9mcK1JNkFFAS+9w6DqriHEDac0s38Ek8d7Mpy
99JqrSq/JihK2ZNWqpM28e4pYbld1quNNSzJXi26m1Oir1E/vQiEltBchQ83AoTg
L0Mpe7rQYUnI2w70HEzJHq14YPgU3xKwoB2P7/yvhZ0TQLasEGBPqKr36Bb+H5Eg
20KHJEdm5zN+sNpFanz1QZABT4gv2mXpz9zCv2tOs4fzHGdATCtr+n42Owzztjs6
llmKsZFxhmzmbzMq/+rNWeV5OHxOV2nRZI1vPhLeptTfqgym3YFV0ehz7R/m9S5D
Izpcd1KPeQfZAEo7swr1Cx2HXXKoMjlkemtDXMnyEKZIfRB6HYpP6Saut40Tql3X
43n6UdDrRq1I6k2niHFogKsfDomqa4s3v74zOr7Pq6qC3USRl6ChKJ5srEjJH3Mz
CQMn8yTChDHOLp+yXrdn4u1Deu6mHcb93Bc2bXOezpDbXMOkbLt8vV5PEeaeQW8N
5PtKmWWPUoM1eNX3yiciyDor4q3u6WPs5Iqm3buqUBdw80Uq2N2vz9iXHy8FDscA
74ZBJfiTs42TMvO+b7lYZ1+Z1QzLNlg0JpEsp54sgcWdXjEv6n3X3sJIxB9o6UBF
bEKlkDQBmfefZAMuC4bHRPTJRbYkybDlayoC57wDC9gkqzXSIGmS+B+RVzqEzUMk
5wT0N6rzU4A5+hAkJm7dDqoSDOsU0rC36Vinrsw+HVr29YhcIiT4945rKPD+rCax
UeHdrlVeHNZcMi28BRvsBLrFcu9LM8XHFHUKSRtgegKO+VBcj12dJpRzXFaY7JO0
cTmCDwGo9kmX0qTBgOZBdqsRMLI0DTQ9Rh9ocI8FfDN6L7NZru18KgQ/j03Ra6a6
sCQ8QzSOest1vIKffYdJmMrtG9Fmq1dUlCtuoxj+rRZFildsq3+qQUuxPxIC5Eyu
X24XZjYWJUcyzhb94Smo/7RhdyM+2RY4CuwQyM6oBT0u4LG0j9kfGYEmD6KuSZtj
whcuP1Nmpaa6k2PrIAkUuKE7saNu73V0vttWg30jrtcK7Hm7jiN//93TxrjbFFYI
yRwsF8VYQM2yD7KypAoZ5V5s81YAr31o4pUjJIOSSo1df4kFj+gmDmYo90QquhtR
jiDL+LdxwNwWDZ9emfG9eeic0KzfvFmAwm6s22TS3pa2MAJYdp8nl6io/m+v5vr6
G/q1+Pj1e5Xu+uWTm/f/XsYVn/InUasRAltnl9gBUL5R4G0Cw1I8OcwgP43ekc59
LGSnzgNbq8YRPGaif0DsU4iN6fcLhkPEg+xfJWelidrKFcIIrhaTekPHuhg3O9F8
7FbIpLDwO375U6O/LAxLxDyUbO8dkRV+P/Ql+OHk3fsFB+DMQBJK8m8rzIiXa993
ycAzIkJDoEDPrP7IzNbXTtGuwoWIvXKJQtO++A4F1JUOPstXcjHzg/BK1kKzro/j
gu2XJOQwj5SczLwjHr9I/UwrISTwr/drr1pp5bnZn7Vt/XE5RrYIYfqgf2ci+ozY
Lvb+4OibkZ5juBjPvHZL0jk4DzFWBKUiWwm4w9W72hY3JnUtwJy8dE8RytLEX+Aj
zeqKvkA4Mv9RtDMmw6z5+Lj5jfctmCiOUBHiKs1DC4SCOHbafOzybhdj3IyhMpeh
19NLR77GEVZhkBkKTuCPsUFy7z9QBjeC4+cMai3K19erltJh7M/PVJscxZHTkPY2
GtkIT/UW70DfvmekQF6LbdR7F/E7t447063/YuvduHrA+6iEMcKH60JpnjbP/4Cg
s0x7If/s5XVuW+HTYPPmNvlHHwa/uScdVYmQ9DSUgUjux1yCZt30iP0Ayfk+b3YP
+wfBJI0uf4Y17F25pebDdO/GGm+EmNekrNdnxzMDmlttpbjr5tB3HvLi4dbeSPTt
urac6AjirnpwcSAvKxxpZfTirbHXQ341fQbs/JwG/x8Jn4cba9+fvmV4l54u+JDK
dTFmiNNcZ6pkiYrxjjAMJDfEw6IM2zmqq5AsJOObfYcbtGi9krE/RKgxsL7clpIZ
0vBOEn7Cl55HgR+U8Uz3YxaJ/yFWlFCK3wuDHLNBQJTAXGp3t0I4ZRMiEfIRDRrT
HlMOoeolokOgnaWr8sxUQd4Ouedihx/8f8ohPq0uNi0k+BgefRs2v/9OAnjCHUHh
Y8lkQC70br+K5YfPH3wE6wv/JUNN9Hq+cZuZyTMNYAAID+SB7WHqRuazuKDvxG4y
07nlkvM1gD7saaWTAGfqv9bGAshjG0IDD3mbB4Gl63HFwnIiUJBdjmm08aCwqwNG
4Fmx9UWotAGXyBLELtkqKhou7Y63c/+k0q9j9vo6jmHKZW+9mVaXWFHh7WIHGZwd
2hDpejTp0BdIDv5XykMEymeMJhm2Yz2QQvM9g4DD3NtDfVVHpFwgb7E1QO5DkxfD
RpzLMm8+tX70lqKQ4WbiLs81y/dt6r/Nzr36jyZn3raLoYEXd1vb7MoJqGV+N6mY
F/S8AQ77PXQIOKE+kO/dswK+xwlFi46aZaYGBC8lKXzOZ8lTigi5L99SdfIskaXj
q9ouSHovrjtRxdzhnSVa8cbpU+n3U/F/jXllxzhmjFiny9dWnn4kIDC3chTPvXcl
SAZGjXMuCAYbuMDE0Y9rRgTf1ngpD5zzr05q7ZpGvMEQ1Fh45/ajhvaC9wCtmD0s
P6TP13QxUcZi+2fquO65KGwSQsLqFoA1HsxqUW+YZI5BzPgihGwnyhfda5kBU1F2
7LDaNWZpUMYWxALtIGPQEp1jMklyG7Uz7w068MnbYbIwxrdtW4CryJz8O16qqSdd
HRP9WTZp91SbdOCQ325ZwDV7hOwxANWR9Gb7iYqC2aqzSVLa/L7tkJd+hrOHO8Se
FcI/iULZ6g9nnLnQ3wfwjh1vlgK042Tfdnu24OVU8f+o6O8o8uqUuRpnTovNj2vw
XOcT7FJ8YdhcfyV9jNUG3BNSQHuQ/pIrVRgIR1wQ9cSQ8y1GlfQkXL6ElPgxYP9E
Ns67uBH28t8U1WEJDrMbLGS3k9HZd4OcTGDJVWkL1sTxJsQa7sdplRqvAUGbN7Hp
rIhVUgrpjn/nqTFKu7bLFsbqdt9iejHRO3TgG0GAFhRLEpVmxnkQEodbCUSIUt+O
xTTwqYKm9exBym6hGF4EDNOR2ARFcUGKGA6SwJdsikShhRJJutLvVRzwoGgr00Ff
/cysWRQzisClvv2HmcPlN0WnE6PS5AuAXmdPmJf3Gqov4U6BxDKeqktYeHufpd22
Mo/zEqYhpZtwYyDRllNU63z3fjHC0nHPDgw7b/NRnqvYB9hGAzxwsg9C37o05wjs
kmr9w0v8+N/ToE454ffVsoJttKzi376ET+jgZWqzBktMeQRXM6Zuyb1EqdwLctSh
2HW6D9GtURiXPIdo8SARa4YvZ9C1s9cemTrZRMeyYUvxqAi2oHEb/bdZUfVkFaG8
cPYd2bPeHDvmXjFh95t9WZP+cdYQTeIAfC8LY7hcaspeLBDuZLI9KdHbxc7RvORY
I222UMl00JFq0NFIkEY7iCP5qadha0IlReoS8sDQVLQPt8UWUXBPi/0T8gbwYINd
4dIGihTIpmjlU0el00XszioAPk5Pzl1u6Byr9UGw8z6ZEQMnGVVEg6bjb508Eegn
616dUcIAkK7clQHcGa7rDaEzxuFgLCDGuKpSzEzsEBQ/NAVoUQA2thYasPt50MLh
R8ZHunEmJvMArwjktLjdNBgHmqdS+5+nkxto323uJ2YPpLQEKd8jVZm7tkNWVxNj
v1+F11U4+M6mmoMj6Vyevz39Mwsm+6QHp9i9LqI96oCVps6QO++bA1e8UESjyV7v
soYPAWzyMPAIC0Vij7syvCBvxTLq0gIiv2lNV1hgRupRRY4lEwdqufTQw8jWVBmZ
8iTlBt7ISpzS6rEoYKISqdFtxtYZc6wvCPAqWyfQ5uVrpiltXvc6MCJR0r/8qRmC
ard2YwheQfGIVhNqde0DW2IW36nuSdZfX/K22zRfsw1gKf9wcyvZs2SavtS5Y5FL
g9rl16WNNlYoVlinmzbTpeAtzhmCQ+r3fYNxBet/ieOh98jcpMXFoKUS5r2e3XNb
ICKWurbXEXjfxlt+FOAO63gLvE0yTY7HaVkEcZ8tQuBDsj1rxajCp0LWh9grFEt2
05UMr23Nb+VU1i9wM58DeK8XRnK0kSjNkt4su7xETyCw3pDVsTEc25OJG0AhhVDn
tuXm7n4+kmNX0llxyJQ3KSr45T69/hsAfHef9SDoaFKSC35kjPXqvaajzL6QbNXO
2UQFMBK5YXjllVxdrPKel6Ymzmu+E9W+rpspSnXSdmQt54RIoWNvEH1uJ9Zad1mR
+ZIlZ6AjeBZ1/qAgW+t5TSv1uP2WwODL121LEdT57At1jls6GNFf3lwD0DGmS/U2
ZNEivIbl5xR5vUEyoO5txkJX5tmv946Z+XADWq7k0z9jLMPghfOsHYgWq40qlWut
7gYzkQ3ung5uLucc3tHzUOANTM4byzTRxOnUCSpjdfjstOQcp6Nj/97gGzHvzzP7
LPeWUL8HPpYyUNwvCJ12RzV0z/JlPEuuvZ3kNgp7kUSZphd5DgwL8rU1HMekyboo
QfbhrrN0RXuaMBG1bd6TDUDAN/T5LiNyscx7l5Yi0ywMKYg/9i+d++kdi3V5NGOq
cKmQ0EacwlcjF45oSUKQEH5rKmtAKlIKKLjFh0z0mNREVRmv1x3MwjvyWexfZNU/
/y8R68gg11ua4/7Lz+P4QeHVdHrCqeRdYdgi98ZP8CKL/gemP7gROIUzLPFjEafq
8zenfkHLGadKXAcgsdnREJmn8CvyweKQCqbEzuIGnvrNVqOjj1OCL5AY3+Ni7jTq
UoFP4d169GYJjeVysT0b6eJVt2Qylrbx8Agnfaz0jdsCTRuwFgrjeiMEeNTG8pPs
v7/jCa1KtaT53ws/pK0HyN2r87OCWyZ6iWwjPx7Ec3FXNh6d4XAj6f2bOYsguzhG
H23zzlZsICWzrJlW4vhNESCBpYRNEGkVu7VskWwrQ8Sb4O5HcKWxFXGyRPXkSzSV
kjy5zHp6QH4B1R5JFJlG2Lo9I0WjlvewBN6RkwI5xzlHiQC2kQrpnstvCZy87KqX
TRjS51UMpr9XnB2NuzU17jihovMxBRSYL7NSABQu1secNgLXkKQuNmsKoWmJfytP
cZolky/39u6+cdJa+VG+eiBHUqYxLzyqE4vwX7FZevbuwqZlNZ5nj/W9Rg7Rnpi2
a4sVc4YseVZrLjCFT29pjPk2hQMIrcllR63Amucxf2NFxXqpki/gQaqwzqnEd3PL
TygPzkjfUT3694f5KPx9PCBYwfMlx8So157IvgsVbuZMbDPhp93WEW3tIUKxxQGS
eW5hpXWvoRBAJKrTOhN3EmDyainsMAi43XulD0m0H+Lgu3i8/TOY8TgfqD8CusKl
xO/gJoDT8O/rOIZjmzIo15lw/l/LDL8Cs1w74k59QrZuipY3/HbgDWP/tydKLoQN
BxNziucFTpYhocT2TaCTM+DvpcbSKg2MBzP6S92G+Nhp/3kigvZQLCdfQHKn5yrA
boOrClgV6SGAwDfA6a5MArvxsq/JasPEFtPv54e1sa+vpt+GmT3n39e3w86I2V3F
c0tKAB20oqRGPF3BGBBV8lPASH5jMk2CPoLBTuyuK6zty3BeDuT4Jl7hEKGCU9+t
Z0zyhJoRRo6P5IcJsKxgP1vxoxfSJksF+13BPy4UhQBbAgiQfTh2zSDh91+93QLH
PSuUcemahSE0vAbglsAlAB+V7OQxGzI5S/m8/GQ0Y12U5Sw4hIIo8bgSel2zfcB5
LfgDQzcRDlibL6/losxLIOXy3wKpcE7dUXt8qDUiXFd8Xug229YkoUmMINyBFzXs
4uN7T6ev0UxOicC4GuNnjyXcM3d2qCVFht9Qn96bVo9vptIgqPfkbMVhUXxObsdX
V0T9atbtsaYau1ouRa2frOa/aJZCnUS2t1vWS0QJCdJsIaZb2M2r9L+tROkwgFj0
autxrXZZolWGOH181+O/slY1zE5icotTEPKH+Ixb9pcUyFUU3fo3s4kYXdxb25LA
xz+7hqn9J8BQk+cXCpE951op+N/ictirB9TynTeuylGhK1JTPGOxUVFzEFzPkWvB
TvIqlq/6YfD07QXNRDgCfutks7oxL5zL9Jftr9foHLZHTQ84wR03Q2xz2T8y+hfS
WV7+z7I5yJmDIdrIhQg/+faej+Wnw+nIFt5zsgJc/OoUkd0PDY1Bm2QY88tdyLOA
X9xpaUejPi3rNj60PhvKMhiDVm2UtZclcySer6hMyLU3dhr1737sW/SjN7Qj8yG2
0uEUM4wTstDLomA0sYIuBI6YFea1924rQLBSxpVdncUbCwuPFg+TcagV/fU8I4af
l90X6A6WaTm5MKUj/tU4qMPIdn++XFOzKDOuIppJiePprpubKYNNEb0npVV9k2ia
/uNrl144+mFJDvcfUwFyZNNRCHmGWgJChM9bgwOy/Cc7Poaq0LHOW7H1RqN5jm6Z
S7IKPbmsu0Ugza1WfYvtLxkxhgjrFo+gSuBp+DRZAYiUWdh4sLeWptXDNIzpaeF7
jwkLq96tHgNl8LIZqhSFICCmCRvJ+hRvAUqDh2FRnD66v0LajtDQfOm4rsPTkq1a
+VOCA3Gl74MLc52NuQ4A2dqkZruwTaxjlduyXesn5mx9J/HGbuXpq7lJrHmg2GB6
aZdZVssFbgscTUhuH9DH+/QwFk1nwFw2sTYIrJeMXFFyLUEujUnapPTLSNID2CTV
OgCzkR2SslL2qTdp7Llf2unq0wPOWKop6gUUNFFumMCXm6+rhjRHWFmEk65O6M2R
hQ0zZtzDHrueXtkYrWEE3uYqL8fIxYUSUOJ/W3BNG3PUN0w0j/KAaElZpufrl48f
BLFCJciaaBUGxN4d1RDE4el6Xbicceu/6+JGhMNg09mIky8ph3wnALH6pf9RMpTe
qlHD9Oufkzi1G2lKh/4oWt2aKDgixUgsv0SUTkN2G+T9kioPrmB96OqVC/EmFMTr
7JuH4pgUlvxBquMyfcISKQsd3G7R4L+UpHdPj4n6Gc+JWb7cSn6tIw4NoHSAGhqJ
GMix/9PNjoPM41HQOMtqLhi4450o3EgSDDqQQ13oKMSg6zj+hDHd6IOvX+cggyKh
RRTCYeYAcSfHTjQGExC4HXCO+0O0YAmBlGCqdh4+4sKM4S5JpCdtVzrT8fmt4OcF
urKPiexkgXCDVqKn5XrAAYAeF2f5FKnBKOs36KadYwrseTTTG5vrvgI1gAKleC7P
jKM4F1WMZr5mCxBE1iexTX/RV4RGndFhRjZv72XEggq0ANXDUgK4Dv07NefCaP7q
bxEcv43O61s4g2CCxLd4FjcMaitJVtjg9LidtLLq6LdzUvR62+d5FyeAsw6JZhNZ
7Ycp2LdHurbah5Lozy8IGmNDslacvHb0UopnVIu7nOwHu/ALCJR3g5r/P5hnu0RA
Rw+PLuPmc/9FfsbgfJt4NOM6tWjwgAdn0H4zUc/QdxVIe+3mDihsjV5c7a5tW2ji
uwdjwGe0cFrWhxpnmkvFev8kZyhlXSVPmtRuY/MPESyi1yfXlFYQWKSoozndgMMx
XmqLJZ/GoTXuuz/lXGbz9/mbXlxDrqKpakVlgeI0A8j4Ze/+ZyOpknWDDsH7gA+C
LVgIfdA/768s39EjjHxzfuP2EfFriYmwINv0cZE4Y9PkdhpQHMg6675GkUzra/lI
EJ/pOKSCwKi6R6o0hurA0ARTG/aQTiy/EGQinNDdVu7dha8o7s3J3U4KMJ7M5o49
x0MTleTBX63z+HIR3AbXiCOrSoQ5GC4bd9K0mvZevISUHxNk6LiQH1Rng0mMfYry
61SVtYP+0ifsuMXoUKrIeN/gD0Md0lAZAImPQH4vVJsL3HyAnC9dWYcp0nBx6Dkr
JyJ3uZCsAbTsnDg0zzNY7xkODHKe1+0STA3K7Oegqwoxs667mvKQyYxdA37PUGZ0
FtdP76J7Dy5zvs0c/0NSXKcry8DineJaQybS+xuzZsupbaypHDnWWPkKa1x4ilg9
b3g5PDoh0LVjji7PuedZlU1HO95Lvuy2XWeGF8yNW6xALZZpfcFe5R+yhBC4opl5
tZXVljPZ3bVQP/a5XpXvbnFlSwOO2zlQbjofd8DxjKyLeLhTP6I7JbmfpLMWzCN2
dEu9p5+PTu0H3PbkAKegcYmS3yfO+UNEdoiFT1uzSumu35RjPA1eMZ1VXd4feSL6
V7tv5pj19uzoNWyi6Q/pMDzMCYXc/jp/ubC/C4mdu3un8BZzuJ+AyjNsXaN6JSqC
oSK50mbmsAgUUZ6rV6OWG9c5VHbxbgImTeXFvDb8GMMHtEIZIgW2NwNEo+X+m3be
dMLxF07zAwWLJEYf5OW6189FTPZ6JTsDzUsnrrlF/z+5Zwa9GpZKgiBYoO4W7o4s
Qy2G9AfCBX8h8tmw5rQJCcJto01LK2ZPQlgP0oDfWeWBgK8QP7mddrPvlDLTlnYK
ntxj7+LUfJGVlut2qKE3Emj/TDx2JS1FCuv+oyfzEcvhdaFwWZHmmTp8a5w943uR
h4SKfJRktWfe/xorfI/sw1OS92P+D/PLh7rvR6s+Xxtg8E5wSHFymKzS5n7Kj4fv
6CinN8JXweLVIGmuX29bHmKw0Y+RdbPHDqhzDylvhlG/eVCl7qenyakcJVv5DJSM
kL1dfZdTMejAItMIvPaPMx+Hmkz+dZUZ289kwLn8uTT86dC3s2/owuj0NqUZMNfb
xJmcjLQVRs10Hya4j3nmEOIkW7vzHDUYwXWPOKa1ExAeYwEn/QYt1yYvFs0VunMH
gJEB0/z1mXvotqdGEaEOfumWdQxlGT1Jj0y2mYg6In2700AHzl1sz0fobCllEzzr
smi6wL5eFizoxNuVLYuenQdCAxZBq31F7v46W9lg+vOpmO01irSyYvRhVWLwgdHq
Bw/Fv1VdGJ2d5spOakxYZJVfypGLXg2PHciYIgMyE91PjIfiEWuqYd+WRO4mDl+a
WXH7QPYS36fg20F/oiOzEMilPq/mdzHjl/dCiRXFVCgWaVZPpeu3c48dMhagJhcW
8zOp2zuGFCegtrsJBUL07ZJzEfrVZC2LpHYHfLWguqII6nD4N8G3ejB/sixyflp5
JplL5PFpqdCstrx6NIE/JB4lu8TjJFTRC3EWEWgnH2eXsTe8efSkr2MJOaxDWvyN
gcb23ZC5rz16j4uLmVUUoF3LWK08bQoI8D6ZNle/m2RdX7I6K/ZlXu60ifemFdFr
cSuYAhbCcjl9CaiXZ+Yrzn9UEpFp5HN018w+n2S+7qlp9PuljySDdBjLCDBKX+iV
dg7jyJ5LW1pMBqcqrIlLzx1EiKohAXr24aQecyc2asFCWHy9CagyPaqFGWqm62ix
nZFp270mz+DHS0VVmkeYGdXdz7+eKat7sajzXl0oLoAkeCFLaay4RE3R5LR0QGzy
x472FltjRkXvK8BKRftMDHif27ysbmjtABv+b0T3g14NeHoNQiU38apkRB5JqKHv
2Dzj/rTXTMw756BqmEKmeK+SHPuZkffSjNt1FQ16AiR7ogJc7h4fyX0wkNA/QRjC
YaRjV8bIizOhs947WyJg0NWbLfeIDpig3Ccl3PDjqoUUydQXjFnEAtupmITT21yY
rZS4D6Dx3GoF1SfbgNxNEyUvED43tQ93BIso8YwX8FqymZWKKPu0OP2JKmQlZdms
JiIEOOJl0B0SOGxXZwJQIleQ1aYRFHpyOmjFqw9cHv9DuR5xwfT3zCz5LleNPKZ0
hFt3MxSRzHCCOfQkcLVHBSsxcf0WCRPvZXIqJMeKOXDR+OmRX/JkIKC5HUEQJYQM
+187xRVlta1XaMey2U8W+4lu+1mzBNh9oJ092wjxJDmu359NjTGe1bneHEufMsVB
BHkNkQFZbJAqdFAhfWsWTdvKOvlJxcG2gh5rkQyYBK5Fypef4n5XXvchmpbEA6lQ
PRLc3GV9WAk1pu1PJ0MpPZg/zrhXkRUfB/ivr0eOuldj5X0JYTnJf33vdeKQU9ig
rUIzz74pia2iRlOIlNjrQ2DaF16L5oDr21UluPvKjtEtOc4Om4uBrw2hRs5bLIsD
7sRONSTxtfM1vKen4rQlDCdRaALSj8jIcM4OunTL2/LVzI/OyjLab8dnS8K4Mvx7
eevQRryJ5SO60P1mB4DuEkZ/GXQiik5G2SpUCfhqp3QnM+g2dSPNRFqhJB/cVG/g
Z2qf9z1xI9/VYmWyNwjR0NLNX3tIZMzoOO3XZ9Jwe/UpVAXBJfpWTeNBqKWXly4l
yfVZey/BstKYtxTzlWduNK7V6CIvyCiDP+VAllgIH2ArUCmEssC2ziFrUmg3nnSa
OQCXhDT95J2BDP5NqCUhzSjEvCI82Bx399laGQ0ZHXwU5ElDTf6FdwjNbbahR4fR
Ien3IN8RcZussF2kR/RwPruL3eiLnO+G8pb4srl+rPkjXe3yCHROWkp2LoKuMMuA
hQr8ZIfTkSPk6Hkl7Ld/S+vOYBtkY0m/peKVfJrtYUHhhuTZkuJqnU25Nqmd+TFf
r+apHV6TwTNDgxK0MGPRqxRu9O+yJzOC4dGDDiUyQ2GVK61I4rc1QmdfdZAefAD9
mwBNXzexZGWLAiWX+3hnVUjFkmTt7ZNsrzYZGSoHlG5IgsNxTH30IxhcZ9BjwHS5
Phg5WbAMKjrGwujDhcZHeFFVTjXvD/9O3fRvaJvp8/IjPgvXwweISv9fvOXjfJcS
Vr56bi9VhMzWJlHjnusc/+a1jfY9D6w2K0b97DJ+nUYEsqDnAq4PNbGcDe1bJPrl
NBULl2atp+ZBrssYARYuJm1Z1ZJewmxMm5c0gVFXdwd3oZjcw9NSmm0XRJCS9gnr
2hii3j4+F8ykobiTZ5DB3fTmmpyBkQY12ZpJ203iN4ZhOKUIab9IOg4HyRVhpg5D
d33lNpY0FkBFKv3jfGJS4ADJpfqLpKSjwdmwozsABkLBZKkpjq9uwlGvkCI1CAqO
Vn76JzWCMnJRTI3lYZWuRtY6k98IO2R1xrsqJKIWRJLListh3rdAOghSFbnZjKIi
BqlyodlIu2Db7Q7dQ0pJ9zd4rNP1iKo14iw2hh12WImJDWgNR+KT/I+GA30U6eL3
ocYuyGs8yFbH9mttw3D7z1xLsIyj/dGzji1AAQOrlNpHcA9TPY5PLj5lbF5/+s6H
s/KumGu/Pj715BYWgUA9RLv0r7QuB0+W/qNOojJ47JJQgdoBHc6R+OQEWDVDV6BK
hUmonBR4I2JCBt3yzpjhDbyY24KLAWA7XEUglWNdm+ll0YviA/nbsLXwx5qMyHFs
WNpknonPlbWm5EnK+CkyrwXQ/OStUlfn2H0JWWsXjUDJ6j+TW8+sfaooyepCkUSQ
ZeEYWlux6OnkY85GL/C6gpmRE4HIdUbxnYBg3AmH2ybSnhQoPxKRbgHLDRCAdFIR
ns4jyU5d1+c4HaQsGD7KSoSkZPZ2FW6vTUmOZl56sGwmqwImoWyqcfhneng3NoSI
VEFHjovgMZpH/fTgN+2goC8RN/qxg6AB4Q8eU6DJAJCVkHeJwxq6xHNH3NkE/wui
/6bJVy0z0vcWDIgKKvnrBLDF+5jzg0iSyAOzmncBbEDqMIlP7pxqM75t9eYYsWBu
WyojJZ+kt/ydXWvtwtjdulGlLfK5IUlv0ek0B1TIc+bk4MJheRgnTG3PZSF62QGz
CZKM/JXPOuR/BTFMQdhDgHq60AfOfofSOBgeClb2nnlaLh0kb9AtFcBWHhJQUbmR
CjzbgswAr6pTudJs87JEVq6NApa3SPPl70l6mmVBnoWzPpI24sa5+ZAt0co8Ywki
mWWRfSVZ73t0gL4yZ99VuhtX3pvRm6MxYUoeTQapkvOcisbHpwKFNwrZH2JwcBo3
DvqglNomzddkuCI2NJzFEAFcDNHc3wEwYqxSag777UNwyVPlJ3T/OvCcO/4WG+d0
ATG11wdP28NQguXje9hnEk3NF9MEUprDjbnlYaskSxnhASOE9VWcv3ezMAnXRdU0
XAG/8TRyFba5zITDOEShA+K6HNG1QJm6oHyW7DSIPRPi9XftOwisTeqXv3+SHjTP
xoVAzXrJexs2vysoTl0vp9UIF8LN7ny9jCP90tzfnFyDpC6f9/w1bVsdURNLv7go
8K2ymv91ibAE8bF+XOxqSm2T0VWyrd7KZL630GrjGbBMH4nSXkoMBrst85OIpgE4
bRDG5mdMiZr1wc9WzSbIdDIVGPx5ozVFGsYvEDl+OBXBFEhpgyAsa3UBBshRT5bX
MNPJVDG6jS5AQOstpAkBaN4LtHLysdJ82vciscaVu9SzvnngZdcNc30ZHThFKyZW
OZas+bLrdrGixuDkVko6tfnMDcTnHTlyPn4yBX5RFQs0RZ2jT1EwXIqxD4BzrT2W
/nFlxXWYQiPZIugP0ajk6Pmkjo3vYMmn86ikJE6iX+JKcB2tnMBvgiktlnIKdEZ9
kjx1nohTmCwgQkQ8MfKl0HdKK+d2JXVJpXQMyH4kWn0CidY8c75RwD8TCOvsvNfw
vTu1LxhAkoW40c7wedQc+5TGiYxJWaULWSlJeRLMfQa7967ORbmUv6WBe+evKrRP
+b51Riv/YY7AmYJyKHNpMMdUx15VNLx8SlGemBss2eoOBV5PvECDdvP4fTzYcJsh
B+wCl27xSUYt0W3sWhLGeF6AQSpGMYl0z41y/YVKPGM9bRwjw3duXG6I8kYP+KBC
koWQJz0crZNuxur7VCiT918ViQckQmyxpdExmB7a9bhq8BITME0JRFL0hEa0lTXE
+YpvvXxoxyS6YOcQdBhN/p164mGCRcHo2H5oDBc4j7NvLGRVNc/SHQOaMGVoaTxQ
nCEfxw7ph1jk1iyHh/hZ6UfldkINhmyZd1ZqZuUdeO53o4rTaHz5ZevVl2D9/cEs
+vZnZfG/ERPRUs/fkz4IEy+e91O3rzrWUroJokHx+Bn/nuG3856J6NR98lSapYAM
lY6X7BkBRrnpnrC/GZNdDYB/dyRC+J/eKUKy7besft+4f5vLyff9lFQFIMH4d6Mg
zgpyczWcF3ejQUm3T6TRmLgKsDX/50ff6DZ1WJlsqj/dVza1Ooza9ddzJzMt3KID
AU5GMLaWtGYOS9IJEkcj0tYIOXH/BwRkvgEDbBA8kqRKHg8aEROFPz5RkhaXd3HG
FzLga2QLgzDZGEe7J6sg4rLM6Gva0VpWwF0vuT+tYboU4kgYyxH7U5iHelhW6Z/5
QTFbYjwg1I0YqtEAokod19hLx2IjEEI51ytqKJldjahxEGUW0N8/RJmcKwiMZeJn
ffUNEaN3iz6+NZb/u9Pg+LKnTFOpGLd39q9yhAMxF9oCLdfuyT3/OsuGlP5ayAy7
jScBbGn8LwXFHf+Dv/JiQPf6pDDSPR8iEGbyhtl8MisGcx/p/Dq/49rsRPIEXBgA
P5bJjOA+eT4ju1vtm1f5StvW61XfPWo+MIhN+lnGzH8EXO0nIhKN1lCGTa8rbXKh
72FeDSXBGqsVgsUSIyd2uQkEtPs2mC2KpikFzj20o2cGrX8l/Jg55alNMg8sWwdU
iLTnlWcjtIXQXLcw5aLWWRE3CmG/nY8mHtmtZOV7N1r+aQe0Z2rpTzlqGZTYaDiS
TguGAM0/xlF2n32xIzKlILhWjEcg1D9daxemsgWyiWprFXE4JnMPqj9APQoYQ6gQ
kpPyTp3+MM6Y/GS1PO7vSn0+gXWcm6wb2wMWgdUR8RsSWqziLYdWMIRjQpvp8PyN
XuDMR72bwOlmdWXgzNmXU4A+pBQb4hgyZLzNQA3yUMVxbuaWpM7dF9qUv1nYSgdP
RFcGuoyoVAUTPcnO2El1dgGwHiFsW3pkvQgQjQG0EWUXaivsndWjnwT1K/twVQ9C
bw5DegBGcxd2m61HcTNAqIsMoMiYdv4UOadPM6Lz8wPzeWNZ664SxSgwhSjILbp1
PHSc03bNjHzb/fF7TJWCFD6E2kC/LC7fE3VHpgr5mkCIqsTPMBiNzkMTkNfHNdZt
J503eew+s+gzR+9Cx1DyqIryvm+RLp+UlrY+TvLTlOBj/EIm0rILBsLJC70nxWLE
ppzEySVeBI+RQWBJFHYLzEyaYwzC8xK0QcYyLdA6l/kA+peuI9R//XEQSR4oqhB6
t3uPB6/ch4emghOH41vwVJXCS7vHGBRwJLAmMYIEBI3EO+QybiKR/oef3ApxV4h1
o73veOaUcYQSE2gPdmfqSAFLTLiPOmCxSzWQKVlCdXxlD18QxNXmRvVxrBFAKTWi
YbCQFkO3ANc6M9d7G4ED/RYk0B+XPwcLXUJWv4sgNOp3OY45P3hnteI+Ij4THldd
89sgz9XMeSTAZbc7naDl9vIDzDeMvFqwbSuPKrqpamY+ZvzPhBalKKFkcOc7BNva
zlONFEl/8d3p0W4Yd8n8tXM3zd8fMU+xjDtmtKIXsR5vL3TV5/xerwMgwePIxHTK
EXt+C9RCJi/5VtRdX5UD6+lYtHPb4hL7etNQapzIPHFYm2DkT4oAlBo9fGFrGxby
4TmZldmM518fIQVeFE4QuaD8SiKVm1yv12LNdzg9ydFddJCb0xaxDn7LTvTB2bzl
dlJPKS22KJRthLSIZ1lkijuBYAxh0vZ2Swzl0K5kUu/yn3j6uRNjwXuZVbPVu3/E
C6sLD/cMF0cppa/8eZfU9mQkv57yphcyytEIoXZHBdVjP5k4wefE/WHrBy/3cvWA
Dii1wE5MFyLTf2eCLw8gVWbtOn+1nQfo6kIZQLY5zgard6KaSV6m5i/WkETuS2sU
KebIIWiOnVWnjtG6K/5EkHOHC+UGXxehhX9LtOmpStX/XdlK34zqXxBVDSGURtAo
MaS5RU7ufUHWwLpb3P7vrxwoP2eF88WLooojUdVnRmSpIFxYHmDVYF6UN585KNn0
X/ipbqNeMhzSINPjrC9qjfIaFWg8yPjJdp7sMwssoyAJssZeodVUJTnDs2hy+3EP
bUEsCiGZXq8Qdf1optJUe0Zp/GRCeJNHZpvyUGHC+OkPuwSZwUUk6TMoAsQENls1
xI8yN6GbD97wUXFT4zdBggwi3K3Q5LhQUHD00sCb34augKGvJK1+jPteQMqe4BTF
eMomWB2yWvLHcDCzMeKJHvp3S2dyBXBHW+acTrDixkW6ihmKfIWc6k307j0PnQgT
5P9GxOs1Cv2siQhr+TL8xe6hXJoLnYCxRM/BOvY9kUSYSeVMfEJw1etRs46yNqMB
iXURZvRmdA7Yk0CaWgEhCLYqu/yzuz/D4I5WQ78EZwjbNB8An6EpdPFhEy5IQcj0
4pheBaQTzPRY+0GH7FCvbcaab62tyDcV8obLP9cR4FwolDnJYPBJhDaOpZosEI1/
XADehjCoXPvVHqkHgp7Jvy1Wg3viIkZendHAjkhC8N/weBdLOFivvBe/y0rk5c76
Jm3DC3DGZUmoUlpTimvb6BXX5fkZ6M5MIWTksAVYNSLYeeekahAo28tpdZdNt7kg
MV/MOgQSP5ywO+zBk2jK65GrJ9npy/EtWAVIzWKz9bVy9Vh22DK4tzTpmL68bK2r
OR69DL/w1HbpfwOeBp6oMQhp0RKdIXwtYLGHShahHaQe3FZw3r7Wd0ICEZNpjECw
TCGFxCLD9C4oemsJ2J/zay4xolym0aJ/HFfh1xUy6yE57FxjeZSheUrW4TAcrtBS
r00UzTtR05Ew72gQ+cUvgklGlbZNmI5FEDSbIj7SoLyYuwzQUXb1Z+keKudWOI6e
hlNBZ1NnLZg21DmBmsWF2iJefCzGfjMqkoZYWy3jnVdsTG/4jpBHZVeZ078VgvYa
A6qT0CA8s/VjndXeYQPCP7WSp7QQEuxKtSMItU+ud24xFs4saqaJqg/cg0YIWH6K
vPBF8NSSdd7THY46dzTTBLvcJuN144Os9w/wN1ZJnimcHTyQvdb4fHQWqEGojv/T
Zp3+8VZU0xroAWl3Dm2TOYrKJBLUIiqarULdhNDvQwLw8wRh4pCxbslxF7G+B4Mq
LHzrnVdlD/Pa4DH9qb4V+/Oxa3CsMHQwufPdExdGodXdcl+br9hkzGgJBnC15qqQ
88lfzOA48YPHl/sk5zSfwfHmNtBF6wJSNqJPy5O1euzm/ZpH/HU05ullrfdUYqq+
YYXlsyGa65tLODV5S8KclJOyhkGbmOkDkJ+i7QGgHtH7TzDxpQ+Ji4DgUV3ItwHV
PnqBzbk8ExXGoncuyFum3qRNXhvaq8L+Zt+rIB/YHhC3Jqx87siuzO1CsNdsJXzN
VReEn+bfVuMB5XlXnrpfbVq3iXW/ETCcLSLYS7+pqdUzfsqSZDkRYlsJt5mX6TQs
eptFyfuUY7FlMlDx00Z4vBCRsw5P1g99M3SFdvNyRYW7zzFIWSfFLnWlP1p3VwwL
Z3Dw6EHKZXv8S8k/OnjFz6iRR5t56cZE/qT5DvpV8Cb1BovDat3Otd7ZNEgZAB0v
mOORHbcEJuRiUDfwPpDdfdUUMV6qJBD/RykIOuiZD8SHiFVSyFLRgCJaRD0Vn8Hh
2iudLMl5AJG6TbJdfTe+ZGzOZcdrS/wHPySRFMSaSPZLApxV0WXJavWRcTF28p/w
uflUrJFpUJNksfbVlN9H2scUSFkD5EvkDX9yzeQHeANpTZGPkiKU2Bn70S++CYIl
14z2zDEjIOEalMvNa89VxUSmAUOJtWlfXqT8HP+X/0OFvhQ42xxn20oFeYd8TyGW
bOxP1B3BkClfvYAMyc06CIp+llGKrzzf4Fg7mvCcVRWPkIYMOgoXjhQvSpWakzkk
9jhCXXETdLRiWsgyx5GtOcjvw9nkBy2B5DAJFnzBd9mwKrD4QPM+ncMgCqtbzeLe
4Vv7md3CEMWTkcoyAgY6TRFJ9n0KunYFDOdJBtG99Ci8T39V8Gf1wQ1bYUg53Oip
QwJJ1G07Qv1G/YYWU5Oc9cmD39zi7c9tBc2WRVBuCkznDCvJfacYruPjjGkdeNn+
yN9iDQkrAX/sN9hD7XAQyQz69Tz5af2pnyvM7N6627rEPyP6qlC+kScK8vZnYbGa
JjMttoXVd5vhh8zAOjTSnRecTR6l1ciF7BI9mP8FVPlu0HHJaxx1GbG1tL4yIYC4
WQ/zyQEa4tVy+u32YvOGdNMnbUbRkJ4XOP6yP1e5kSn8mt4VguOEavnSW3BaPLtC
tAAFdbaE8EqGmhFA2SzXYwQ2kbKgbl9sYxwe9t+7dB5HOsfucwM7XUU9co6eStL8
ou4xKtx8AM95w+njr2zYqHCWiSJN0+x+LvQjlWdo/wjkR7rWVfTdNkLZM9q7BnFO
18+0G90PIBqhiO+58I6Jl0/MVdAWJJ+b4N63VddyUvuuvUG90FMsFr5GCYoxyFQu
0lCxYaaZa37FOEhspV5DAI5BLYbqohJStDTLt7uDm9Yg+U2FNW5g7+coJ2Aa4lVF
YhOB9R6V/249dpPPP682toDwwde8/QahcflJoJYFNHUxgYGG2YcYVYbuYFL151fe
JWEphhqEhc1PWaBnGPCOVNm+CRtipr/aG1mAwAidKWJD8n3lho5wxToYEce0yOjI
HBy4O9IUypXZcyPOwP6ZSFSME7i11IlO95hM9c4L2H5D6r1lKqmnSgWXRfK7Rsdx
4yRzPYbXKF3fTOlezNVrWTrOlKn3y4f6LjNEb4A1s/cgiOFzNF6U55L1apLxaHtg
yU+kyW6tzztgSBZNCDiAbGvGsv4HFWRpfGiVk7MbMeCYfJmp5tlHGplQHqtQ7X2V
3VVGS3XqX4uzxttzEjh6+aqL59HlUPbWB0B+Ihcn39+AqI066lVjltl1wtrBLyLf
M2AQHlIR/jjovqfLaWK509C3uyUtyJJAov/i1lLxCqIwdWISEw1DmV/gm0itK6vy
57lSoHuQsdAKLSMLVlZ3mPZzx8iCdOCZknTs31cYi5O5LGtcfMwh+EajIn6uMyGt
b4bpkLrJElq/yGdz2JG23Qilvz7UwVBcZokxvHFLCEuqc9golz2huDELL/Ze/CSR
+PFN/E5xNK3RVPRW/rPowRdrvhz5fdq0Un6eKTWi5jVzA5BOZe4G0xCU3wxPeV26
gdYBOCDBqe0vDSy2XIYGfvkBylsz0tJsPS+NrJj52INlGBCcS4MQDhIPZqH3qk3H
o658IFQdKcfZY2s3fjx+iuBCP5SzVVBvD15mJzbTFhoBr+uhE39cJMgB0V7xXNeh
MJC9zp61ORQUjxMsbnuyRDJ4HC19Aqv4cbomd1N9hCxL0UrZoUaq0C0s4zV6UxOE
1yg/fywlZyVLN7wFHHx8ET3B+DG4Ydu99A9o6vic2EMZIGajKEpjWL10aqspO2EM
HGxLGRsM9F2RD5hv8PWDYa/Tl7gc68GE+G6MqsJFEHBlivrQLLUrA2kINEx6X4DW
Y+lzc4osrgKANlOLU8kEquZxAMI+j08+xCE2EIdEo3muTXVp8W1WMolfBrswbJSS
vAF3enJ5BziE8+tSS6/GvlOYY+MEnaZQFOgxjJnY91HxdBOkRjgzicPhwtKT5C/R
mvCTsP2DcH+w7EhduzrOcHCM7xxtTAHOglmL/exnvb3JHsTKe9/5CVNKx9UQQA0v
9X6NltqCd3DtdlZZzVdctFz7YIORGAn894Z4Y283dz/UdJF+Bv3ypdN3JIk/e8jw
BQ+PmzU6FxBPzn/Ctq1bh3GJcgtTNu8srU+xLXNSMUGJAPB8Wp8QNgA0SC8k3WYT
w3AtdHU9oaGwfeSkWRnWh71Buh5wTQLRT893eclsf/i+917iqZoH8NKWV8Dog0dr
uKvhhltlzwc6m1tdU0k+hETbDkZD2XSXIoE8SZTziDGR6Z+Nzrqg35mA3NaiYV44
vw1ALsz+GYsp/vjk9FU6HMOaVIXk6/J6Wmjv/LrNwjbFIE2uR0CphneGHnsVTMdo
X2dLOFi1fPQbMExHMUrvyxOllHNfSggA3VbElC+ylRjoodkrb4zBMZyzRiYXFT9L
DvDoM1pjXaZUj80LnRbgHBedX61Y7MCUdaeLI5ObJ8vFapj0J1Afwc4eD0+hr6Sz
IO5FKzqvsko36qxuLHZw6BNOlHT84WRfNESrWKGHyTGCbDgdGr0l2OTiARIfwzab
DmHhRRyBJ+d122JC88vJeEA6Gfcba7OXLwwr51aGb7M2b6gQaS0d7GQkM97ncRDQ
1YXGWaJR98AYe0JapfFI6QgDcHr01H+FhFm/ayEyhg0WBN7lIL/AL43TKU5WT+PZ
mR2dJS21oI7TM7j7rqCI2v5Y7yj29IGTKHWIBoMx/vDCLWgjkg6vEu+8R1l/LId2
xTPa7DwhM3lF9GSnD5PgnYvvWj7JY4eMJE6zHnRM6pdL0RPBq5llhurgz7KPJ2bH
HGmmhdFel6y8R92rzlewXVhPxcrsSPBgME7KlVwUBjwTXbKWeGZwgbODCuvrUPRw
BjEFUO9dqsA5OGI232P35QFADp6aag3eaqXjYqAUg7RVnL/EPmi+7j5WJdBI26uy
SkTAIxkY00V+KRuc71fAVzA8uD+obKcpzswNnQH0ZXrIjIaCBOcYBUbAC81XGjNt
Zzdt7CNhS2poYy3m0MwRIBIRvG90nRE8gXVc23RtXGdWMyuMVdaWA2vDi9pXyaYv
VNfC/1t25eMAs5uUjl99RKncKV2mWvhH3ZC0uaLCpu3DNR2L4rHX11Ljx9YOh1N1
rx4MWprZl8e2VE1rz5jOnurkclTF8ujlL7kCd6+OAyTSCvGe1sD1tCBEXwb7bJtC
ngIPWAutIwJEv2xJ6gMy0FF+QNYqzatlKOh25CLEggbLI4Vrt+wS50Bj0KHUejvz
/hfAr65h9XyfOSjqMzZFQN9/sNxRNwUsklYEWD7H73lv/aQHTdn2LeGv3IJoVoIE
mVp2eGd0ieQy0ZVGTPceDPqWTAGcU6ECS6y8LyGc7uQ3+firSOrFxAoIitQTNQB+
K7LfJpJTHseurgi/tEdclmZyOhCCPzEQWtsl50k64O7XJU83SJeSZ0t+nvvgFZ5B
ioybK5MFoWhrnRTi0QH2PUh6SRo2dpmYooOnZUpjLUmIXyrYjFiIjMatGfqvFcBh
kQ4kf1onU9TxejHjOGNKTfzruzPvHp0fpThMAaS0YnPue716SwjCYt/E3/0CKgOT
pedLDTklQz9tpqIccS4Hug8sgdBFpz0D3MCRKfgTWUsse/B2FCL0P48LZk3T2s0p
V/WCMw8DPtpQyWDZcL4qaNrV6n12yjgSdZZU+309wCbDf4B6jir15JgU35AbzEIr
nqTDcOYCjfxzj1m9V8Qa288Ehmvk3sCzHsd4nFfVCjYHPXSU+6nlHqYzz7uDk7zV
5VM4LRL0jAqkhPriGchfEQLyswYxKhdULgmyVagSSZ0cRQQPaLS9ULX3WEZdJ3Xl
nPMhntfbZYzMZ+YupGg1P37QdOsVj13fDjiG8DNAzStVkrL4SsG+rH96+mvNpkOo
okegilsQigw4WQK67uivTudrGsPMPMEF3+D3SdR1ABlG+0vopZHSB8+Ww3F5oY3L
sJvTciRkKFgvFWgdbbIeVPHBHrm5PaCTFDe60Xp+f9/yj/SIIJwbpRZCEJ2nx7Fi
E+LpFD38pfhZhFck9NOXuWg+lNAXl1VaLfs6KnyZw45Yu3DzTcWC6glNLbyxOKls
wcQUkKdvWUCS6dGcu/yIyaeJZ0vDWsWZI23S9xKLaZQv+1yubsEcU3JSz0iHCuax
kjx4RNFwogsyBSmmcWzwGY6meC27zU4loauhgpAs6IDpGUH29dW+lJY0ENa+JwgO
vqAzygKnFNaG8aPgXiD+gomgYH2Sw0n0zSaJ0MOrkEqxCcK/1nXVPWYS3qjos9CI
995QydmsvEER33iDbenziMktoNVpKsmnyoQMc+96eAkQucq/25qatp8MoTePfIhk
hFwRxpQ868oQq0YEaQzApj9HTiSIZmtJbO6JPjJNzBWxF08Sr90QlKQGIRCYM202
ZPK9FGaWXQuVElTZMM1jIwTgYd2vOXsAR7qjPmr2xnEffGoEx8qyc+pyQd01SIKh
iI+TNz3pJaGeP6eFTjKEDZY+cPXG2sjvJsVmNpHjXuT+qN2TJIPcqdXzUNwJFJhz
QRrl6RVyfubDarQMhukzVGu53BLsggRu5lYp7O09aZbxxjQpVQoJr/byAkdoPClD
pNfpQH95mRWJ6pvhYqP354K9L0US7L75Lmfwhhnx9DIjCqJCkFG9bQK7Sf5WNOxu
eKT8nwctsf0wVSdvYIP33A2bl9U5ZD/rqVPfNK9GDXVx2jK6qqnKzdxI2xc1cPyq
x6Iby77qjrU8l0m9evt4XbGbv4wwKNB0uDOz57agg2N8jaKu9g2BOeQeW/juMxRs
1sJk2YMZ7rTDrGPSbbKyRSWfkOVp2Ck6BCZV41XbqVG8Ylm4wiRvLlf1s8Bsq0RS
SSDXsTHgMU3cNCu4HoBlYj0GlWNtZh9Jq0s7k/jSSYKwRLPd8QnRJHiLuzCN87cl
XS8fhzeX0lfozfoXXaIdTJGU+KdM7AvnNYsr+ARxO98yQqrXZ1gRfavowDqlcDo5
WA+5kBRgtin5UOozwBqO8GsgPYO6ukGbxVjyeNz8wGIRMyeO96hhKpowZ2EsarVq
figffsMyhZnvDNbU73/TJfeo3p4LVh3JbW2Cpooa48GwNoiXPMFVLgYNFos4xcF8
Wgmz/XtPnRpTWf8Ru4nLs9myldnTLBVhuz8wshDevZLhdwTJG43pEjXwLr2e9lU6
YTL1diEY3XczYBy3OEBwHp3JFQ/JcKkgahyn8kl1/fcgaF4a6T9ohGXxfaRW91fs
XSqng2xsnuaGhJf1qkFmj+RuFm+335TfgKosqAddqMxz1L/SuiDwW26nZVwvkQxH
M8LVxiG4LH0hGXBDb17dYxN+CG4QfQ5woHt9aShEtwbOoaiy4onGAvyDmjrBbEqq
a6AdiZa2NAMXKnsiieVwHkOcGj3jW/yrgG+EqFYvUTqEcpHnCeAjOm/MjBzUcsUm
S+VnyBxMK0wgmIfDx4CEhR0lKzM+7KUpnxCa/XQi3X8y9iwtEySsmatnYXS3jroj
tjAUNLb6QHgnIWASB/9Rs5Adx2yPcWs0gPD74Lo3Z4vkbVIjQoNbWsEK7GELAXLK
EVagDbOCthh+gdWyugWTZv6CUBrUFSp6PkdByawnupV0Qw/HDmdXJ0sTNNBUpacG
Az5ryXbQGCvPvieuoEmvWYLtrRNIVt5ApiLJv8lM+B+eR5b74sHV0SACXFgnMFuD
6qZ8RJepFk7ZMFHo/NmDEnq/dlulizbayzvDMhN+iNkNSyWXHOhjZ5G9vOk5BJ3/
CQ7xqSFvqhFy6kzHoVg3S3YNvZH55PkvH4NYKfOd1JXZqr8MqVCHnE9clKrFHJ88
rDiifs8pDFA8uHIHU5FN9dKyAtSr1n3F1XY73c6VDv5bXl8UcqF3s8QXrnfWksM5
qH4dGmV3vSlJJMheB9Wxyl5p8UFLC/VVd6CiHtICfDEOFZqwlzB+xv9hJsEAsbAs
6Zy8VL9sRqd2MdinwicICAr1s7wrfrkgMmxqRmhAl1vie79C7S6v4vzNZTXCWuAL
1F5Rb7m6e0FA+FtAtM06RsMUdBuoATFckXPT1KQgpLEQs4Es6bxdD+8fxbBSPX90
KIFIVGlDXb/jsW2S/gNefhgxsppubkGewtiE/ad/TVMGnuF4u6/4oPMxv7olgtq8
O3PtIW5vHgXguIgY0mS48863G9vWOWAdcXtQVvjqCLnGG8m9S9fM+ckB1mfeek0K
NPI5cMTJ2yeW64fUYBbSYgP8AZpHUIv1gAcxDTFW2yuy/98sntyDpnLHsOIK4KaD
NG8HHsY9krgYyNzjut8TU7M0RmJDTDSpmhQiiZqoRZ+BvynqImpLUaWxTTvHMpZu
m7UjtTxHokUEzLQLTthI/4kq9CePpuzbZ2X/w5z/4VTPUNjlRqUic+43ckPu62FX
E7DXaXCykBbND1cTpbRPPW0joMUWUjIITsGPtQyffGS0PlzcY+Qmnlcs0kdU96Cp
9NPtpTICcSdOq1JP45780ULOdcBKRi8Bsz2fel1rbTcL9u4rnIYLs7/RUCPodr5k
2yoBjGAVOyPdsqMOtFBLY25vXWRocHzYZYCYTOYrnsb0/BaIVqEK8vLR077tqb5J
cTmRHkWzCJPcnALKRhzGztJ++xaLM9jRX8nYl+NPVmxvkIrl8Zk3yOv2doGJ63Tq
F5EM5Y65vzbKVzSwKwyqS3XljdSMTmanxcAbIIrAP7/W3HCQiSjnqYtvUfZM7LOv
TKPoXeGgpfKLkJv5paQENU22Gl43QsbXClp7NjGXSutC8G+iSMPNU/x9h0FvTFfm
9gd4GsIbPJ+w49sy0w9pfUPcLXBDC8KJCt/1PXhU1iUXtdQrXIlNhQxOlLOppmZi
jQoa6bElGAy7Wkr+kktrv7oyP1YlZecLyX60KNKHmgAIftz2Npr+7GzBvYs5DzD8
xmgptMxmRcVIGYoR+08iL/FA7xy9E2racCevB/T4FodK24wv7+0Be4hXr5nSqXVo
c6pXjyreKB6tj2YRiKVlVdO6f+QqMq5I4Hztak3pnunsiT/s7i0BwsPv5jD1xy33
VszNJeIqWnl1czuNWBFr7zgBMsX5UJxVg8HrhdIJvnN1KNVXsWpA8qSoRNKvpHKb
9zJagjKTWgTVYAm3AOLPG6Vac7wUtzsS2XfPd2O++RFAJSIgE1JmvMz70xIaIsSU
fCNBnqLBb8/jklBk7yG6vlciGYS3Ze51ALUSWbkJqYVAwl0fc3BCOp5rZBVWKXuq
XdP0FmgueFbG/2K5uvP3sXQOM36jFmcpwkFWe5cZ1Gpu7qUboY8SfnSipCxMzHy9
ATyu6bCOK7vEFWMW9aznkJhDt98+OZVf2qMyPh7L7+tcEqRyfr4Ufz8C527/po+W
7Sx+m49earBSN2vBf1QktASomVlpvgyO4W04+ikqBNKSmGJ7qVuXc5NfnRFs8YTa
PHV6h93Sb/60c8exA5IqgMDUQ2lTeO4yjna1xqYWF10JRnF3DbrkI1DmT2M05P8h
VOKeurUKTeHZQ9kQBFtXdU5aprVfWRvdutzbEWfjnDM/gHLF4hzlR2E6AD8y2p6T
PYBQVf4eANFGGun+Oadk+jZSaH3bBvc7FnQBeEKFxA93wp07l+3coZr2ziwPlIon
6kAkaFsM/3T0OXDkuWnopc4qFnFtnu6BYSPnqydBKHv5aCi4AqZaqiE0MPWTrkA/
DAHkwIviKTVe+8t+vRRbw+rv7LpyQyZAtLri/jbCw/vk9yrmAb6yS8k4eNIGs7eu
fYGR8yKr0NQgXvQMzwKbAK5li0/IhG0g/qGJ3xc/DjJc3wUN/HK0RbQU1tTOIHFR
W0hVCR9V2Rn7xf49JKcNH1BBiRLupKqXc7rtLraeiO1uy+l84BGQPCxPJPDqkjyH
2A96KzHC1Yzd2K9eWdxuc0+dbuCJEgP284SWo4AxEBPPdYJMRuClq9AS8q+BtMsf
lMeq69U1MiOSFaQUQd8/O/OO5lfpwvV5AIw4MjyRuwqQ2+b/WLHuQ99br7Fg/AdQ
TGGLD9+hWUEaCqmUPtx0R77hLVmppgU2KdwF7n+qUzu/jJ5PTuoQnijSjb+u3Sua
Jwk+vQtjDIWFh/GDrGkl0vDEwxdD/GSWKLsquQYmZqXEt5OzwwJDmfWjRcXhM+7P
bwwDDUjC1LlXpT8DXUeM+CGQtXbxfhUaIwD9OH22Uo45oXL1PmxEVVKgCzetSmNY
MI5hnl8bnyUOZN6M2AAJyvIAcR6XnEJTH2aRNyJEHwnUZof2R/JJWcd0IigPWxq1
FcbjGJ2dyU33GM/nk3qsd5cRSNMBoElV2chcnhL1Fvmbl4H/V0L3i1IfdMloOwhc
ATMGrKuP6eS/lLj54o54qnWtzbQfMdpwpeEhTeqzowZo5fm0PW1d9SZFWhazlwqR
nHLjP0sA0n6ahsrqzeuhkZ2domTLtyn3ibz8hDn/FGEy1IYBDyGb+LpAYAyYjHqu
SoszZk8Y0x5nQqlhxpGywRSltRrYvDOxPv3L+d/dxDvhTxvsaIjo1Oq/yTJBqUAU
CF9m0OFXL6Sbw1lYzMu/cyxwmCg+IhDwa22UEm2Km3mN8EtmiZw/3ILKeD7fugOy
z+dpt4w1N2pycnV8Zn4qgHArsQk2bePAFnriCRvLyffAvyHzMeesVmvjKTl8j6wQ
VoeFSTT/XtVVe5CZDsLcMIf/sES1sa+FcB1MG0u6KVZ1breMYUgwdKktbov8KxEG
18c88RVRUlmUvwQye9M5cjgOfoYbv5QIrx5QodzaJyDE1wRJejmh1C3AGoIvzFQN
4V63NBGSHCA3RARNsdKCB/XkJS70hnzJOb468dLfb+CYwmjD13hpO4JcIxORtJ8W
5Zz6HRjzm3H28EFiCdb48GnV0PoYMj3R5uO9lKzowIVWpjdXcLeWM82aOVLMYb+W
qbwMhxG2DGup52TlJavp9qvtRaezM6xKVItgWcIivVD7ux9avA8Wqa9IL3mx8K44
qSLP847mNi8A9oh0nMX9KRc1Bh4lVeY1Fu2K3D72cI2ewD3oiWcsLlJ99QnSD7a2
VNVV8XHK5Ef7RDjtXkY5yTxbfMv/Pit5Nb4XX3CG+QpkLCZoCVfzW2hBg6iUVH9z
ssPIytsPkkONJeLFMZRtGRDbmK2aszezRPZCKaUt0gKIIkNmMWleoJ21cC2092NR
gG1NuwLLOR35wNQPe5oPLYks2F0zRsyhxiXSqyVrt9WTYqvXqvPfYZ1kCJO28xZY
sR16oz+4ejxYHoSMcdx1KkKllFzm1IYuOs6LW6sA8phJMRgWDKLB4F2GLLfIk6gy
E31W1sqpOxQxJ0rDJkY8+wURlN1vhrpa0V+3JJIA44I5MRxz+PcwB8dbNI9jqfkB
Gj+mYtDFyDhcv8beLytcJjtthgUQuoaydE8ZblSwsoa+zxEyclsN75Wf126SdEN7
jR211SVnR9QCNKp/E8JNEVGXW9bRuFXXksIZewccTiqhW0JGwobAPL3v2n7twykz
ZYsrmdfUwBgoiDbiaQanOZwQPf9K1TE9jnJmNbOko41H6zapR4r3VWVmfYGHVh1a
NJA4UOYYaeb7qL+HFB5TOicGd51wawgYphxox7pGMn+xeAV4hvP1QEo7zEnMEHAn
oeEUGCM2Dqn1KlfFK1Myd5aWWzyc+VGpsezwDS7/L70BqxELtkxXgCSscho9HNyM
t5VqrrnR4F43cPjO1xvnYhIdh/xfTBda94YdhxYRYSgxH0aWMSUeAn0TxTlfczg1
4+j1YmRLhgKLL0Awfz4KaNrvc+bZ09Np/9doKkAUu1B/+gRzFbvKAvwVN0pvzGjI
zviYkL7epwtrzuiTGPGCdAOmFJhTps8F9eX+glznoMSgYGr8DJYfwVfz1SdqdEvc
1HHgrStkPLvjUyFGCfLF4XyJBu4I1MIr7sxUr+XYZ98ppdhL7W0c+gYcanaGi8ps
trI8tZ/joRby15/xjPQzF5hCAnDLPa0qOuCuZYpYMHfX3zLGqLMm7fu5FZb+f0PR
v+fXdccKa73nNr7xaXr562B+5cwuiQPext9zNccW9SF1KCqKgljXj4LtcJ9oSED+
4v0+NglkEdWrrK/CL4ujD5tOa+EC6sJg0Z+Dl28OMQQpEkutf1xeIJdcKSnE9OrR
BwFYRCcsa2dR6MK+pRhVrkok4Xpl6NazsqW4FDPXIs0tq+xI2DrJrF8/A8uTRGJZ
UXHfsDnoHnd22ntyBjY6W6VGhxmFO8nyEjX0eNK3lIpPB88bRlLcn5Cxh3b9QetY
t7RxJkgqJ2t+0RIBRdLGStGd/4IdQbtAe9IgDdZPLvKPyVnFHQpklh2cndS2zvBh
wKlLyrX6tyOLBkwyHjThQH89ZC6GepWmCA6DXzwSmuyLpiFN4nTZmcvYIw9HqV34
d45p/c5oOCgaQBi04t9uA377eJjwih9sDYYzpFcXka7cIiCU5IO0ozl9WE9BEULT
u5NRcVCuLC2HEyJoAciZHqdLCPOwxzuvW67z7q6Iy+ITxvgVe1lTUsIQBwJchZo9
b7smJjxwF2cqs8qCmboWGSB2AOvIa9sUlKY+8BN+eQniTKbevwI0kF8VZm7WtaFS
EbJ2OfvEC3H3Bb/PFaMqoiKnM2tX+61qVJWx938Hhv/x4Th3ACcf3jLbDjH9tGJk
E5A0SGe7VncN5Kgu5dR1KC7Sn+rYPTII0nkcc9xHZzcAppYyuuiHGZIBVSryYTQo
MLZaKXyxwrv+/O2Nl+C5j3SZVcALPI/ZrF5/6oF3A/drP9X7GlxzRKCzhwXB/hHc
dwxUzzfSH+f+qP29Mdpo2N8Gs3luvEMQwGBz2W1eCdPzvYLC1WrOAqWajgSa6Xot
3F8Q7wjhGQA7Q6y2g+nyGWFfqbHdMx3Cc4FFCo7fhrSZdujru5jPQLrdzq7Yiywc
cRhgODQZmQ2P9g8JW+ThrCzLBrpC9eNBb15VC2VGmpXbir+oxjBOBHuG7G0zk3D1
QoCd4n5r8sPWW7Fw/QqTtbJYzskS2KXuGom0TxroYQyIJtOzoHiuzI2ELsPA9Omw
N3YasGWCk+jBSqGoccTwjlRaNgzAYrNsJ4RslpBB1Grb8sv/Yqx8mSXn7cYNmkUI
QNPiS14j5Dkb2S+QvpeUoXMjOdsAaHb0pZO5qc0TcC5g4ssCUI5DdwjWxpZ7mU7V
5Fn+MDhoGEvJ+luvr4F0BoBjH7jWvfsGDQtBmLkbKio7O2jQxbSyd7QGPqM3hrOT
Jb5+pgE/a8fg0C+bl8vnR/oEEZ4pVKXTb9yZefX/azXROzZHCQrjBbfZARPl2Avf
XyMvf95WRVmsklZMhEehEct5QsEeIk5cMWcRCVmOLWt5FHHn0IT0Ho+svF0vOLbO
C2RAFAOL5W1Thsux45ZS2sT4roX5EnadTGKVlepFYUWyAukNdOOPyPVpwpSeGfb9
FguCI4ygfyBmYvteYbdeyyOHm1LIPfC0jahhUzfX1BDONOmdBMn8JS+bvtDnW+dR
MfuPHGAY4kj2oNJWwYwns8sW3MMCm3gGmsOtEsqfcNROxs3V2F60czUAQC3oVqXW
BUHwLz3t2iec5DexqI78jgqvQxGsBEOhsJPNIqoNwZ1tzFX8bPvTDaHhoPXY22E/
GooFEvMrsPZqQHTVOiN559Gsv353wGoWdGHYbza/ZUMkbd8m2/vwwWtTYp2Jr2pl
0OFVH54Ef1T8f2U8fgyW5g+6NPd91RHy4O84X+dE743R6poNqGRE6it2jKRFmUUi
LOHoKYpydi6Cx+H+bXsQ1gBcvJV8Ztt2G7+NZF9x1khbaM7/ufhwqtPLPMpOOYgO
psMOhiCMrH6jPtMRJpPKJubuseeBKvpcxO3XxNbz14sIdV3IHpkSTXJuyC4BqOx+
/k+EndufeJI3SBlUvL2eoL0reKmw93g1VnTJREMWOqNn82gaFESM8CFc3dgOuJhn
BKOPcYw+82ZZwG0FPz5M7LbgiD27B6ffsPGsoFZhRfctbrHYWcAH/Bl47MoN5Id8
rs0NCIF8NsJjWL0QITk0ZYsoEfSJ7EJSLTjGBCU94bW4qVnlJEST4X1VoQ76r7Zp
GfmGerb5MJtsQrvcnwfQLgvGYI5c8GpKjwAsZ8mxiWfbnc9tNYjHiz+Dovzk/VUz
Q91Hw5Tyr7LntWrERqSPNQ8P8QzW4+0zeUV5KCeZakgM8GcnaaFiqsG60U90OOn1
Dr2Lg/PHLoxKKE9Fb8K5KjANX3y3YwUGW7tyAzXR06F15aKesrR4HcVl5l6l6Onu
TNbG/gQdBWWFoTWt4JwJVmBhSL1Ohle7cfL6fn+q259caNtHJZNLMwRdjExwDdOY
v9/lXshJq54TfoEyLEA5lRMDQb3ZQIcYUPaSVTKntUGAAMRdnGoXBuVqrls7aJbc
YZiQOLcKp/06EgTbgq/hSlTlWHTu1m6lHyNgNc2jCDrUN1YVLngCeRD316Vx2Ucz
3TYSJ7tSN7cc+yz1rfjFUArlRjO5lTIK2O/7Tw/GIEMLpyqKDX08JkMgPvMQ9jHG
5G2tKdwsik5psKWwO4NtBLrwDTExJ26xgJlaLPdNuxSd6+2S6QCr4UYKsnG+A4Zn
IZ/rHNly9hqRKsZmLL6185jewPTvAfZXZmOU6IphnUe1lLfckHQLwi6H5ElxZoee
4RohAuNl16Nc0NXo7z1J02GZefuSvGUpG0SaZBrmHTDDmPCUpBAyyFlypKeWi92L
y/Jh+AKkrUqc+WDg9bzgEQM8izAqJc4u5u/U5dbv5avQghBop7oBPa91oPL+eWab
n0OYqA/4QOklk4Og2JV8spFhY3LYTfr0/X/5tJBH1OjZnNsWX09CC/KoUoKrEl0w
P+TMrrzR+EZEatJH1QdevklFbJ5S7qtva1eqmRYmBdVsRGy+w7jxCO+Z4+XuA6iA
fzStd4A5f8lEDor6S97mOkrLxUPxAmnusf7Fq5DrOoKwguLDb3PsDYWY9BcPTK0Z
QW48CmTiH7AN1uf68yMzpdKf3zF35ErG1t/MNOlGrlnXLiBYc4HdZMIwH6/rnW5h
H/bjtSy6ZRBBMxN07X8vXj3ZHnO4pBBt9o+4qd/PHi6wycXMOagafc+Qf4kqEFXV
4qhJuVlDCZQFFt0a21AYluSPkOqv1r+GEkV5/f9UQXx2lZ3TdJFYIA6pL6EuxWUH
XXSTBY5XWsPgeEuThevxazCSiFDdfMrctjp/Ca0MCz8sB956+gMvlaX5upaYBDWk
1ZnM4uYenX680wuFtCDjohfwn7nz7llk0swRIgN7xHrXK4Eb5mVi8GKE0pcVgz4v
8KNL9yEpuyJ7INZePAh3awG+oy7dmX/LFGAE/iXDLzcTii+TNkTj6QTAjcq0+KRz
jVGxbgrLMdMwzQMNA5uwVLjws8KNujjWwzvkFSmnGVFIp+2SbGHZgwRKZed8rcC9
VR4So6s4sY4lCyFMzTAXFkk3BaTtLWmzv5aTHtKjvhU/1W7Xe1LxknJBo8NIj/q5
0DEKuBhGrb/RC6bkKSEkhz1rx0NU9OdHveOEbgEeouz6u+53IyHKxdwTtG9VEMci
YwgEjRPJtfGfNZIRnmSQbrMBpd0cVBJ4tyxFbIlc/lSSBKFxNTQlP5J6ATG2IzwA
15SvOkvaOhdxRN2+WfAWcOEtDgE+XgOkwpBfrc0YL36jfkxd2zRfKO7sS+WbMRXC
YtfidvAX+6xtinp5hWVF+pVt711YT06d+id0wk9P8Zcz+D9el+b62XExzbXtNgUy
NGb4JuHjfFvoldkedUoYGL15OouoFYvCTNgaAbX8iYzrVVqoBsx7OIDOUxKr/lGM
B38GgWTDBUBQiKs3OWxSSXKm2FtU4W5oK1/V6RorCJq4Bfp5NnlOYtVt4zSUyYuL
Hfiw09xb6Iux4T+8jThTtQfrUXQPqnzLhIvF4aJT5/7rerbFipm/eq+2uoIj6r9U
ZEr703tmh8EqhkYoVcKq46wDAHO/6vtr/U3ips6c0fBnZk6oslsl1zLabLvjtkR/
uErAsPkE8bLE8qMjdk3H873fvYPTwNwNh8ffePloc43WVAi8Dv2LwR4nIx41Ywgl
EtZZpPuILLUQwMbKMeJMlEKJcIR15gZ21b8RStlNUDHJ62siTDSoQ9rL88UDfHls
uXqrAwOlpn0nXPqnnr6FQTpYD3HZmDuWeUw4H5s/Uzp8HWavL22JfNR30t1Ol7Au
7XTDTxU/4tOwwII0zU7INZWesEr4KNVcqNwJm59OwEg//0BOxvkMQt6S25b06UHw
FjrZcLkI0gqT+hII9XiAwZViqEHzgnGw0YAVn98bP0yEidvkWTONQnsk8x9s0UGX
09JumCp4Bgux8BSO8irVAvCRDcFA9ndaH3pVAH/4hcO1t/jE8onDcTfgWCGIzqk/
QWYokHSS7sfeaxco8F5BVt34BDOCPGVtUnNkHVjcybkWtgItBY20zCuTyYkrq1gR
jZiUAuEuNygOA6UZFKTiFXzd5oXFtiibZRN7woxAj9w35mTNPfCbzEj+yoVbTWS3
qlYdKgkGUeBKzC7EGTfuzluAs7BjCs1n/uLE/2szoSpWARA34F8Eps5GIKPt5SxQ
PnsqveI0Y3t3hWhYWZaat7EezLQGmahiH3eWSpUN+3EGDSuHnGG3FTN4A1bWIqtA
vqHSM31PQ6vmZ7nmZgyU6H1EY4Eo4G18M6eVx1omOFgzlBpa/+BFXtmkzeP5WfWk
/gXlWD6xTPF++h2oTFhHDiJ8hYA6scxcLFqhpuis7ZIcg1ciDhdpoeLrNbO+kImT
+2fA5bRdHaf80TVwlYo6wsv+NEKNp0FR/OahGqy+8q52C4cTCJbZ28FNQqwKOwXF
XCrpambNPDiNbDLm4Vg8Ry1BREib60wRtvLjOIC6hFfeyAUVQ8JuCV63HRgtZduK
/7e0yjGB/XDWnNFdxKcd84D4izh9JVmCDDRaTWJpqQy9m+CLFZoVzRpNSXEkBvoz
qDeiZTEyCuW+kPetj9ZVaP+SSPfBJMpMUAVT2STN0ueZBm8c6PeVoVEtXWoIcaP2
NxcPQn+f/tRh1iQjHda/a3p17Cf8L9NhYV0e5ffjFtamG3SNpv7R59rd+0NOfnFi
sHMR6SEzA9yOgo7uvDzWR4RRIFCmsq7belpg6B1fgr7+chdFbcFU4RnvW3afn7Fa
vKWtYg9+YhZwLskfz8wTXYKNW4JfgScuNabzYDmKpC8UOHxaOLMS8lGTTgAGBjkm
vIrrj/qYptnlso7IQ144+pHh371uW929JMcuTstu9+rN+FP6FzyI14L+fTLQlG07
MiNmfkExr5Yb7KqR38IE6MzijOByd29iCMzVcyeerlwCxj8/ye5qRvcrfvcSqX5o
glgvKIE+KOwBe99OnCLTxeACVs49s9X85pxu9D9K9KV7v9BO7MvA4ONjezNpDuRv
TJw4A/EQvQe+YeF5tZ0wtEcLPwUjRC/I2F/D2DkzX7K2LPn9OxfbV2djLNIoSBiq
Dr9DXO8pDvMTJDvEqv9ZUcQD95xeMQYB/ngW+cijsQ1IunaifY2DaTOn5CSqHnVp
DnNVZ3pU2Qa5NIFeDp4rPZwSN9QyyxEp81a6hPddAedCSFes0HW56OM3JW3EhK/D
8eVVcMI6nybGKGYQKfixHNIOSDPr5um4B2mh+2yTft232bU8/jKjDGoh8EfqANGL
azPniHatadkOLZIXs31qGmILcjjUltJIvSTHycjjsMv02jkEa6S0mBTDr0X48Ziy
J7dC4GRPa2Nt8F5VWKblkXUXPODDmtv0aUOyTFkXQbWHgL5d7dj6sChnHlNv9g5t
OkuM0MPywaxEiKvBWu2F6yMgtGYbM86PO8YrvE0oXyP/jxW5AL/7qX/aiILDbF0M
qteZBQPHAoxQ+EA98X9X1whXra06JKA6pS4oWQU0FshEESFJiuKy8RzRA38J9sCt
ETig3ikVJ/rHC/ibdjd+xnTFAadhnRfKfbSiGsSgrzlc7I6WU1KD2SVQMZVVhcdO
mQakZzpEWRkeiz//UdE5TbFp0nIurFCeETjm3qFoWurIELtUyIT/5rf8HdIKB4mi
4U+eRi9Ix6Kg/W6XV2P1njQzOOXsMNSwrxI7Kl8jUwYuDDp/WNwfuCVrRDJWVy95
WljXQrCPsMO4qhZgpFarNQsvUb5F6MKVxRQK3c7jZCueENv4ATj1XieU3bM/Z5Fo
iG01EtJEeJIBCYBRONcZZxrzVucthn6sDqkSI9Qp5AkYBccozoOOm06r53MuvhEB
M8QKSEFOBYk0nVKNVbbFg4ifhbDRuLYzlL4Tgid/KdFfpQgXTZfOpV0tYQ/n7/HW
R9Nfl5L1VEow36PHtCrqz0oV3m/Zc+sGyQQcDygR7JhNBYWxdnUHrRnBGyaDYmTC
AJUDDnTIkjNV2yjb5miqnk91nYPxMnhWNF8sVGPh9rf75XR1fosuzT+PofONBiTc
GgU+5ZE2FUJwlMfuh9ehyaS33thmbemq2d68HvDL0OQBkk0g4eJIAqcLsPxi7k/3
ec32H1jp8EBsYzNtjnIYCoxFIoKO6Oyv8XBLD+pPCj3BTWvK2gWJgWUCYH5flelr
OtVpbXy7h1uNcxtle8btinhQs+pNB+0+17cwGLtMhXBUDtNGrox7XKLYxjIuTxfJ
PZwsO1C+hm7otf0/4qX+L89yA0i/sC0blhrf8y0t5snA7ceKpNVY+YIjYdapRJ6W
l2pej4AoqsOKY4bhKf7IoG0wKttJ/UMuGjTtfzpNMEVlzjcE7uBvVI7uwoVaKGlH
DqhYQaX6V9jJYuFC9LyVGrcM3NH8YCjYeMLwm10Ez03rWF2IvS5Mt5oxVlajfSaA
ob3tItkNQaogz5Lb/JUq6SdnmCJrszM5HI2PvgzLnBixKCl5L18kOyqWdEn3CwdU
/tr0fgFKmRSblWuoeEgGIVS8C7VC84QIk3XcXz1e7Qx1t+lGVhgRPX0PPoGVyfin
rg/QCjQ0r1wH/EtMxEcdP/syXjUBpsuYQYrIRfuQzc3oFCltqzQ9ABKpD9Mxslla
aCmbVEGcgtOVizWr5wvcpP41W8j5flsXAV06ykU/YfrkOWhpN09hMdpl+3xE15nj
Cyhq7WnJdl/2TCPNW/JjO3Y73xMj9OPdxpkPSHdU2lZb7mBZe9pGupoGiWXQzMa8
CdMBDBSbmi2dmOOqDj0ZfuUd5lCBakPRiS/h+SHIzvT2/iCGU3xBcGbvtAK8ttiU
mHRwqK45EvQDoNfo2vpiUQx5Njhj0RseK5cIgXfy2ihX4GncxTeSEmPbTpIPoELd
KPje+3lxn3b1oUi/wRrfgSY1zHzCeAgx1rAP8P9UdudB7jlsZb0oqkl9lyqtwb+H
LzJnVna8EmO9FvxvlIwpN51gt/5dz1SHTQ+eflX3t5Id50bxMKerHpWhYw+QdLPN
vC95palMxP7OqGcGMFvIIHqtN7Txf30DvoHHbT7giaa5inKLPVMXgZ4Bbpr8Qf7W
uKa9BilzEl+3BiGxXfZ8hrbqfbLV0nl1HXzGJ5by+FhL1lJ2sxEOvcC+gKOjl1Gr
PTVRVgWfScpMZXwtil99YZJ2F1Xpxiarmk/QbYt9Te34SS1QnAS5Ew7aPh+sNNCF
mBSbTxB2DTnjvjdBCQa163aukGktCx0MAMSZ+ToJsz+tvt34m4rwMwOzjN9f5vnu
jyhznUY6lWx6x5O0Pycw/P3ngcryMgKBaPS9bnaQkk8aLZmDP02hgp4arf4JYvWW
8byDIHlzL5Ga5DQFWQ7F3Ae9Tij9dO8kSyj1IEt/KD2ij63J86+v8gxGJc/i0fYK
bYYXduDyGPiah6OmZoaelOVDo/Yj5AFT0eS6sw5SGpg7UmDvGjJqAOO/67uV/Frw
r42GpD5VeOb0fZcPmYrLubI40JzZ/ee7HHYAjSH6BO3CFmPpwxPRHR1QSnc82PJ4
dE8nKkqBaJ4Tgx1TLBvanHZLTiXPH1B4lMNVUVGQATdi1ag0pABMeoo7hB1pulrC
PuzAz+g+B1TIST3tFnKKfPbLWq2Z/n2JHZyORIlwgldwTWNhhzF8sOaOldu/A3NG
rtbcXjyL6rFmnjTxOvCKNGxfHwoyDZYrkENvXLZLxYBXUua++2R6n0ObHRxhJVNN
C4Mm5RMRLLiL/0vLnEvVszx/hi8RFTjW82w6Neb5l/Ka4AwFJPZygE3r/SsIe59x
0U0CRT9Ek1QKDFgSC1xA4Sf71AjqMym+f8jRIGpOXX4/j/hMIa4FCHGxSdwqHJtH
xIJX8CJkup7C08Su3sKsVcIs3Iyt41fBhafOU0jOBJJFLMa+DvVowX3f5mzgPpAO
9cnJl/VaMxHUa6MpqpQwUHi/Cp/ZwEOtQ3NAAWRu0MAWDfASIyDYFCLQvh7cSrl8
njw88xlwigU6gxTXdDLyJIbNgilia0+7gyQnueS0Fg0Qura/ONJ20q1+KXGlGHdw
/T68BkfTQz3Ni6Fjloif00W40Fa6UmKRLg0asFSkZjTG1x1o8w/Wwma/xLg426wC
31ks8VpgB/EA+c/7ByYikIOigEdpZkFxZODpa03LCttoBNgquELGRFeKIdXNnRUb
7GY/s2RFnD/Px2LpbaiyEyHqd+/ED+3Uzu78oPDJB4ANuk/J6e2ZceciUKEYomQw
jgSzhzPOB0waVg5KY33cBBv3rCJB/a8IvFp7RbE+PDz/CtdueHvA/eI3o6goVzh2
t2NpIJr1pEoNG1aAnoQfOrpNCzj7SMtQgvElohc6fgY6ky54eoXvf1H6J6Cemv9d
JYTuSqQ6RqjkOWy1vcfDUYUH+gCmObTFUbx8VxYsOrRjqO5JXq9HHbllSRvWsMZ2
JSXw/0uNW4A8tcV+eYj/edFrjkez/HZBfdXpW0URIBkeAgGzRZdUJn35cv5ABKcc
i9XojpFYptdRyeWvs3QfydLc4S4JSaAfHPOCeF1WjlrhFtYf29lQl0ZED3F2MBZD
GvBld7svMyR/KnuiTRY4SjoAg1HOkjmoonE+bNYZWzJYPkLctTACDXE56YVLWCdK
uVx2orIn/PcB3GjgXFvMAiwK0cMDo/YaUWurjssq8vPm03JzZpJ5qEQpDR1Zi0cg
/fL7rBpTdwl4Cxckiy3gZMcdrngCsjgPc0zZ2C6GRfVhZDoyRFTNgl1IgtYPJwjW
c9j/ZZZHxXyefhIpZXnFfWjkrRehgOnH3Rr4K8Q+tjt7Q+2rrz02lkiybpf02jO8
YOhvmxCGMciLeaIaamkJErD0HwN/Olw8W48aoG7YfJEJJDnh02bwQMmiO6V4NU2r
30pPSge3ujpMGP9xSsCf/0AFRTxvfM4SaqLZErLR50v2AJgDNidP7f7UVmspvhq6
xhQ2qoFSl5iEWruqd+VQZOyMptRWNrMvA5YrX32bSYUSMLRp98nvu5ccx9Yqu1rH
cOWKZvSB8GNp1jTV/Qf7MdOTCejdAFIh0Nei7AWXed389YZWepLQfVs5s4Mu+UsA
f0fxaDsGFX01QvBqCKpCCLG1Z4aTYhuhITgil8KLNRNs2posaW68dUOgSJu0BiCb
O04STz7JnyMNj1gOKbUTSBQji5jwrcjCV6Hx1HgqjE7GVu0vmr/yjmlDyjL49Vl4
uieNVrm/BnDoT8V6wKNVobMbnr7KaHVcRN5i88KuRVPCmAc/4EmLzadHhDOiTfF1
pBeZhGgSfkE3viO02NBoDuTKm64/YTl2KmWaXV03GQDVPzjj3EYirlUqipzhJsfY
JLBrU3C171O6x7YDUfyqEaaF1ptymbjJQzhmvgYuBnOWG8WX0cpY6L19pan0uE/A
/QZOVapDZtcDrAWG5dYtiW9q7hlnlba1L1wpIllvUqGl4n4HnAufVy3lGys8bSll
LJmrmJuyREt30Whq4dR1C4XwrFF4Rn98w0z69ruUdIK601FwPUFdd4G66r0BVOE/
1bIxMFR8LReoL5t8kbVpy/+wkprxexbHT3VEyHRz47ZiCwri+JJk+YRSgQxKI68h
+H+FCli05R1CrzY0vvBKkVl5Vi9j+JO/p9G1mfqL203WoTB9j0j+5aQSj6JZPCpR
KSSjY+Il2Cw/jdfp5BLEaCdLUAkPs4eIvDkU0ieFulo2ilvsFHh8uJJR4GvC1N6y
lbDNif4k1jTcd1Pz0XzSJcXMusySGVAGTcvQAVY3Nr2cOFlYMiY/kALWsks/+HaJ
qu4XZRWK+Wq+ormGqI2+xrvjvmakYOK2/lYAGimjZbm9LYKWCDfvIpmzEcg/Yjdv
2pIxC+VV8HaYsCPb+SYVbAlME6YyZVq0wRcQ+uN0ADiyQa1CXieYVBUBx7gcrM1Z
LHH7WX4eLOnY7N0YBRGgP1lvKUWFCyyKLd7bg4hiJC/+c3PP11OMu3IPewUCXsKZ
osSVZC0JKOj/lxu0r5wMThvkgZA3eSyOXTSXPIfup3RZLLgAqA7O4PTw1C9h94KH
/dttnbIossZl9f1ZnLKbu6wv910yfpeP49hwA4UurIQX5dpW9Npzt4MxfI8JvoT2
0MLrYqlaQ0BmZO5lezoJb5a8okpn67UqWijRXwIMjC9IvW2SxLJC/H1CEopH5nTt
GSD3lic5xCppd3M7BTM1kH6/mB9t8bW1j59MNhlYugTUHdJ+dcQebgpmx4Sr+1xV
R81P3R4GPNzIDsdrv9fRP76cDwXfYJw3UMktAT1QzOnPYT2rihCAjwmlf/jH2bGr
M6+35JZ7lGNupX1o3HjpS95X9Lov7ZrZPuUO7FpLrtXcVR0GOQ/bCzOQKh+tYDXu
qb4lMJgI64k3ykEd9L9J48XpMjTQKW7ZuulF13ST4zUFlv1UtYSQuksaPvXgNKeQ
ToqmMpgSppKMrmd+pHPl0jzw41zxTceMznMGJ9H//JQeCg65vNbFAU6XsKNjp5hP
i5ETQhqTFOv6ZDiQ8xx0ne1d4AGmZeFoVsWXY3q0HZTYYWdOQnwOAYge2tydAUO0
V2Oh4tQRxkU+bD8GpN5VVMTt+jGg3fHQUg4eIXoNHp4lnV10Qy2DH137CHVODsz4
GqPg0B7zUUFVWp+WBPdavNs9zVT052Z3sYaJ5SwHjIg1283QqzDX4fSHzn0wkHZo
JhlS8PimSYjZDWFPltvGC2AMCWGbiRPX0XS547kFIjE1xXLeY3zPodab8mo3RJ2g
c5z/O7TqF12WVCDmDYBgLWG4nzfytSLnK/kr1dt8cf4/RbgSZUXLrfmX7ON0FE3E
lZa2ZtYrTNVilGBV042WSqYqqK+pu6JLAu9IC3H0OKZlmu8JPKboxmPL8bBBgOY/
fI5Hc1AY5KFmJ5plkduIsS0USTIePrXCdn07EoBswkDlqFzArX7geg2Y45Ct4onE
5Px6hTuBLW+gZZUPo2TsqNpTxPYzcoNE3krgSnKO72Nmixr8vhbHhbswSANrGc7+
p7gSYWdx8O1FQ2r//IhTMrVEfEgkNoWEOVf+lNKzFgs4FELgG4nGI6PisVVOfYjs
pbIkFDpNdOj6KUefAobAsPMhtGXlkE9SU5NL+4MJZrbiP7jy5XWRmblQV5CbkNSy
A3+TSZZ3JF1ODboYSFJnDEmQJ83JiCB2ivKTTfP3/2zSsCyuTKz3CpEzTdcVTf+l
hEVf5KYDolV4Aw5eQ+KREqcVXYUvcI8gvpyWN1iyhUA6mZl1aaTMrym1yI0L7EyO
NavNePoLB4tnztUhek46MArSCI0f08ooiKtFNNiO5WHO5aTDTRN8MhW2n9yCgJhD
3ifKP17vUl+EVgMpXQisNarQhAV0+toDsaZXHNb62pcscJwsKiw6+olfIglmAOJb
0KjvA7JEdcm53aIgymMs2YHpCO25mFA42ajHx+9eRc0AAq/VZKXKgD1TAXAjJsVE
p5a9Qtg3Onr9H139B0V8k9sDZKiLM5w5sEueNMlIVK3q78VdF4PTAwlzqjeBs+Dh
IwPw7na+t3c5EcBsFTEoxhX3AUkNZy0ffnJRXqOnwmiy723mcNX44iF5P9q6PGNM
X0XJkjPj5chGOAW4ENabsolMmBaI2MXo5SqhY1+ZyRFlsQRtzkQ9G2I584BL9IDW
ULb2tZnXIB/i3YRGgpFnfhYRoFT2MBOK7EAuWBQvv5/e+s4PiZhL75cwjIzPPMz8
wQkBgFJ6Vj/tzHA2uFxFlyEhLkVrn6XvC78y65hzkVdo9LQjom7EEfu1a5p14X3s
/O3ymWaGcsgcsXqKqqwtrjX8rOOPqOhgxhZHasXDfqLA1AWQZjv0EanIDXVj+nNh
9eQGOgXRE8isk0MCSn6i/W3NYIE+ba1OIjBo3DF7aY+UlSEprD6RE14okDZohmjo
APD8JqYiNCUlKyGuKVwzpa/m1nT6JR04SUMTpp6GPPcYA02Asn6prqO9KKgvlPqe
df86XA0P5zWLp3ACUWOa/NzlkxuB8yl82J6rYkj7ObURvZSNYHHiFbyObZjaVTHv
NqiOOi5NLx6ZhmqjG4C0vZ/matAK1hFne3PCQrK2sUJ7g61M151kEkTvLM3dYL+h
B8bRBEFuX/dGxotHhp8JynEYZ7KZCRu8kb1YT+MYkLeeySIQcJ2uSaGsp2x2qeb0
+RQgk8QDfmKGyM5ZEfyT8oJLH7by0SJvZtXCvGx9EAyrcF7DzghQHtjSdeooWyEs
xA4NzJzujFq8Jk91JZm/ZPOwEA9GjjTn5A1lJPaX6lOre9VWmlg+oDdS+LVJl4Nl
86HJ425obNTaZ1KMFcKofsamwexLxuiW1GhbuKMpd6FLxJzYu5t1IVfmBOVmNdER
IZ3P/YEqt4djDoFeIKegs1eKCMCxwgKSmr/EMeWfuaOjVqQV9kV8tljTlaLjtmyZ
q5mCVQe0UObBC+wzmo2Am/EGjpR2AMyrWJO5J4e4SCYr7LK9gsJNTa7xR8pt11SD
c03JOvn1aIlhxTu7U0InkQqd1PsoV8xlTw1dVK7zA6bwB4J8jzHn2qT2NOs7WV3K
9rIev8g6NjvLvMw8Akv311+ZN/OkQJEkFmSa5N7pNdTJ7AXRbXx6jvmRktLuYzIX
PtyXes54RVFR49aL2RIcfqH2Vghs8P3gA0xeCatWSxorJTmZB4ZpVv5SwintpcNV
xutVcYkHxzThCuQJHxpTi0ZJXHzmh3w3g4+jTX42kIwyztjLnZbxWPPg3jjC5TKm
c1eOiLKrmYNOib4WpSR08J/xilpcncj4FacDOf14pn+GiU9xIhlTDsR0U3of6LCd
kbhQ3Mx1YL6ELUfVjYvOCREk3YrSyLh2KC9qadaYH5r9lMd0TGk+teFqNRGmVfZ0
tJyxzevLEo12z3Lj71RZDhb5XLXz3Hi+KCQv95pRIkONXQvZBSYEkuifyWrJFDuB
7XOmEDPbef0ed+hyvQu/mvwzioNUiVk9V74oOgO9d15RTHmUWcdoQ7m+o7iVDuOU
j3i92kIfdZ9SjxFmw1f4Yv2OkHSuUwumqrk1oIL06ykPtHqLug8TqQfVgTfpCito
8gLSBI28NrLmqE0i3t2beIbiDPLgORBNqHCqdAfP5AQbMqYZLFKIfXrb272BkXOJ
y7T3fqxqlDVVKpzQvYcLQJgvhKRU6qyWkcZbwS8P8liDgUeVzjE8lhkAnZ3op1LJ
Ru7UmPZ8GHqfc7S/vJMjSamLLD/6env/yLPSjgjJs7deE/zqT/yGGZ5xpwXCEPP+
fUK7zOgYGvDdyUqXiPqe0Jn6e1TVrmZRaJFtjuoM/gBkQs0FhgtfaUpnBS5rjyMA
B5MhxPILspNi1I4lZrhrcLCIorrnQ1YF14Gd0c/YEF0RT1LQ1Z0/KcLiFJll7174
mlDGJqIsfthGUP+V7Ua9lKm88lGdF96rqIA7mLNsZc+EGVow9V+ah1o7aJQ6mYfC
SYmrDa3QgwGVmthkrIYhW5Q93N2TIKKxDTWsZQOCjFzi/vbLcXdgEABBZiaTFtO0
ULhaPCjRhlq6cpccFAYWJ2ivwDcJpIy14hOv4IVBhjfV7lQ1blwH2oKiJJ3NvG+D
i+sV+AvuiAE7cUlzlelr9hT8W4ehwfgTYJR3ubKAFfAnOaGPQd0ehxNW6Umuk5/p
PmGA5pOIhMSp8SAgJqpwN1QtQQm90AyiXdROvtAqslR3Gkm3BaQG18+LtA0vj95r
L7rT7koXYI9lQadyNF+DxOf1UlNnvOIrN/4JwszC3ZpXMKGUWa/KS2RAFpL28A3S
l7xcpZ+mb95anQ1a8ivWaJdNkBjucymzwGym/g7NS7EbxNCULMlok1niSAzxmq5p
0tJUPrCzfwVTcm3bjfzDJiXRRHB2lUB2h+oHkRdK+Z9YEJ165Tfae/nOVX3VVbJe
UytfaBqM13ibzuiOnRR9KJFDObXaXDCEUCQMKvhHAmRu9AWP6TOSBFSZJwCY6YmC
NOlaNViyMZ0+yL7HUvg0nCNYh/o+jJSaSSgO4rxU/PU2uVDUQWRh1E1BgTy2QsEc
Qiw9tp4Oo5i+OGEBoFrPZQ6ZmLnKfpBwnrz4aJ++2lg0n53ddqzFE5yBRZQ95+9N
Sya0NKphZjiCPJEbI6rrtdt0BD1RImxWRhwggdYV9p3lKk0sEfAs75zeWlAbnbAE
9ggvTOvCsQNh9QPU5qw8KxGjKHXfeYctH9ZVMVCVU/12pUKFVcICU3So7hjm60ZR
Tve+QB9qv6Zv9z6rWw6E6YTtk23nEe+jrz5s9fvqmnr54oIbOJBfoNsiM1UHgP5D
qgCPtlcYklqj7qZT5eiVtuNe9Ic+UKXfHejrgEXp0kOX2nmDO7ueFosxqAX2BdzQ
2Lpx17VVdsZfE8w5dFe0HaCfjZp2Cbjb7rU2POB2Fo4H1e0KNW6q0XmeEDypcjoI
QcNKqwE8ma37pPBwjMqiWAVcVqWJZ8cmiWUt8DOOFGfnxepIqdpGS4zacOcQx7t7
wdWeqv85iUvZnAZSnw+0wV0q29SqyrPDqoQRApEnH/KJIZpbg2qNy+9TQuLitQuX
J/VphUp1eZsTK/+QrKCRlQCXa8FiqSyu7NLt28h6EfI603bJgf7sOG1ItfzRYICG
P+cUbvdDuW599+YsZwkXLa64KrM9z74kOn1APbLcMexarRAcr4Ft/1cRh8TDyZ/v
U10ywoQqpa4roWF4lZVA4dkD0cebvrZMn1o/cFs7TVdTKEWJDJQ3Lrsom1Q2Was6
BLzrv6nEdtwRUIB+SUW0yccTV2e3DeVu6+FXLPBoX9xriL6cNdAcQMusA4B0IeyH
Wt8sBFCGZUfeIoqRF9DcCuFHfZ8aDkfqlig54hvZokOpI173jvRvHzmhfXOkCGCl
RkdaZ8Q8b9eUeSbhW2mx9tbDU5dy2VZDx6ARwIGcibDKjArXXByYNtWP1PObcWeW
P1cJh8rbY4r4xO+ConpauIerPvo/ehuerFwrHTN9aTCCrz6lg02bw6roi5OymW5W
EwlEdatI1Bhs1w/BPChTFH6sOs1xljoyYRMr91Zj77CoVL/JhB1BVj5HBnoYmKkv
IWuvMQxSsicJdw6hiRzIs2Kqckux25X1LbBCeKUMFBLfulutYfCLIVKFNjQwPHrR
QusrzE1DMSrlc9fXEIYGJEVoZRlN8guARyDX83rGUS6ij6Mid1WHwWhjvPrxV5l/
8usWlzbxL/H6GqgxKBQWjr57XbiQJIkSDK9FyyskKF8cjl0W5DjVLpu/xS6xHZNK
ydy/Ri0WbqMv3cXxtVfVUEG8OnG4ws9lGceT6Px7DuxK+vZyXzNEjn/imYGPWI0z
BNoa/9GdE3i6w0uLyNi1QAou/A0dRzqvVpW8aHjyYqiiPu5jRuB5yEeEbYOcCDFj
u3kbEGU0ILBkG7fv2/zE5kpkE9CyEPPQSSCYDk6YfgL4YLal+1i6qwLgC+VZO1GL
yMz1SyGmOlEMYMxSKZCey/3XgEFA+JNW37jD9zROTE7La5rpr47bjG8AcvXQRS6D
BeoJ3IhRKWshp97tR6XG/36WZZeCM8X8lo5WXg9nZ9NH083ONKkqIymwebD8G0+a
dDOVOKA/tqUSo7Ld0ufCprKAktJXibqOgYzy9rB2G9TgtxbLe9LL6uaCUSA2PYVP
z3t/bYJQeA4NxGBRkjdVEi1XtvSFGeJbd09zzFrJEtIS1n9zcwojegRwIsT2git5
tR9LndyIeyHAeronfhU0MkkMbJIfHS1/nWw7TvzA9CVYhmtoCYtgYaXr4slmq8zP
qDu/3A/spEyt8ynKOby+Cr1Dr6nS22yqDTp353FCWe1yJbAZruWnYSxm39QAIF8t
vNBLQ8y9UaQhSbQCWWqO508n3UW85Cg0JFSqNojf9CQmMSOh7lvPPSrBjo/u2N64
gRCxAjkL+SStNiQUUZolBqpfmqMkbvVBP3liUyR9ofMl86+IjwGOKrDUkyJLsyFh
WCeGEJRilmLb1R45tROsbyzzQWpVdo/rDFSRwU2ga4mfrnIYmZ8wnT+ttMnf5O2A
us9HMNJRoafiJrkIFFlHqABTGmpf4EQWC607IPilTrg1G17wIhy6C5IFZe7UiWnf
PPjrYUcCo15nlzCE7JI/C5WZJvHpbkgLMCPviUPUwmmT/B0ujAA73m87xxbCB2T+
pkfINHwWmS0ZGxom9xPB45eZXovddBuASBMgJIbHlaDkxuQrKBMsaHeca5MW/W/C
xlwQ8FLfL+Vl7wh5YyXg3hnLnAtVtKwlF/cwn/mSRxTOPshhyVNpIjfmbeXgioJt
0OMj9D4nMb7cXZJm1gNajwRaU1q6cGXsnfXISgpxxK3vlAKesgBC5PgVOsPMUhmF
ZAJQKYp0aTFUn0p7SA7Epcp9oSCJjk+AngB6uo6y1vB12a5H5qlJ8O8BMaEQ4wvT
CNXAqLCXh0rAsqbaemi1cAQHtXc9yqoV6YEB2OF3aNjOmS1gUYjcrw0v+MthCmep
Hke3YxAZpMwSXc/z+Q6mZnHM82tj56scEmZI+dboGrhibSxVcyo3yackBnqj81Lw
/bWjTiqpxbBj2+7Mol98TOGQYwHhIjx5LHWs72unkzGWxHiZy3uljmG1PuUut4Fi
K0CW6BEiQ8Bn67sdbEyJ09e1YVoXftM0LOWJdhcjYHgxxDtGHAd1f63S2V0GHnc9
F5c5eUIgs6Mi2Sndi+jKIJ8mA5dEb8qrfCVRz5xWgI3KsIbPKKn9/qu5D7yiIp3/
kf51q3OaEh48QiSqNbFfYzjoYSOkKCfuB+jLDxRlxqtppVRUnTzn8iDTlCAMfcWV
JiCTi1CaiQ49af2K6qzgK/wBYD/AsrlVoz6b98QKgogqtfyuleNz5WjFx/AX3a77
s4GkqgVOKGB5PH3seBfH1WPSwIpdICTPZdlQgdmjdJF+Gbw7Zqudo/DE8bdE1HKB
HwQLGA0EOum34/zq4B8g5mKYDaGAWiEkqpkolpg2iEj/PpIWlKx9gPZXxoUD/8vy
DJ6wHji9XI+Qq+11DAshLa4R3wmG4qUtOKl1hio9madVSF2mrgmWf61T4nEv2LA5
OptnimjxlBran3mIvnd/awPhKYRgNQ2LHmYOQEUzL4J+I2aV2j2pML14mlLFnaIf
Mljsr6Z3pp4s1QyWfciIYncl2fOs9oglOqIHjsZgbb+JFYC2bc1H6zXYGmBj4qs0
HKnUUOyU0828k3Hll9cgO8MduHQzecBgtV2rfsEgTMUTN6BDUv848P30IMj8erD+
tALWuskNNf6lU6iInsS4R16Xmphdhj0m85Pt0HJkkvDdjya+DojVW0FofF5iWAWR
a1DYiSe0UpXCxMdjsc1ss/jUv+6oVGXfHqmjuXZ5BE8+x6I2LJRRDzqaNUGO9UTf
vBjQbCulgc1rr29L4+1UjpfQKiPPXVpnaQGjYG5EZzPCFk9wpK4d7Lly4CP+T2or
ZwoMBE2ax21fctYV1vx3R1MTkJIPULWdCEiD+3XNZq7paofHd9TpkRCSBTRoGoYp
eUq9N6Td3rWBjtyunqIhyvnQqrc9/YN1te++ru3RuzENBTYyMOVTLpW2xOFFujM7
Rg7xbT99cRZ+5OiPPWI9aANoBtICtkGje/gDiC3i1c52ARdPScwd2N5T8gntfcSi
tLMrTtRs/lkAYt3F3uox31QA6K6K1S0tbm9+OzGy4jDe6Yrt2fNumopOLXdi3ZJ+
+FznNjGhmTtCc6ilYONpGqmeEFtuvT0YdN8zzZReUkJltZNtpzs5gZ5gC24m4dJK
ECuSj5Yt1vZkKB2dfotf62xfPCz1+DE2o4oIe9t8dBtqM4wCMjoIA9fjXfih5VEJ
HytWG2ItQ/QFxUQXDJr3Qy3T+eGtIIfFluojeOhvxqEKkM/D1NElcHLFc+KcXD6l
cEd9jzO84YfdjroTE0UlqgANJdPc6/7h4n1NNvjhcsNdY69RSCCJxqs+VACb7vUM
0V9hH9TIk73kpy1aBdcGISh9tdn1mMQLP/sgJDyVbUcwYLOR+NR730l/nSUGqnq8
nn+gUleBa2sCDB8GUP3gXHcT50JAXPhzqTxl7//vwHy7K9qABCdedYK0zgPhGFAH
IMrD/s6uc/50nsdw1fSQCddfYK//Uj4DyhBWYj8JXDr6UCIxFY/YtBVlgvLf7qJr
eu5VvieqRx0qVmus0o88hjSWiMlli/r/Vparvt5r4uUhFKJhu9ghHed41TCpnf3P
UJUbevT8/MyZgX+jsrADwXsloHBrh49WSIllUAPlHSGGCG5vEX7sRVB2vT48EwMz
EQGk2j8IATfS0+md5dSOJWLwt30F/4eha0vXpAPpkCWYM25M0nNuREWL0GnfsR8D
wj7ZLGgwmwKKINSmsDxZd3jvEp0LS3VeQSM63XqYM77AzTIYnlBXda6dmW6MMZfF
fl68d32RIOtkDoEtNxxRxhjUb2agwth1rMvsK/3Weww94x+ul/arCw6JgfdPwcYy
u8rOPg0EJQBGsNWWezia8prZQCmyevWRTrYh3t6rWYZofuiueSz8wKUHfeKxxcXT
spMJHaYaCCmPjwNsXDMHRr7CajwLmoo4m62ZxszfqPfzMDXYnt9xUPJt7ENhFWPA
rpKVgsrTym5kFSuduF2ywO2/QusLTE+gv0qCMBzBm1kYtmrzhJPEAobbGyg7eEm5
C0R10pFXX2VshIlLvq2KtSmezx2IYJR6vY5NMrKzVRNFP12myeRKKk0s/er3ac9a
cLcKNMzIhY6Zc+03NR7eqaN4bHU66T/e7MLdYTVxVXiCUnXbrlYA/RMHAFEu9TkA
u/y8UUwxJx8i7ERA3B03FIsUbEKClW6lAHqARQ+vr2yFPQ4bZpJ0v3WkhZPZx1Dv
sNrEaRVD1qtc/4PNcjv3Mwx1EqfhshIaRIQlbTM6pSnIO4IUXHeliouhjthZDr8M
2HluqhOFBi3tUNDeA7sI9RCUZBxFLa9CKyLoOEK4kJJaVVJE+l24ZanG5bs9lmXR
haPJkYgcDn2sOyzYp1y3cYOaW7FQmxAtvKj9ysPVr0O6o/VKc8YJsup0EFEpiUmO
o4Momr8qbZ/HMwwXZc+v6Xv0jya9XbWq8rkW4/p1go7+MDf81UC3WfD4wHyBgXdo
AuJBK2/1cMFuot93+2wp1Zdcbi5vGs2DH8Kxb1XHZ715532psIITen5IJupvoP+T
M8AQl1VTCn27jFTp3424wAXLRwka5/LYC09Kh0PhTfI97OJC8S+MsaCTXngNfhbF
SFjcBmKajTBBRYPfIv7MVPx5msUpk5h6Mmwhva/M/c/78FuM9Q0TtRc4baH4d/q/
sZ/FoUgUOnml32vLqoZfp8LsDwFCdHLNZ+FglYGXIB267lh4jUiaRUv6tyf+GEIF
iD2OvAfG8zhJa+LNM7uIc/IcN0mzy3Ahtvp6RILgO9h4xM0DmG9pmRx/h8BxY50g
jz599SKC9TiCBErQmAHTWNL53HRdz455ahGF/hLlTzID+1g3B7Jlw9AV8tALnaxY
LjbR++v3k+IEKPZpbOumgto0+c7LTQ0dfVN6+C+5PyEZLaypzSr9xT9tWQi+GFXh
a+BLS7ySCe9r/S6F6AgaNr+TBUegJsOLyMziQhG4cuK9nIJy3rYwrJ8JscuzF6u9
cVcnUBXk6ohPcxp/7yTL/ZxnqWG/3T2pSHTlUL8Y9XUf98fYpMDK0getn8i43k+q
qyFn4G0lDToo6mxpnH29qzqufnBXQ6rMOiAGa19G7vaHGYwO9nrXCZJBLq2b7W58
GKF1rw9wk9PXmIp2mnVk8cPlFpEDZp26nywXFpI6TbVcAoSC70YxvD7IwCrkMfLo
fnMa1qodHo4AwcLd+6A8zvRTWUgp2boNkgd79S1gLr5UDmErHvvS0ILEASlyq1cm
WBWf9+VSqf6MCmd161tpPn0H+Ybllai8ev48h2PWGNNc1SOaYYlnh+vH468/2M08
c6JUu8axhxy8om73suRKMUwQTPWVaKiSmH6eugZPxS1gE95/tL75EyVEXqH7DNHH
0RoGvwuYF89Bl7mi+AVsbEWPrZJTlGf9/fNYKm4hVPk40kpOJJIKqHeghcY4Ti+a
d7Ky1ZphFAcz6BuTYV/NPv83A+DmhDxmOQSB2tKpLv8iLj+ni5RV02u5FH/1Qjau
KUoFETVTgueQm3Z9ECXHzw7t7iEeMxvQsqiaU4wWzJNlC8ftqkq3hulLAYBy3KnW
aeBRVLcuwkbpp5gUBLc6i1ZSiUhFMNnd1E7j0WlnUWKQtX+7CY0ElCcMoR9LwsP0
/PNF345+yz9ef38TtMgDd5/aolj9xCYj0yudBig/cP1zRIFWq3s73H79icFmDHQP
0pSTQHQryWCmZYKjt5IahsVH9Xbqugu85OZ9UY10wlXylRePXPfvX340X2QzKgR/
VUJDQJ4CRITpW/Fj/4/CHVIxheos5G8aHUgVsmlUwNmc7q7SSMTy5BeYfr4Si/uP
SUZ+j6G1xzu6F1cLdtn5XdhRm4KJk/pH7pILv0jedhzGPOOvrsiHS8JWJB7qsntc
UZGz1/NN0bQbRcP98dLaH/3Rj0fx38Djzb6DMWqpqAq+GtpVNTKfZW8PjoJnWlkf
abTJl16JWxkRu4Td9pwgrXIV5yJ5NaN3SIgjUi+KAityyaO2QS7VakIYGenkmYo4
oOPvPW+3uVRNfvtgRvVc4vgE7h63Jo3GH605xZh8E6OYVN6i+9fyK2OpWXBZd5Fb
LkO3O9RbMqStkqeFhGHbcBCDfaRPz6Dmf1Fpr955Ize2iHrqtXrvjEAR8YyLFBJ8
uHkwYM7lKOdFQzk7/3BYNXfbOl1WRghYzCiiwErKLJCBIl+RAPjqljnWBGpFn0fe
vgrYuw6H2gRWsTzG+DAvMrRGh/Y6km5BxVexza/Cnv1C6GFKUKmEPKxv2kfp2ADZ
7ZJ/eKOYRGDUpd1S8Om2urAS4dX500KMT2aWdjomJVJ7Lje8kyJkWI2gNfvD49yk
TMEMf8DRIgnk2gjMVPHaBEo3Pj0keZA8rxPeth4UC0bX71f4YhNo7er4COyR6ITV
1pNRqD68vIj0jhUx7YjrdKryscPOWZfUqE7HJAVuio8+skOgX45dlq9Z992agJnF
VM3YL431/0NDq7+d4wDUzZntNTkxSJFFF8hc4DeFqzYXktxbjr4wwHE0SMlQrTHe
ZZwN3etySqvc2KP+gFccwpP32a4OJNC3ekKswALd08Upti79+f4MkpBp4v3zMmEA
BakoiiXkZG3QviVhAo8v8o8RZL3qRyPZSuaT1YUR3FHRCXPo8D8KbDMqXl1nyFMY
l2uCU78WFWF0Ljj4U6ZVdBspXIcYl0E+J92jZW34Xs56QpIt87Zm1psQ+esdDWYU
cFnXgpb00pZ4zfL7APHMORhdXzIvW8z+R6G11KnB7u+3t1uzsFfYPPS0Ft0S80Rt
Y4pdP5i2L3phGiZxRGqNjHntbu256D73DULAqi510yKOODWTVgSptNjcl1gVy9bL
WoFnHuRgrnCL2DremrTElOV/KLhG8gK6aGMDjqZd/66/YQuxaxEQlI3mf6t+2F3B
ohlzl70tpoD78rpo2DDHLXBFo6gg/R56sC+AisfNoe/FGe6LxF2ev+9ncjOUAlca
id9AsW0JWrQ9Df3JeQbct2pTF8AIV1/cNIaFwNhoNNTBaArTYjtnZO1NDTOToRK9
cP7gjUIT1d9rDPZZo3Q9JW3E2uUbW2TZosc4i6IIUDvpA1tWql6ezfEvA4jNVbyh
Q4huvKx8WESu2LC37aBDadW5400U1kacNar9FuBGefMSi7TWnZvW7HHXsH8EYIA5
In9k3Uw2QfILD66QniejwI9jerjIfTXPFn9D5ZlalyBBHHoHyKOKOlkZRo+xxIRt
Ckh7l3hR96HkaSLjutwwQEAdtGuHve/+AbbOZL2z2t6EuYv5NabgL/9p2f/G3QBS
qp54839CkTxygp8N7ioWOKFTmI2tewMBjnlXCUQUKRmmHzYNYz4EqUBx/4q9OVKe
do48jqumiqQhpy104YXiRZeITD4PvlPH7glO+s6E/WYVOcMZMK8UqILxHlhVln7R
Jd1ovNKjg2RnngqxylBFJP62G+5kN1MqRtxs8TGVvLvVkmCjVSamFMU8ai/pFcqo
dq5vgd7/8wN3Q7mD13azy/2k3Usw/r2YuFnfU4nV3NsRZYPpjCkLElRTKLhIYUyB
oTNiEoe/8SZLxwqNfQ9W5+9N/UcUqy4Ow8GL05prqGQS6fOIfywdp9dZjMe+yj1i
ulDCmma7vhhFQxqeWe+ILdHm9qMM/ZdaOqKBtStsFYTMwpyWW+4+pIOUceHoF1Bd
QYm5nucaoJRwHI+RYrgCVrQCXbaOWdxkqZG4Qp03MABDsmkXU0G6vArBmdyzqxrc
IETm3AWM8108RpupSltTbV38MGH30kCHJ8smos4CVqWsRQ5z8zQhURhRnZIx3Pm3
VMj8yYwap0oR4bcnbUcj7FdwGmwZy+tR9B/x/s71RRK54TgxeKEMlZSto0USKxsl
/LgI+sjaMF/49uRav1U5hWB6MNn7GC3NkWELxTNyJeRRHm22PXEydx34qcMVx9D9
KMTtTg57CiTL9NA1KZW8lfcIP92BQ0WuMYVDgyM1SeC5rMKdw0fWUvBgsvoF0AzD
abqY+P6Tz2AgiaZNmWC5Hr5nSubdA0Cu25FJLNYeDg4v3hiDR8YPlK8tZ0lVyi9E
q9xKG+Hewy7CJWdytJtLgD87oxrnQOwGa9flSdfagYH8AId5FpyzCA4rybK86l72
xv7KvZLO0/V+GfnD+SP4atyV7JBYXDLA/94ZDWwU2eGy+5A4SzpkfHzEUh9rYVLA
KQcecf+j6LqYE5vqMI9CTR9UDhw8MAASHbdusFc1kAkASxjPeCBACcfum5Le2HaX
+fRYrazZ0aL1oFRuGVjWmpozDON0Tsv42HBwPOzkiOHDDFcQ805E8dT+yX9Qh3Wf
QxNaGOYPyvzbEDi99WtkDY1VF2aUCM3po13cj4CHZ99XwqDHNiHgmXZ2IUrWkcCB
8pCexEhW6ujWHpuLqnXdSe+tJY79Ba4kiGUfsnHyhiK53N+PtssVWuznrhfvtDWi
vrV80YHinVPgZllDacksfO3QzgaQuarD5a0pBzHegKuMIy5ZJyRUaWJIDMDF9FXy
Rx0a3DIby40CKZVzPJNDE+rTHNKOI7OJGnkUjXIiNL2aCrO7Xjv4CghV4w4JaZGF
BYetSy74lDAxP2acREQHx+DHZ2YXtIJp9r4/EeojfM7V66YrGhT3jrbp4aR9Jgon
+ZuIYdfmBvBBk8VRvhW57X7E7oNaG0vJlDKke+8ySo2fyLIOA2+4JdRrLtc0kJkV
hkjQe22Cab0Gl9hkz5W8pBxuUJgOkoqCWkCSlsQb5xLDpNxcmc1mM3BoJuYlJnLg
wf0JUuAhRvEWxgasTaX+occAnN5pUxdTbRqzKIF/f27whKoEcnVmOYKW6k66GP5M
1Du8CEPvgBJdVj1xJS2BWnZ+Z1Gs97KeWeQQA8GlxXSCcqWf/NqrY+fyBxaCJgk6
OqZGSUev1ze+sbDaSnJLW8rUJ011ZUpzDpVzBWqBCfJgMSq6DFMbtiwOvjfTKv8g
nVwTjnX4dBWCM//kDNl0sxgM47ml5Kq69i4P7tCGkT5XgasFFSFiURN+lhwGCdCN
YddSQKa9JByJDXq9KXFgDVjbzv0y8T8/YyW7t7sMXt2lcUanXFqeQ04Am3RU86pa
vRjZlObJzXqywiWtNl8T4O95D9Y3wLLI1nwHVJ2RKUduC1MuSqmkKEhNh7hkWg/f
MDu+7Rw/7g95f+cxc8odihtfwK/PExyZqSppQyTteKuyPBH4UWM1JfIDmCocUtg0
U7b/yFwoTVBYn8TPIecaXECT80WZpgceX/wAMBuEU4+qVxaFrmVrsYLTW/2i+97z
d3+2nrTf/QdG26bL6LoMeJVo/2pBNcGBWYpjmB2UitM7lh611o9Za4ipzk+o8fwb
TEAEyY4HHaJSQQLdU1vB9QrNzIevppPxFHnoByVY3vfFdJ6Hp6IoVgwO9Ax3Wsuw
eEGi15kzVq9M+6gBozZyZAFbKHirfmL10QOv6yu42bacnpL6oF3ndhsBtPSa2QN7
pr0n/q6OP8fRHqTWLxzrjBNvfC8WUiI5/malJ/QzptpEeffVjFroJj2evvtPwAFm
10TN6lUTcBHQOmdGwDbDeS9zBUdzKlU2i25CEoMpWSvAx11bb5zAAYUViQ5uF5VU
3shB7G/RJhkTUZvlsg71EEeJkGdB5riTwvFWBU05EVy+20sCbhL+QTMPhkinSeOr
vSJOoyagoHAeJRAPH5+u8+FKSk8c2suLmTQ+r8FXeC6Kmb0bsU3MFuPUfZCFty4P
NDQ7ewS5aOARRhTTc4YHQ7zxBLPYzAVR2kIGtA3u6Cag0DNLNTDBge1ixk4O3+2y
MFMkCfzsBUT94XJVyTp3DDtS58geof6AooyinEvfq+qAA8JvMMs8QD+xtndKQejN
h7072vhVSh9ldDRbi1ogt6tx/it9It2szO3a0dKBR+aeQ7UKSC5z1ZoDIB4ZUC36
3xQK2bSU/jumrQxYVO5sN4nsp0GtSscc4yxEX3D3f4TkF+BgzkBBqDy+i6ZukM59
XTTHpGDJJ603P2AEcWbikAaCO6UFRSs83E+t/gGdhTuESd5HKqZBNx2tXps55+Nd
ihnqT2rpexpswakVfm9t/IwEMf9/LmfRvbBnPcqoDUdC/En3XzvmsmOSi1owNzEb
cvg7ewtbRZ+02e8bU8OKBIOxY54w+Hr5jyGSTnLj2ldW7XVSJEgYoWJzja+W4FYh
ZlUvN0Y1MmX8iwwtuSsORJR41Ogd6TmM7shr6wrvH2xxorgJ308r43B1Awc0agil
2+f1/dh9tv9psBpgv9wfqN7Lr7hrQggu36YPHi6LVNn5t0OcgDt2L0Zs+cNxnsMt
Pw5KWcXre/egf279tl3tiBVppWDj+MDTVS4iUjiJFufvFWSlQTr/mFprnZJjItXY
C8J9OEIS+JuuxN1bhee0Kf/JyuFJhGGUYYDoRY1EimDhzAT0tJGPD6EcxSyJlVM0
2/pC+t+lgMp2hgha1Nh5b4XjdZiiUwjFdUFIJ+HvbHiQ+HhTzvBAQbR3GoHBg29m
YsCmXgeATDXlmfstzkYYlROvsaCQLi80XZ76JmflhOnYnvBnp22krH+bnSMyfjlE
VVs32XGOlrYF48bJyCd/REl+oSjuXg13QbKZX3H8jRmNaH45mZIcT++zUc5frxoM
MRQVhW8J/Cy6s2XXiXyVr9ucdHkuk+OTaNY1SgBrmR/YrNOjo2lIJoTNDoGcSXud
u23Lgf+HXh/8GIML0vfnPu0HFxXNsGU9NOIf/Q2OqM52hVgra6HUGI3MdGiZT1bU
cbe8cMAdg9af85kK5hLbQbzvp5Z70S8h+oPkkdVBd9OVTM1+8aNqgz+dsi6QQJPU
pNBiYSoCWJjIgwUEYW8HXCDMbbOc6toWKPcWQ7luXUn1FRuzolq0xazl6Q4p62HT
BSLybavpCJ4s77Ow8uSq7+VIBQSzIq+3C72Ukgp9Az7gnuRxGguJHGJx7PCSleys
MwJAMCMCiCOUByzxpxG1IeDVFXPKruOSk9WmgypEhm+xOB/Bfg6Nsb/F3iXmnXgt
RGjTrTqxeJzBQknTXQml1OEvcX7CPzGY29q4UC15Pcgq9jeTVADChpU+Y522M3n0
S2tqwwtTCa1Bz0AHOtDUkrwfrY3sQyRi2tHcPD+w7Iv2+cx9PWkuZpV+a1rQAeFc
VLrKSqI/klti6xeeE6L+o1AECC7658en2rZfAStnRohaFSillFuQb2RYIjktJDOm
km4s1qx7JvT5spP4mw8bIYoKReSA7wfiCtyXU6gTP3AmJJSW8KOfsZlYCP9cBXuL
ldPwqOmapZau5o/rCiN2TdEUR0L8hSGdc8FNk+zcteN7nJkBIuFuFqAJBB5J3IFe
RjEom5EcF2HQP5fgS/47enxvHLo3ml1NyPufKtfYVKn/zFEy5bqLz3V7MFW+U8RA
4uaVXXYuj2s+xsNeig9dyeWd+4Qlu7fSZyM5BcmVv7hU+iF8YLXm8w4V9jJ2uKfC
Xpa6Hb8drk6f32tL+KH2KxOTz2W0Wbt4vLtzIFZRmifTv4K9ZtDfidaBNAeIk1Z0
OfBRLE5zVFNajdBizoCtLrdOPd4QwAsGvLaitMY0Lun/VleDx/mxmaPkhpLlP6vZ
WocEn+3n5AVIxlEmdzZBOiqRQP8g+V9j+yMzMZCw65CgA84QYgPQHF9uYAvCxvFU
ZjJoZXRhkP3nQn3YxLT9mn1AiKuesEx1FzgGFbBcoHYUF1pByiLE/cyXOgEWDnXx
6zVvOIixr1KAgHd2Ls4Tvhja6vQAVMAFNzhvAWEZDrfQC68obvTpCkyBJXUDZJ0c
pwMeBB/a+2redJ3FEiylB1+lb2qDjzkkmslftEr7+hSg0kMnN5ttG4s7P8vm11yL
zxc19ZO309F7n0chgNpSr1tQ9iqBi7ki4Kjj0jkBsNjFrrV2dLinmYpsJAHmZ+13
sFBRJI2c3GOouG8Nvcfs3A/Ehs+3nb+0CIqWTf+G9OGffm0G8kRRPYYN4L+RpsBK
Fr2JfqF192TSet2esVCEko6HXs6VMHlfOVBn21HsSxworZy9P+GdajhJYt5FM9q3
cwtRXGYJkTohV8onX4KraLoRLuFAI6TtL6rRVBP9foq3jOZ5CZ5ujutFyZoPNVwX
pFRvcjESFL05DBKuF5STNixEFwcZzQPzky2BsDgdSYa8AbiNSYd6Vlr75sQ72hMq
tPjpA2ZEAj6vxByAdDEaL9p1VR/FLn7RlDbJaqT70852twsXqv5WwUC7wN1lq3qn
wcPlr/qVrikmw6FTYKVvw5U3/hL4IqcGl/DkI1bebPI2XzBV6LGKS4/B2NXntfI4
VvMRUbDUUd/IkuuN/VOwtbBgXqy6ahN3nMpBBX+t43bMlUfKOHuDgZNz5MpGRk5w
00WUloHJa7S6hHVzgVTmc3wnL2bpX/J9MDTEisogoe7VOEnPTzW95AjVmlsxdCAL
zRallgAU0JnrPgB91o4jdgDeEX40tWW0B+/Moo8VcbnA1w07+nvcJ+mbKRlq5unn
XLqu/Vz3NRAHvuJnqWqfN8JoQy55GvxDWxHxTTuRa6Jh0L53I/Sa9+BULnEcVW6i
/haIQ237jaP6nq1W06uKa+cvMq29uXPYDR44u6tSJyZ5IGcLhS7+09Uf2VELBi3b
trnVDGoINXzpCEp0p1wdRPIw2AFoK79BlApqrGqU7SVjewSfFccxHXBnCv+DIsdz
E9j74AF1JPAjTyfgUtDLsUGAaOGPeJkhlrzC/XAP7q4rXG4e+mKcxn6uczW2O6zO
DsM63CYXZYNjHkt45SygwER+lJi6i/9qU5/39wEGVegCjaQIgNq/SbDVV2Iw9OhD
PfGOZHQO116kpJpyE1OMlAYl0KEHWN+OKLs3S15LErSOtkFFnafBDiwUgY0IKu6Q
EDKgNKghgfa6sUH4cDkWl7S+KgBQMRh7MwkNMaYEPeIHWiZEI48cNS4fOSk+oPmJ
tpoiDJzrUkMVz5ORKK62/UykkcjzRx6u3K+HnN66WNeycjL3zSoInV7zUPR9/kwZ
JqZIz/uGqWcFq5/FSx1xhXs6ancaQ8Xew9OvfapOKPpSucbwsoS/fRf7aks50VSV
6GFFaO6WPVDcjPORGX+vNu7FfW0w0xwjiCn+o17sS1h2L6fDqnzCabLgr0fcEZKA
3KFLBsd2TvyAh9lri2kSAVg9ldvJOZ7pIZ6nlLK06HdbySzSg0sxsfH5LHxavjzu
xjiwRmR+ZuvT15AqEY0YMsgmnn1yow++mESiMgd8gynFVKmYIRnTTIqNoy3m7VvV
Ec7SYOPdgx+mCiAHOUCPBIgFl1gyzNyfMsuAuQBI1T3bU/LGW55Y52mUPkI/iod3
KF00qawO34a3S5++LLMo07jn793PhD0gq5C7py2n6Kw1ZoHhpHicdEgnwOaJzPF+
Aql8/Erlnv+dgIkHYI7F70E6AtYqvMHb4RkwQGrP19RCyGz4REAWBjl1vJc7KL1J
gjmNdjOX3MtZoT3gRVjoHedB9Fm4vCInLVtQ0QBPpjlhjo2o9Ha9GB7SN7h1NC+l
f/oQFBN40oY3IBLXqkSYPj4WSzXG/zf464/1mxjJ/eSZjBVA42OhTkZXUylESzXC
xKde8+8yZjUBCmpNeqK552/a0YFsw8QafmtMsDFwKcFEwsuTaJkX0yBx+rJWj8Yu
oiEuc02bsP7KtwyuP5hsOrcy5Lc1QcBS0kFDVBLxR2sJr5NrEY5LagYY/+dRIZsa
ZJOlxEBfBziAZnQTyEZuXe6Oj41LsNDzR/DZ2vA8dAksN8EnW4WLAb/TZWifgA7d
mkGkUytU13xe5xWxhcDxRbJkUYSklCtptrWlIyER0v8QBxHGtOXnrVwi6cMBo893
+5o8Qed9mB9sahRrrA67bHtMyI/HoA0EIHPTEz8HnSHQcZWYGpAkW1hc1/seu62j
LaeIWFi5SKCPDZOMjvfEsbFZu5RwnbQFZlIDXorym2oWHVvjcNEc1BYn4VxQ0kVA
sloFyZfLxTIIIG2RyVZoZHW2aubIep8N51KivhNSQu/2zLP7D3ROM/XjtSyPVHUb
f5oEbeCR6Grnz1M/cdkXYDkmFOl1cEFIZ8JTqnkXY9SE7RVpMe7FMjd8Mf1YzKFE
kIl6IrKq2OU8scZL/WiuGfvwuqld5I9AamAQBBSt4a9lHslJHBdxfjpeszupMORw
UgYkDv54VCCloPE78h/QCBbb+4KIq6t7AqHSfNKrYppu/A8EOy61JMUnJDzn5bev
slIGDFsaQqNEK2lGw/Z3XZSAQURfZ1o9CcfPJX1QihpL2dZcCBGKQmyyU960/Aj+
Fu2XLyAhJdauAuDXoD1lH4QyKkGtAZ+qvO6lXU9BJdEU8lu2c1nSusuMy5aFb603
M0tp4zfnHbQ92/n3QWzkR1dosdK0xMosrogKHh7P2zeCe7ieeo+eaKiHeKUWgM3N
8bGGXOVCLo4llpeHN4ED6RuPyTQ7A+pvZtMqE+s/0uzQS4JLXTB4BDljED6Dfwux
r9LAxT+Xk5R6PbMTJAkzTjs01vhxYm9IIFSsSHuPh53KnqVrrOrXrFgFfskKexdv
OwqvseU7HYkds7dGfBI0xPOowlJE9YahjnXsngyhMjztkflcS2Gx/6X7sr0I0Q+Q
XZL+K0hHVf48o5sQtjuuk4k3qadIyez6zDHbGX5ai5l6nBDsB16Qw8l6ZmBNTI8y
3DSkaf5/kZDcpsn3bZiUX6FVLVF9iedTf9ueVVpiLoruAtLdTssCWAB7LeOKFEN/
Z5jUDsXlx1QA7Ul9Ue8FrbI01t9k/COZH9QgrnVbjux6pd1OixD8iCpdxNgZyaax
p0KhPxnfLBa3og+f3HBGL6LbTdOftNV+RElp+N85RONc2E6HZaH5RziC8zh/RdVR
fP2k/zvo/H0s5q39D73HAR1u5YkJJ5s5XBNQ3b/p4vEJFlpOx6uIVDlxHUV/x67F
FXMv/tpBwhseXbeBTqibEf2VfZHWCX3sMUPDdZflcqs3kMxKGnhAnUsj83LNaGwb
ymKR4RvQ/eIdQVyEE849TNqwfG3/tXxqXvg256TQIAhN/WpTcvaClEbaa64h7aVt
9WHZOHCmwlvFrA+k5oPCHlgUaSZJl0yvrCy318colSAodchNlJhhRcDxXqdJHxH2
PnOIt0JG8Y5XgafLroNBfp1/8qRrvLcMq2V+T0lM67tNi2EaV0hW8kVGWRdnsdZo
MI0CexZKfvBMd2VbvKF3/6czYhX6dWPduMz6nGqc0M1Mrorv/9re3vey/yLxZrDR
YgDjI27l1SonixRWEnWq2LsC3K2CRGv+WqvMp17nlD5+K8I/xBzm6+/vChe6G8oF
+sTXVGA+CoMBXQimVyKoe2YLNeAkmewssvd9az4CWlk+qaqLX6uoYAtD3Wavf4Up
OUpMO3ZrKKfjntdZTcZSq28mhSpv7V58Cfqx6t0iuvlR/bCr73/VLcLNGCBVzZ+F
7skPqZM/v8FRQtVfQbylY6tK16zrpp+Ndgq5hndTanEu1EbrJxWLw734MX+dONMw
o4oodT6vTz4IZIZE5e7wTYoxFKpEHWTJ5RiRKxn3dkNoamwEC/2dFze7bYrMizXN
msF9S6RPZngu8FeE6LnVZAeCIcMXBanEL86SZAQJ4eXPGnYQFzS/CjnbwU9h933+
VOkiqdw0H/s5pl6NhsOk96vWvAvAkfC+fB0il/It/ewBrGDj/Fd+GKtm1wonMZDF
aQeAoqT/4y9My6er+EN5dpeP/R0//CHPieh3sv/j0xV/gPt4LW32IqbDMfGXWH62
uZPX07T902f/BuhPm6oylminLT0XXbxUHjVGc1B3mXTZy+WohxGfW3xQUVXJSNgX
/hZ1m0Hsy7e/bIVLSVlgcwiPf6N3mDtB6/3UPCBVQOdfWLabu3FTxDRyxVfCPCkI
rBpNHXpljngWLarj+8panXkRaCK359oU54LQKCgV4A6hdPBrPOBQTYlQu98d/nWd
dBPSUiQ1wYsatrZCtt+QNNPzbyLJPBL32BfpSoQa2d5/sjXhAV2q2NmbNYR6RYfr
Ydj3BXpnesFUPqHD2/6jWUKTL0aC9aC92Xrtp6IAhccWdnhgeXyWdemakqngLazE
vD7ttYQPUDF83D+vIRYBszY0oEo9uDVbEfTednLSHr5/Oq3K5W8dGvQPeRFq1xe5
wXV6LMMOTJfajyq5YPSFJhN/BJVBOxVdxyydqIcQBL2lmcB2IfZUo5mLkbk+cRaP
7JBPDpI5AfdbVwm9zp0klHNcz3OBd9OnordIlye0aDli0HpFNEYf3RrhkjyQt2EB
zZNojmlN+v+WWSsZilbVhcgLOnrwSzUzlilL8IU6d+dm9YoXwKsraNWZrAHQXXhn
qd0xf+9z8fMt1KDByistjqSpBC5oTY7aZjPzkQH9o1YBWdoDzsBbLeFO0syeQANl
RW/DRUPqzNcA5WL0thvD9Kgkr52r/PyTPKvQYQ6e8yAacE/m8ZzHAUrI76iVzp6M
ab33+rTS02RGZhu/aeGX/SNcnxZweRYpTc5D5b79pj2ci5nJGaWoTmhHlaf5jhO4
fxoRU0p3EW/92O6pDgIEG3qjdZmy1Jt25eSVlLsQ20tw6zrJ2Iz6LiohLQu6jk62
k94aD6RCY0CaaZCHGb2ate7+J7mqufomlNrGSbUg9jx+qJ/XYOVxw3+MglWmJqFf
M0yVVgHAanxhfXOeyljKKN7rXljYrr3RAdWY65q6lrX6NsbeuwMQBHdxNc0cnSPY
G/+d+8ZgPMyhKvnSNhAOgaFIQjWDNjyeNaC6LEcN0r38MoyrLRSKkMG1yZTjuIS/
SrNEYHgWmUTAA24sASXYl4uVYcC5pgyIoovIEt2yTPDOgqbbmskp0aoEjwegns0L
K4gdiIG6qkvQ0cWhlQYOSi40jollyneQzDufpASY7yeKipHj5iI1uzl5lYqu8++a
xkIfbVE94+YYxr2WM0qdlkg/Sznx0STNWbG2MMGyZoQdD0WVQTw/d8v0sELVZXMF
1wm+tgn2t5Q75TR+W8R48n3wiQfOXxRsr/mz2CNfEKJ0XQxRSc3h2St8essSy9Af
OKciQeRkTaJtKEtcDu3mJNbHtxWeBvVgD9b+/CAyN4ezTa4gukkYo+2iscbZ9kQs
PYnUQ4rbnoYD5wG+SrViwbdALPEOpYGMV2cOKUYYZCCFceo5YHAI6jEIB/TSU1Up
KT1aCySJnWwMD6+h8RM96xhSy1MYsYCts9j9rTzECAO04c90VHIESd0/z+BJTAJN
iE7hqFulAFpe1agXn+IgsEgyD1Wo41BQ/jnQ5aBkEuQq72q0UM6BxpWv1fAW5yE2
rcG7XrCeGGx7fbO2qqCJK/kwvG3S+DQp8mVRG4DNpG5iu4NM2UdCIF4tDO5cIt8G
VvqWYRbyYpgbClZIUyf3QYB864r6kGpRpr8hR/6Bqu2jqlkFohNX5L9LKypbhEcu
R6nO0v9mqCEfNDP/9m/6Y5FHlGJCpjjjzE2tDEFGvi6iaqHdiUCqhP9NXIouzuQu
8BKGXJ/L2gWr20Yhfr3uZ5uwG60HItV/lL9Dz3j9I1wJ4eJMnRp+CI1KUzWehY3F
RK1LM4q40N0N++LaGl9ehXPz8RBDmk9k+HrsVJmuQNxS0Rfry632KXAOkmMYgrZC
0mpFse2Gnq7oeKLolPUU3FxVIzMql6G4Ny0dPyMJlFiJnfLUwJMf6dARDLi2DHFO
2N6iVPSm8vL/2bg+6zpq5oVnCDi13LntpB/SMla0M+VQYdh5gVDAmtX3FEaJn2j/
LQGi8rgnA2R1uNFnpVCgiNfQfbAvkvS6JBbi7/sW0VZWWIrpbJuLLR50eWFfbNio
pmQDT7P3VaFrg4sy7H/gOexrMqk5D7fkYi3Fushrd7io/8x4UOQlV6dFj3nEL6du
FN8orgGl5Kzg5y0jwjEvOsKZ9/Nx33l9ExTqdHV+ezr3YTGUs29A3W7Yi5QTI/9B
NkvyzLLz3fRqpyzTy9GYDgdiOAx5FGuohAzj+q/Bns3CueKXYI2110KvPYl15+Bz
p8FKBiJ9dOVtHnFtPsAd+CXrJp5GP95HrFgqYAaBo1/RDviwmyaftpaW6vZnUABq
Gi7CFhKUEUGl+/iflonb9/gZ3/HNRIB/H0B6oi2JIfspLR16lZkrdRPxpd+y9/Ga
t6kD+VxVpOOJCZoV65UdyMJtMpZDKm1ydY49geReXtLSar8tGNa+majHAevuNAKo
8Z68qeWd6WZJCozGL2ZvaKOFHKeLLwVSGxcJiq6mbYf/aHxXJ7Ksjcf95O8/vScm
GQspaRVJrJAS0ItpIqG6WyllXvKobym362ZlnRBLnOUS2Xrb2xRpOCJ588/G6ZYY
eVJhPPd0FkS/jUtZlzAyPDd9vXK2SZcK6NUda75FJVkUdkudRTF7uV75lrM8BJtY
m4WLGe7TsSrDQ431t1EDQyfAo+D1B/HjMBQLm9b6TJ/Ceqdp3CBdK528C32pL475
1Eiy0nA6gEQlDCkknjkIhivu5fYFV1RgNhpAq2nBV9esI277uEPUcNYIB9tYq+Fo
hRBeukR1pHCEV0GfOAfcBBG+zpJjNgTIGmzkXwsWEWUbv/T08AMWmdSbosZOIteR
WNmvXgzNoEqPhexVsmlKarrjPnEsF61KCGSiLX4VfvbMsiI13yyjjezju4vZSdJk
rZJ8OmY/U5/thMCwUlKNgU51UeLdsmPciju9+GSWdvKXySIHEJSbrpzloQ2d+CVM
eYK2sr3UeW+eUUPgrNudsv86qcwGQ50ufmIdwYp7PUM85hBBvDrqKDCNGk5JyVvJ
zQXBY60CCPpYd2vLSPBVp9WBUfdPchtfXXlBlIyRDMY4OnQJf8HhXV7pbvSA0HCN
in4nqpe84HboA0CPWQEJJYfvAeDrpnClYCzmkMdpUIlLS/U7ok+BTIsuHQJVNqor
XmgIDdr3x0cgcygu+8Nfr+D9n96geaiVrsWUfGQv8E9kIAl85WWRPmghiE0b3zgo
56HhS5ykwCRpQESQtvjtvaBnuefnQd9G9aa9w/j0qf4f/onlhC4PtS6C8AYAoKXq
/np/BUpXrE5iqp06mR62aHEjVdnz6VqL3axx3ZgOAmGnpFLhzSaJ/egocsQgr8R8
REQ6idDBD7oC6knssNs8K7p0VbrcLD+JiEtmL6NkK9th1bTL/z0jwNxjZ91OTMcQ
2F69kMOa5/cr5VivUy9/hTzNMIY8vYw/B4ZyYIyfbVI2sEl0r1PfAO50S41Es+/9
YYrEk5XGrXcFqaRtX0V/JosSyun93R1M8SEq2MR16Pz5zfjJEK/ohAXNFT99ABdG
iWpHZcros4GilaaR2Tbt43p0kHyWYSOtnof1Cdmt0i1VEke2MOOfzwhwKo3JouHq
ELsKtBnX71EGpVilw0qpBFHspTtJMgKmLJIi40cCUbIYz/WOQXsUHKVDQPjaj+11
IidohKnbgQTE+3I95Nh+s+pCXyX/9CVrEvt/lPdilhcZecPVW6ddpcL9ohMs04Sk
DU9+P9mctdJpJBSUDcJypSsGy/I5TS2CzZPCp1sOII8aD+RiAK1psAeyZ3Ep3nTJ
NlqmqmYQrr0Zg9m7q01jDyeuoITA8B0s4Q0fEBYU7KtmODWWwrvz9FhEE2lycfLw
WrmaHmkzYv4BLrYRKajXq39i+eyJWhQVT5bShjgaBYsAvJ3nXU3WMJjkqwbyv7L9
mIndcPXSRm2lB0nJpCuSrVjHc5NPHB76kqmNHNHqZcb6LzsMChn3S/1JiN9E38Jl
UI0dJt3567XMyI5dqmwSyiJr+K3/ZPtUNVmVBf6/gUIGHgXKcKktwyJJbPdBNWbE
XGlaljcBMsuGCdLEXL4CYBQeTw6QZSIRM4hXidzZ6A7XhB/A0Cbcn09FL9LrmgQ3
wIO64kubHm4puo31NaMIpwIY2yfA2tmQc6igjmA1AEv4UC6VDwFP301NxMfTOtpP
12jIkMDcfsVFpVobR3ytVQGggdWGfpBMAzcTPTg2Nc6PrWDjHw+DIiDpGTwLQmp+
+Be2MI83vRzQbkrEgmBS70qXoFD5EP11KcxVQDahmWWZFBrhh9hod0RpwgSTNdC3
SX/nNYPEaD4A3sHu3m6Zn/RAN3HD1Ww8gLlzCQxNinF77gcFBkUX4Yhhc20YPjM2
rDH48uLpD425VYU7w2xFsMtrMDmycmW1deAqA09Rm5G5lynPdC8jm4eS3RDJqz0E
QflMk973VmLBG5CcE7MDQwhGjxi0T8006bYsgXzm6q/5Fj883Knciwj2gEhNz0xe
ayErzzCBhv7Ld/MQ3nQQ5AktqNniNBaDuoQ4gaTLXLnA0TwVljqRdCO40oX2U3/O
yWTFl6fM7f9i2jeN460oP9M/YcrpYNo1j3I+/hS9phIv/9Galc1PZia86WvklY7C
0v5HZGRSfF6Vy778rc6SWqtUXlD6J86hg9MHGVK5cdlPZb/IlAUxI/765yoRzXmE
g0bHOOlWy8sUb6z3wUfgo0WauZq3BVdg5uYDMlv7F4PJ3GdYXeWdifWrm4LKzkr7
NwebDOGkUenI+jQRfGoXd7FFF/8dEY+OnHVPcl8e+N72a5b7k46R0/kJGMe+c9P8
2ps3yj7VjM+pCBWBoQomy1wKYmpe3w14TP9jOZxYBpnoyxKvcymT+MZ55zF9KjZu
hY0oknEQyf6eGCEETw+NQSCwYma0JxcdngNkd+wby1BAgoEL0oRnZwSRnFOFWZ8M
cKPscVpsFNmMCFsSRQV6J22K8IjtejiFzbfGtoDp4IjkD/5Y0xzVXwcUMz/Qs7RB
Nh4CBebXqe7EChYL0Fg0HLa0u1l8Jt0RRNQhInjViUua5zt4OP/vT4BuRoJokd6M
Czbw8OhLckIsqoVPG5oe9d2soR9aNGgIqAI2QZzp8Yy4R5gk7SG6lWgwJyXXqDe2
nOaMFOokrsgzRo3IHFx1qJ70O4funvU5ESYOvDakcl2T6ZxknzU5fkjbYMx903E+
SZbQS/2U2igiws9xp5zot5IAqfW2KkQFiQsYxjGglNxpc5bL2BnCqaLiXPytxYmq
VmGWtYb+0w1w1o8x1RuPh2zNxfPu1TUH8SrujwNj79SSuwrVpLvL8UMH7Lc8gogK
oGFF3BX/xaxSA8xsVMFXoFRFPvUnXacpyDVBSWbrR7MZ9GzJq7JL3W2tNlwM4Lzf
MLROSrFA6CYZxl9N7GekyCLRk79vgTE6HvO+F+bDTnfii2pJi3SbQIBzRpdlFAfS
9fQB6vBnL9Tz7l5FNwB7yySc5pJWUNs9jZp9sGyr//czbcD3UXzWWyTDQwrzc/aL
6FEqCFIo588f1xEBRjyQ5WNJMn2goXw/RVRIHM49uNiP0xVqj+6soOPrthdz2o20
VGmU+52nAlpYADBTbWv03D/MlH33SODctmTCCin2fW6suZ8qLi6ConhYn9rrXold
YDwoMYHe3tp0Djs+KfQmmJMwgZymUyVCf7/mAlHOQeWSYWlnIzSqP/oEGvVOUe03
SRzMnw0ZkODL1rrEH8cD9TFLCFlY80bSh/0iEWLDUaMZEu5+sRAVXrmYlj0800hX
+tiGyvx80j+pnYJ8ST5QE6blLJuVdIM4ds3+I5DTmD80ct7JiGpumSzgTzwCgeFl
kPYvPEKwjJEsEvyiVG0w+ec9WnsQlNr9YKkkYhKcRKZAM8gqkUlT1pQYhsAQypyC
Ze8n3NEoagA+qjqVKmHvPWKw+nfDd3oFMn39Uct/PCHSPJRsEsZZXGjpssMUPBSK
YzdmFHLOpdHdV4VoZOeQWlNNiKa8jk3+Xu4+LurZAz6CYPBkkhpX2hVci+Ezju6H
PK4vIGLAU7x9lEFb9X9klywg2eyLbtULLsXvOlKieblmmg8V0AxrDI1a+BYvaZb+
6sx002XgOAsP6m5xo4P0ICKOPr2Y6DXA/3dh9+j/DDHJxkr73hovznFFfMJ/amPI
tRURA83tIOLlhMRz+NNAcO308mdYTWbHua7wxgSHDyQ3YoVoy4hvBg6QlrZwbkcx
X3ds9DeJ7EMl+KrtD4ykOj8PyAdAgFxRHHJEWbsBRCYEZ+Hd0rpSNEsCOV/XmdkO
ytN9rrgGz1w9g+K76GBysUS+6gOZ8u7RAXwkphsjeRK4BuWVeeQ8uNMdbIA5XGVl
S//d97ojcYcfIECoS9RjZnO8l47UCmjYaHqnEYAnfdtc/prembWaUSWuEzYAyLRO
8sdDBbsWSLCK8GIqukB3C3fig+yWBtiM7BOQYZaWkE8BfS0NwSfZvz/A8ZdomPlj
xXb4pk9DxTHPXmgYJJevju7/LZZw9d7BgWx1Ubx97LlgHEXZ4xNj/e67yYb7O8kT
55MwrpWMyl2r7CztViM48RrVjPVLGioSUzzcAvFXkKaNIrQ0uoTJSxonATD7KeBi
ZLFWJQ2mIcTV/6ZqEQXC9rvXDy7U080FMJO7QSrZY8OVClQpELDBYDaSjXNFUnhs
rvsKEVocCXHrpj3iFIYa2VBCBzdYpMDZkupkXdUwx0Vmm0mG4M1SxOHMeap11K0b
lIcQR6x8s07GxKUgTY3REqvkWQ4n4wUX0v8FgVeOTfv++ivgE1GAhlcnywDeO91m
8ZZXXOgUg8+tPt+1V44tR6pTYpT0n2nWtO6a94nlGItPNV3iuI/E4EIOpyO8EXIb
7sSdAseXqKSh9wpZ+YCm9wye3K+ej8C/gL8PxiQ+WoVW22Bcp7i1Pc0JEgyxZObS
4suftj+9TxVUYHheqYW/47rU5KVlZPyMRzHWnNZ61q+j/bFRrY33gxZbo5vlR0cj
5DMwj1Vvs8/aL4FLrDs2SLQ8JwJf458mRxu7YTchXcFelGwwdfgSfMt0rVFOU67E
rrSb3BULzztE3P0OBtvOp5G7pWbKCMC9q5KqLdWtUjMAJn5C85e/dFiSPH26bRKo
6dcTobk5YbOTAYa7do4E+MRfD1PdebxGmGlzTfp2MNScdw5XpIi9HDQtPDi9t5p5
sRJA2xc059BA05oRTFvnLhIwryvo+ZGi+8vsskfShZyShOeztSEeGYduCJTMLTcY
oqH4BmHqGDcWhiSZLkTl8npBNIXXnykpUG0H4iskU3cMfrczJse6H2QqB4yAqEJh
9zm7FCMhhbinanjPsAZ210niMjC9mrF1V0VfDhCU5NrsPqgjq1kC4LCNUVDAi4GF
n81FwYvGARNIrptDFD+4J5iULvvu3s/vBv4DhcB7SXYGm5AMwyl0atQ6FHFkfl8s
zxgdFK2KLniUTBNvM7yOw9wyGwSxZW1QhgQNnN2Glb5JxCeoe9ArYtnLzgv9KOLE
4cMeHmpRxv+dmw/XFa/cdY1j7H/eNz0jA+XBNVx4m8pXE688Z2ygDA/Gdl0OA71D
XSK1VTTtXWZR0WR7qGhw2mDA6FT99Adtu11fT+kXCbcfOIKwoejdfXNE81rdTwrn
q5GESDpaoEPwT1yqs1gh4/6kBK4pEsZT/RZP1tzmU1KbNTiViuLk9wyfej8ZBo0P
LOF3B5mQd4lYto8F+2aOLX/lqh8oIzHc2ed1LYpsT7shiquKQ1vqhQm9mvw0h1gj
Dq3NxDnBDwbdTSp66xaAmEkiw8hEGtBSeARFd64qwb7glAj/IyffuAGjsqbqcFyv
A7J6QNtvU7h8jnssbqHTGYKz4huYnacPrAFfGj8nVLkOI4WUicuRZ45Fjv8zpJF/
a0JPECGZ5FkxT98MUBvi3sxZdAFOH7Hyn5JxAeJM/ayHrZwyU7SYgjomzwzsWgJt
33wKZiBo2w+88UtnG3lYXPtTQ9iH5BXKxnDW5IyGIWvm68oSfkTZZukvUqFA6HVB
VqhdDMqplmdF8evCo5ao6dG/zvZsjSqW3VzFHM+yypIC4rURfBMbyv2F7fsBftyA
sBSObZjIXtPRhoqAn4nsJjLxdMY4iACQnqtESUagbovEmwMeC42Br+eM0yWlhB7D
2u1n/E0Xpt9duyfc2doRdjMVdOuOXv9mPsm7ovhIwuW0WUWSqxkOP9vdrzEzNv8A
Eoy1fr1fu248EDDnrjoT/pEZmJ7HdQ0KzAGM8noaPD7HKoT1uX2k/FcCXbVJlF41
RPwKTz3SGbjCzoaaesknqaGh/IVZ8J/+LF/R2R7mhPfJ0Q5gIv+qKqzRNy63pQsB
60RotK2pAbB9muPavexsqZl46tIXQFNYlrRJupvxOxAxWNN8cHWbqDjR0TUn24Ps
+B34mt6X7/bk1eBMYSMchhkDDWznVG2pnnZ9Nb5FP/tP8Ab4+FAnKEFXHIauxyLg
lWzGRwhXKaFFG/splkyOQGAxytRwfCGw+hjgfW3cBXUrMbJEG7Evs6VbobbOTuLe
yWm7bppI5o7U2XGMWdKdqSnYbxdQ7IvXXV1XGbPEbtqkcz/u32eHS0WgcP0w7pHQ
vq17Q8l3uFQkW+4YZWQqB1s2nzzHr0dS0/lmjlh3/46V4nEweUWHvdH2j5ULvnvZ
jKPuGTF1FFWy2GZ3w3if90MZ9CmmK9CjxHv2QybHPgt1TjDC2+yvkioDqH326qjX
nck8ByItLY70+Sei2J7hGNjSPXQqD1NKC67Emo1EPVmO4ut7BX+GzuBzUhbiZpbe
dNVEmWeTOzMX/I3golMwJ35w7/2Tm/+ilI4wcHXJig3AcBFwIASKuTfJ320Nvycx
YYI7yXT05M8JbtZ0dDbtlmI5DMPHIyZiw2q1X4CKUvRjIRNPVgOZ94oC2f8mjUZI
0/r8a3AkO/ulwLNSDo049dLImFrSCD7CSZkvKHmfnQUjo7bliVewVXnFp6+FOE13
GMikLBHJNMaydx3w2M2Gus4SOcYwGjNMNw1LfY7MFVvkdKllpk4wCh1YDh3A0lI3
bVN5d3lQpzNGi4eDkCKwuNK+GGs4OHqxsAomOJocjj2JCg5R9OcJRFop0B+kKqPC
WbJfSBUH5M1yY5nV8HY3YcjjuWs0JO5+q0s5K1IDq6h9GpaEJE6Pbp4bZkC32X5V
2Vy/2FHt1yD/jUr7jVBwZZernH26FOZDg7ji04yK9+oinpjaUbrvrMLu8cs635N5
+da2wvIq54FSsbrBcP+UB2zZHTLRvaWMj0QLIwSy9ieC1FUffguO//6o/OETErH9
VicVYR0WQJtGTVsKrTEB8fb6f4aXgrhRfWlF9YtdDnXCDDx+ZdX3ClCRY78EcsXo
jMQ5l5PoZxbfbLZ92xbI23DkC0UK3kaYJPfLL79iIgXdZRjspFsUv7ywgQVta/OG
LIOq8PjakrdEnJjEnGZjCG+GO/fh07n2V87tjS66m35Gl1V0iNflCSJu9U5Ysive
ioO+nRLO4CIx6VjjvIWHdGMmWIbuBbtOgjXpAEb11GZj02QYpedN+F16XADvF+Gt
sqT01cQ4L/681AeX/k/DhLZ+24ARBc0PcSJEVQYFwhB2yJAw5pulqJf2Fp/+3T26
4jjwqBmyYV6XqlFV3TsMruCII+YW9QlCWvmiPiook1ycCQHGOzQpWi98TCAxZdve
POiTfgIjVwyd1NgUUQKh0L/bCmFfTNQXoAtWc4pM2Kj1MzcIAnqQ6S++Kehglrwj
yY5HNXIw4qspYnHgxDkzxiTWSmQXZg5FjLBxA77rp5pPbMmZ3LenuYGlcy0VDXYw
vqUoiPgqns7m0qRM0lYFCtKAHh+Z/Sa7RK91eYxaZ26k5EhkfSkaQzA/tAVF8r75
jNCbSyAj9TS8WErNUrGQTVNoba53Yn4UGa030XWaWZhZr7IeXXpK3nAda059DSmr
EF2b48K6Vt6kahIeKXioDybZ7aQlBkmoewiSdjuzRXB/plI+IMMHwDj/JEqbmQ9q
ZAd5TIua3LIyh9orZdXcqYAM7AQDnizyxv9WmfQ1rO64vPHU+s4FEdx7f0IoyVz+
gLt2g6sAIUt593clAHSMRMXBBx+Dsatm9HiPrsIOJ63q/YoEPYVRjFU2l6ZS3lVG
pJM+ULS7qxazFUzIzy9uuPSbfyzIGScMHCwsuk5qC41z3/tVneVq3pCLyczBXNo9
3CbRF91V6v9aZZpzdWONe0yNGtH5yNu89mw5Tf97b0CnnbAGB8m7V46U4HggyCJm
PhB5slRf7fH982Xb8dyL0S1Uyzg60XiCAeCmTwXb1o6KFLrL8mZIT80hv3vIMLuO
EzPrs9ENOh8xoYewJdIsgZSSs7FkjYxQroFe5O1TcngQ/ZBKh9wBGJupS14ekubA
yK3C6q8pDkRMxkqxj6hSoZjzzQzxI1r/nibxHPop5lygNgfzAOPgKde7kKovDMpW
DIi/B9al6mWWccrwnCfnXa4FNstvtjrma2gi93wMByWy3BjLrek24G9OfHQjU6xJ
7hYGOvm/e7caB9GMvpwe76x82pGVZuB8x/IkZQEARWfCQOxuhV3Bp3arH8yOcfNZ
Ja1qasOaBdH4gkPoQle7kIyUaGO32aJESUlfOOaxRYeG7jCFp5nbWsAnnk5+7/O+
6NK2+V1CTtnPI5gsvSUMpXUpa/6GN4dYTiVhndui6czHRIlEfesHsWRbSK0R+iPi
43XdHMXx2KnOsixpGzippAsgrogwMZChFi5aOAG7GGuyZ8Vwjp4a5SV6RqspJb96
5QRvpwqXlmflB/G0JHWcYLoj0AilUnLLrzOv+6IDmIk5fJ1dd815XxxHeS/9ahpa
PMm/5XkP4BEVaBRCjzQPPJ9RYlHGdfjHpo7PifYPrBOdq1c/zglN5+Cu/ZFXZZVg
XEGGTg+qo7Nr+hGVYa+pO756iq5zElOvGTbVduFU1aCYicK13zTSckjCtxbRoOU1
CMdZICVc/HB6/qmcuTWE6yiHzjB7mfP+4GsPgo2IQjttRzdafzNey65BNLHZMtNC
eQ6TjOkHdkKy025W4pvp0sYHnr2/SCZ0Ly/uNXsxziVxOt1YoKkTlLCvlnWZCyfO
jObcnpLdqnYu/0OOPHXBpJlnAjjC04BWITNeRRaE+e0mkYoVvCGo+olMpsHcdElK
2QIQwOpVgq01EIzwNe2wb6HiaQqqcAgDvQvQUkxRF51P8hJWsQKysm2nztKMRvJo
Oq8Ij+yM/7pWrtHytBrNBzECm8JUHHlnKmYXmogC1p2i0/3mjjiZO4xpaMB29Em5
QE3xF+xHqGWcHDpI0QJe54KFrj20LsFqJjQnvMGxXUsTTVeY3r1TC+x8Lr2NDLh2
cWN8paHJ1wXxCvM6z6fw+E7NqHm+DaVx92WMILdb9JRoQjaiqGbCcY3ozrzhR5SY
C0UcIWaVYrQFNnA9NZpRmwTVMT0QkTc6udFLvTJH0x0p7tJ/g6tx/UbWP6BTMnGu
37RVEDoVVPSxL2Z6tqc2FcIrNxcLXqsNI9FDSsaTqTgwI7cq7vTc9iq9qV/n2zES
1LJBy4c5BQCwARfAeB50LCWVmi7Y8vxzcdB+uPPY3RNDvjMGCGMaQDJ+moKM0/GH
lDER74DPQ2qq0TkiLyab4DknupCIM2fJ81Qw/W2cYFsxJnBOYTgOgOz+nIJvP0TW
WJVrL2vmQJySZOJ6c30E5KT742O4hXjkXDV0UoeKuL9f0nfSKTCTwB2Fxqok+h8I
sYCetRwB9AQa6iWGDHK5ED/nad3AS9CX74YX1uI+liEUVDbMtPdH+xD04Ipn+nvg
useNEMP4/BJ6QE6IWJ7QSdHe9PzJjHKW05sabYh/z8ECWr7HMDMuCMmQsqLe/0hn
Gklu0K+jZLh7tPwijPNhRF0ZRLsWQWhMvxP99iD9jz2Ypf1G7wG1hChUEGi0DBNr
qpoTIs882k93frMeTs0HgsO8v74zOQgj5JQR86QtRvcas+jiP2/irxrgJxYkkOwl
DjoEDQUy8hzRXSBwY49Px2xfPYUXc9dGE/3KpeuexHzzb9mJjxR7be84o996MlVn
wvPAoVQLGyt6/aQhkX/DdEZp58dJKe24uTb1ImmzUZ0hitRs+GNpKltZMzQtBvk/
Qw96sfNIRVdKbRG81WJR7h2on7JxBP47stoUuA6PF81HeXcPMwDVO89aPIYj0yHY
pOZYQ+zTF6vL1r9vxfSps2ksXQnVpg5yplc78XUECvixV8WE6HaBpJ6ihUBj9BSv
LAXBN3NlNQmeQ/Li655vuD4lf+i9DuLqlqA9vjigeY9KRopkpdA5I/gOVnorfabX
CQJ3O/Xjj1irus+vXS+wiPut7QuIRnz8ESKfOlVYWZK/MUZ5qoW7PVo2DxMclD4t
vO9Zg1z5X1CUQWseomcpI8HRyD6OEKTLsMs7xYhrRq1CnHc31dkrgIx74XdszQev
CPK9qytlm8WOO/gyTXc56rim2R+d/SH4AhdOugI3/q0eQWgEfMz0G9+Yp9EFRZWu
d09iUfx85y6i53TyZvhN+aDGwqdKODRCBIJjQmi8B/IxRyP1l6z4+1rmXuByUSMs
q/7KjcsC+fsb1W0XpwepoXYcNZEwnsUO3lByzeXwTB325S/MpcidU5XS+Rlf92LS
DCWDgNh2eGnXS3J1/qL5svOy4v+66j/64xCltUHkSqPMeKprdcI1Xau73xG7EMT5
a1mEumBdSZBXfGfLwBFuSZDNxzUDDFZ295AYRvAKTXLSLQS4BHnuCQVg5y3eXP7i
TOvI+3kapjMAYxjEKig+Q7N6LMTrGFrKDkmTsyEOQJ7VGnMN2xreZCrvF0OKGro0
b3w4yQM09gxI/tjVrRwthjnJvhygU0x7Ue+yXM4Q+6yvs/8RUoEf9QeiSdUdOYsu
i4l7f+pXc4NK+70R9y2cSMZQoUfhgPpKs50QmiC2durbaTIr7QkyKrKBig1EwtuG
tekYYUH0FfSA5CMgZpV9QSmCK9xVoi2wGmuq71UILyc+AKGi+VQYWcQLLmheefcp
LoW+kR+2YJCmHL96h/wLrnXwlBtUGQKotFnPyO8qaZVYFeoM5aXRF9U3YTm9TR4O
SKufoiaY2XpveXjAlHVR2bEzAEufZPBttxDXiWb9BM+lYrRca5WoOC5GAC6VoTDr
ls9V/s9CqmdnG6yNsQu6Fvepy9CKtr32YrvRimk9QwnDAd+a5EEbML0uv490pJwn
45xWlFoJu1UrujNsxK+gzGZN2PQYem3AqecTFOat0Juf5q6SsGDnYAJm873kFbxV
ByvhPLH2zVV77Yo3BgVb/hqNgkKy75rzRygXXHR/yv09dRG7crlDh7hK76XxymF1
WAP6PiG/s698zvdLLPRDEV16LJYUaL5JcJl17XlFk93nbkwnTs9bXLx0jp8x0f4a
NAsPvGvgRjoKkiUDK5YqJPj3iTOb0WuJvuYk2klyGI/wkObVDbAA2dHWRKAaUc71
6ZS2gV3Z46T8gLmZ5BBFplg5phefLGyjlRJmDPtTGiwMSrIfYPZUwrbmIXSznagi
sQ8qad/xeK7wloOUCaw7MEea8xYDEM3qRoGxFGzjYg5lqAdoVdR5JDSYoiUWsyNp
Z9Up6P6KRBdVy0vwBSNu6DpAABndkOkH0/ythFFKNxGPugNx+tjb2hlJoXuJ848p
A3Q4hYd+NQjoY5O3gMTHMfvhZi7SFZ9Gb0TrhlgV9GF9J62PNYxdVC5bWuERVMWd
jS/MngKMPXh/kHxRI8HH13El3LZZRU0+2lFW2KiReNE1CVFtdOby88LJ8/99xurH
01i4/V1N4BU5n4txPQp7F8oOqxA7Ue3ZKffsAviZ/+r/0JwMw3jT0Sk1TV30gebI
hEyhwEMP/Ys7grKB95yPJL0wEYhWajALoT30VisF36D6e7cuJ2bFQAkzVbDj9pSn
p0cfZ+Lu/+eC07aNhdEOXiHoIAMpsreV+p2d1Y6nfF6vGW0vEOKtg9RrvuL2DAZ/
Anq+Fk+fchIQbpFUi44Zde+3FSlJxtBViFTf4xWNGmGDQuN3+hWe68g5c+BvACoG
1llj5C1hz1xFhlMdGFA4nICP94LXJQXiiVeCZP4Ll9KcM6eRu/ibkHqhmwFrN3HQ
h7MQKwu8fEpSwOoJZhcXRQVYEXqAg+SJ2hER46WBkeiSoFpNIVGgvHUQsTFuAcRu
iEUgXuQici2gMXxDLlgG+CiEYyNfrCCgv2/4BT2W70PIB3Y23xPBDW7+JECfVZjR
mq4xlFBCTI18rA7TGq4Y9X+8FhfqS7EN5dHX8gTOeODScMhY3U8l1wLeQ1mRF4ca
iCkckOeSIlF748Kb28KtKWFNNFZzyyRy1z4bHFIqFUcmHCxzCS7XXy3YY+qGd4g9
Nbm/d1GBDNEcWrjFHLfjgu7P3tGEktp2167M1YOYOdRhdh7rPO+kLm4n+aekHdCT
5uExbVJUbfObe4J268D/iEs6EmtBeSJGglf2SsssdASR0SfU3EHSjNhUwFSbt6LX
+vCH+GS7DV24iv3EEXQ5iCtsatQMnWc5iRAsV6QZ/yEDKhjL/TZe7ee/To8rPtUl
TqEY7aJEnTYF7JXFqh1bSemf3/I6OEdAbIM6V9rqpYUA3Ewo8P8488h9X+O9XYF4
1bnkbhKGljVDjf1jl/umMfiTP5pJnaifazEIQAUNDQF4NIGav06bsd0ag5nUb6Xd
N1SBIcHModbprrXy62PHED8V+0KR1vSZgQmWHSomDAZ6vAllY7BKW4d5oh+Y6gDm
eSxy0/enqNoAZ1YOPXEyaVC/saqLziPluReytGKq8JParI89QQdUx21c4P5DNTys
o/qNx8zhzHDfZgUEzhTW3OdVnjgbYLURmlqlVOsm2cQ3oTPC8A0aR0b7un0Q/8gp
2ZKEjrdSfoSUbFm0mZDD01ZgZAazXEiMu0u99HyxCNH1c/q8K3DEDNqPi/hZfGrn
Twz28aQ12BpgV9hVvg8fFkdftrqYIO0dNCkfXkSPhAzdMjghq3fbv9V04EvschVd
3BjYU7FGtJe2pFQ5l7XpHzA1Ramoj0zoJtunAOU7Ht5A8dhY81zwRYd2MUNOwh1a
oVPSMnXBmRDxt4kdly0yMIbWPPopjw9tAQNyOxeQJGdQLxenrs85yRHdBxBk8rHl
MYZgE1ZxcpfOjMtZ5d/Bk40+/XwSveA0l5WgdJkRpBnDEm/aQFzit7SstXP+qaZ2
+J7cNl8RQkfLptSwlq7gIRTc46R3xYMdaUKDwYkGtfN4AtcRhXoXb/WVQlv9iDPl
6ejtSL5H1Eq4g8x/MNQ2X4hi1Vqwti/X1CKZjmH5aRZEui2xng7RDnxToaMhlZG0
wopwE4sSy8VLNkvs5+RemfMbbmdcqMntGstxCpW6mr1hIgTTu1N2i821x49AfipY
pJn+2q9w4vfixkRQtbwT8jXql3pezg5sT5PblC9GG/TFnr+E9e+eWhipdV5xAbIb
yqPBa0R5OjJGTtQj6f7qvR+xqiRWCkp7c7XhyFpRSc2no87z1oEwBJY1/9YeBIW1
VTRZdCqQvl9smWgXN10aRwHCUg1sa1fTKKHOtGJSvWO2Fc6ioRjdHoNqcPkJC4Zq
ElEmQ2h30WIctCa41Ovcl7YyAmoMoccHWUbLc9T4oOooTyuz3xYblw7Rtsc6FFPU
Z3qjnEavBpq1ZBWzr0PJfcxBhq9RoaRO+n1IozOspmAI3wgaviAobWgtjMWh4oCg
GTHokBmt2Ts3HTVI/suYusv3qyjbKsIgFbpivUzUXoureesPayTcgawu1gTf94iJ
8eKmaib2Z6NxtQThBm4nibhLrhGppbjUFDa2eojrHtmgNPqaev5uOgm9QL57+LVU
klAx2E6BRQt68YjKBhx884jI/nnF1lo80I7KVqrJw8qY+SWPAhSSaka5qYizK8+y
J3TGg/SRWgGwfSgjZgrMLOHiAI2NbYzIbRzRuuzbj6uR60xxkFSgJ82VLfPb6119
RF23CnDnRn+LL8MXDJTY+wCcC+gNpouce2mDfKw5BrMNVvZZaevfJFvAj4hjwr2D
KfkjMbugby31M6I/4t2pHTDI3l+SeZDcRZ6zX25ooh9JCFgti956vPQ44LOn9jMG
c+8U6AytxPi3YC7q/Ynnm0E4duFNwFeWZdiylBmZOcC12Tdax8oU9yb+Sqn1K4CM
fb1J/cEF6OPsEasS3Bivl0pNYPikTBbtE4tUITXDmM4JbTw16E9FdwkT1XaFjs6K
8lUAklI7avvUUqE5hbQgsWmeHSzDfGD2e47tE9JDhEMj6a1w9FqvSxYAkJGv0el/
7oqBSWD0KtCwHh7g9ENrY65wQ87nPqKulOiHpZTwTTxkHzIl6xUZp7IfZpWmY4wU
irqKb5QtTzii5ICnPkggkkb6ktjmLykTDa5iSbAIC+2Wb+PhDsR0jMyOD9lUl7OW
yxDoDkvkdDxaVA/UT//xU4txMybIEC5dodRRlPJsCzzTwqcKML+9oUV+rUBZYKao
U+mpA+vUNeCQD7NZJ5h+HtojF/gDCSnyZtnDkZpnKrmOoMKh/467e7ZXCeI3KiA+
bJsN9z8X25CgzX7AuqOm0R30fwpM0hqGrD4Wy1NCiO0RoR3dtYUZXcR8FAxlukyB
c9dM0vcV06PaGYncaZ5Mi+GIQCuwUPx6XQioGZE/k68j+gT3dEwnAE2B2UnyDF0t
dOmuM3xIXtVvV8EZ9eqrhSE4QwVdmF4toppCiZuSYTPF9MPnWBD7aDJ7EB0Oq2xo
Y9qDD1p7X/oUdl7IES3exfV4Y5327K8nAnXSGc446HuWbgN7AO9NKckX5Q8OUbQn
B9yb7vx5B1QFo7Q8PDYZFM0+A2+u+t8QMB5Z63w2RHx9ZPcyzWTJAczOnsK/RFjs
9jCSoT2FpT4OrH13Jtc++sH5CKaWIuZYZU5dYbi0W9gEF9qrb6oosso5fYeoW+oS
65Qlm5M++0umBV/n9u/WMo8aD583XxnDp+mIUeine/Hjo5l3ltp51W+HZkqJgfvj
NOmbwM1Jbn+1EEr4KjTV1ApvKFXoUitJCpE2CsFAB34I5M2foNmSC5OZk4KsrOnH
xY9wuRWPtABIog3ChyRUc+JlAe+/CbfoIE/bapUo2YdZJqwIV3HrIfnPa6quGrhg
iaF0ycU3sgIWaUKN/vYtKeR/q3QSzQEzIIXoHZDU/ADah1dq2fczU5pWNNGTp9rP
wfP8/Cxhg3Uc+Z+G43gFxgIUOYbl0lN6Q+7FzQ+TgsvcpjBRO2znEGCV6aN+kLvv
ZMH6mbRDnGbrh+PPYNwUZzXiLPxWYNjxOnV9cZED/F0wD3dzzVCawBbb6JppdA3W
tgysRq5R3oxdroEqWdWpscIlYXqMKUUCDsqbvUSCiSh18WbULINCsstch9M05/02
iXrjmOthS8BmAv+H+3AHq6gCEQtEeOuOy00kG6lMthME0lJUcdZlUoKvOdxubtgB
DU7/yHRIdpaK/r4vy0qhENE4/UQGaWonsIYDIXbvKDm6hbUmTYr+ZavEfYOKM5CT
mhxNd5t9wRCbj3DJeaOvphhok/vDK5pFkVwUicl9rq+j49QxYTDxcWxcAEYSh2y1
OoeWETPTmoSGXPVXwzmYjSRka4x7bOocBQFiyVD5GqDlLCxhpcEEp4qZZmSDXAzg
zyZz+HAI/yZY9hOk0tFBQcGJeKCVU/BkYyTnQYat9OQPp81aN/BM9XtJmBtM34xb
PTmRjeIFK41RZx8PylkRPDxuFN6JAIzaU0AXoFBiJbqyOSBx33VhWqnSAHSALb6P
eulekxpRmiljTAD269XZ2kG/s2uoivUuPQeqqT+bCuxl9b1UxWVofIr8/+FRaLH5
CXPnDMWmAkaOmiB6taZ733kB4lPWpvH2dXKcUWYux+oALqpG7dUNiM9t56X5RHAx
k7Djh4XZqN1T0JSymCiH8+FVrLmWYIesvYmoHisdAyCvRq6jkf4vm6XWuVUBjBHW
S5kILPHJe7Vms77D50kkPIQUNW12ExaoquPhzZv3akcR6AiHSWtMZwD5cXULV6ZW
Qc2ydFbjoBHoPeO9NvpUM6npHgg9yl02g3GP97xQ9zQ+uDwJi1DQcqz8+iZnt2ll
XotJ6W2oNXh3MM22EgN0+UWlagDNbKxXAQW2Cl17EwIc3u9ZUhwQwW4aHFpaBJ4F
dz4gmpJD7soYS/D8Z19iT6KkdfwJff0UFIHqCQNicd9DSFOEg01dx9Ru3p1Iz1TW
btMm8WJmVFewNVLISf+bhUlCJF9wQa2SCq7JEwaw3jIP6sGvTU1SxlVOUI+yi8GL
AA3D6WNiRNEhgyXvxQwkoXIX7NBA38fJb3n06DUF4nasLDAqDG4JwyNTS41HtFiY
/3bLlyYhjc00mdzMvit2yAk3OreYVPIPbmlNnT+9tJs56Uyut4DV849X/3ucecya
KdtuAnKwj9ogDmG1cG5qBeJrueyeBj0Owm4IQILUSEwmyIAEbivqeGMGQz1X+6d/
aV4vmMKioQl6y5gMyvR0wgYNmHyuiiF9LAj5uWHnP80cznKtSq8mAVo2YAuqqNel
nwyRDJnn/f5dRrEjUoueP8p/4DlBa//TalPuZ7gSLFoqsCCCzvHTM6zu1tnx6u2M
G3suHg8AboxgGhtrKEf/kpRIWlPTaWuJqfVaggpubIB8/JoJHaAcOf8/nn/Dm72T
RQvjz+62SNkmKDT62vb9DgHB73CPmBlX87HK9/ghaTnqQH9qbxCSxQLlfGMrZQHS
EwW+h+JCEzhxoCx2O2wle9+PtuezwfYPvTy5RmHcuYjm7n/dMgIanVNX/Fl/bLHS
N1YqVVD1aS8W9GGg6JQRofxCLxf7Y7tZ9dwAGFhqrSCTakKwr5rDYkCQLGz0rGBl
Vyi5Tg0mvbiMgBYde11o6oEfTDDL61b4wVeC+w1VudQ1V/FPD2E9QqJPQsINBZ4T
V4/TC2lhvlMKdekdCYRepUNmjskIakOObJMtBCLYIiGzIT9M1BPyU8eCeBgScuUA
GxJQb6nLnjhrbYfTUv3rjdXLszkpAvOrSVf7tbUDA0iJQyWB7FR65aAgpA8DtNW+
ZSRpXJCURxUzzWGK9d/GBQa0Q8NfhQOADKyrmOKJ1YOJUW88t1qJ0lFfP0d2e6EK
FWskAgT9FbWR93JBWfFh/tbxTTViIPnFZHk2kidMkcC0ZA34UgQ/EuHjzp/01y23
OXaj3sCZvz+6NyRbNxUE1ZhIeAq/fRup0o3UAz0xrxgoRHzk5BIuutvIXEQ19Sdu
kIL4KHC94yXSF5nsj0LIl0/MQGm5fn/h9swBENkCS9wKFqKuLCEXMccv+1azQ4uP
EvFQynr/dbjbveWSmCW2AUD0ZDZTWuTC43xlxKc2AXQ0n3zBOH9oLmjOdoseW93R
342yn0iO1azqGdT3a2RG6pTWw/3DfozJxcbw69r3Rhpv0rJ4ndGpVJLdQxv9Ape5
1grv7jsETI9XF25eJHoewXq3x/XP6i0XHlw5y7hW3RLVwNZ5OOOA4SJavV78hQ80
atyPYMva5669Z+9gkNA65MtJozP5WvhAeOPu0JHXeN8QnbogXep8uHc2ERJGblam
lXGyoY2GBhSC7AOC7szrl4I/hJ/Op3xGL9OsOwKKOY8zADTJMmsznrSlEtdQTwuX
pnJQk6SFOjdXpcj4WbAKDGPUS9uOTuFNtX+szk8RjYbs6yf1bZH1tg5npz16F+TJ
7UVOpmXHjrTVgIIoPamuUb1/EHha2tlNLPMeBeM20R89sncZU6J/G6QnE1jLEjzd
jijdg/VH3WuR/YK7kf/759KLy8+vbSXCQfA5uUDO8yL/e90oMlFQA1+F34Y9Duwv
mjCSTs+BJ6LS1IC2+C/QdK+oSvSKNaOX7b8a/x5cX/WpGKKRsbL65uDySaIvWtXj
PAZsGVThjc0/6z7TEUbnawLad+O+Z3npu/0MLGYQ79aS3Oza/Nqb45o+/sVlQ2ck
nFrhkKLokMTGHHyjAPPezJCaPvK95zeieKG3QG79NVkKkdfstqeyli7/TD3n1A4+
ZjZaGFEMB4R4jObxBdLp/nA+0cQR01GQkLYT7SBVgyJoZyQVxcQhNmSfimqop26F
9D4j7WloZcCW9RLumNYEJYZnS91YmaDlsjOwC3/ZNiA5ziPjnbkyNogdgU8KEKTx
cMICod5KV02isKeF4RVyJ7g471mqDgAALEueUF+9Gxm5pTw9WqI7rFJyb/xKP+EU
oExww6mBDNdhruV8beIz0rDZ5U4qSuKR4pZm1jd3hp/Q7SZ90g2QeA7+zyhMivDn
KPYnCunGbSgOGjfALrfflBCvrnfJ7WiLylIJgXNSBW/dHib/6OSLy+hH5C7iLfL8
lukpNAAJ1grVTeJdluLVi43Nk164lXSoUM6AnZR7pMauNYzQgbJ74/gLCRIjcip8
t+3DUpQc6M9Jy9YypeOQ4LYFCoc0v4CELsnV0IEOdI7U4dXoWKFbKfnmeXZx910c
WfDzibDjTnLVEWBtSXpUNPkoSxZKGcHW9dv2vDcZpiqR6cAChhJX7YmDRMkQtEQn
uFTwFKi2lXMj/jIKXjf8d9OdkR9F6FV/w+EInMXRhRqUlc48y/jkP32OkrWGpa5o
5/0lEf7GrkgnRymh2p00xVZjcPQFxWXzdlAmbgq2vEj01JiJVzkvUmQjLthMRE76
nC8nt92MZLnsq99F9ZNCEUvPbQveSwt4Rl+ib+ObpNg+8XAYULoRDAwDnrLDPQYV
h9yw5nZkPo7cwVjUuUg0Iqp3cV++/V5Yj+hqN3f+bn+HviOgwq3HRLhHcOIAFhdE
dDKTZQ610LNwexS0Q1+GXd40SkIJpcgbcPEOkbLyWpK3EVG2m0IZzSGZ8RtOxoc2
w2otw+/rTkzfG6mNz9TD0kojJIy1rKCJgx3ov/KtvuWJ1Yh9YgyKGDRG2qX/5Jt8
VOnPhjni/TBHTK6DJZd2K9Z0fvwUTpaXZtZhhTad++79Nec1tmsSha0VETKzgsmC
oHZwhL6UmhXDNDAl3OJCqzXxxS/D8e2U/PBuJm1PmdVfwHpPXOIlBthyJ+M+SR00
JBCLTxoBweRc5tGhHyJ27l4t+RXlIzJWF+2zp/nX5SB42npecRvc1XcaJum1tt0q
PDdzssEHmXI8w6AybF8fS6v+h9IUr3A+86XbnqdnNDlR8aPuRz9+rD2D9LmxAJd8
cEDvkIy9Pq7V7oWeELf8VDP7Ez62pQQmOMQV7uUFNN1iyfZy7OTB//sfaD20E8Uf
2u80zfe6eanPZ/jI7VhwLNy5m0HDDBe3NQKap9SxigaJwiLP+O/qZtc8IVEQq+EZ
y22pndc0GyHMcv3diTBoR+phjujEfHRDVEaMY/q1qOhBZHNkQUqUWhe1ij72mpbk
Ur6VYKzGP+nhoStipCirOeM8uGj+jZjonkmcrgQQjn8/GtA6ZTK43gnQhqsw/5bM
3H25KDNExLCKO1Pn12+OrI82m1Vm5R31jyQP7tj1ZgyLWnw5iRvizQzVQgWkO+so
zWhb7DhNMurPr/O8MMX3sAJhnIgRy0YZ8SevT5oEBSyySEJV4K9OY63wrTGCHaV4
DnqZI6k2kIxQFeVZgDgnrOMnWd55hqIfKSAz9GzxckhBKUezuZeI7KZOcHb2QNYp
LZsJwssYWGrpD3iuFTU+Za30tCBHCM2wMLULu5lDXdb2q6bSM7W2xJvceXDTNxog
v3dcQDMi1DNgKWpt2QzfGt4e2CtNADJoZFFv+ZxibjzFQavqpWBYTLE44IrxGh+S
HItoBOkUZHAOfvtq8ro2E7+1ypiH3LocClTPi6C8LfXIbv9+PLGAOs8GKNrFZAgW
NBr3MvbnXo73y8BzNjRFWPxGaKfcc7tBCwV88IHTEtcYhjWarQNNmRFgbDw+m1l2
sALd6I2lVMIZ366jyVemFXbyfC9mMAbCJG0JLJiwN9C7yz10vCIX8lqhGBf49az2
rjopq3U1H2dQSf5qXfDMLxvEFvmZUoxQotj03gjWTEUsh1kZs3gZPKx702pFWOfw
ZVhwKzy24apwIxT5bWVKCEfj5zdMKGRFD2QYFznib1DD/B4W8lYLChhvBLrF7lXe
SPTODg0Kf28H2gN/qdQOMgeONjj/Rw7/9gG5ISiKT8By0zA89DmimbA25pIgsaeI
HD9HBoL+b1tztq9wLi81d1aHQpJynruUK+/vWtgZN1Zf0k25ycZarhnuYe0zg00U
nHQDjumiRritMsjvHAww4po9l54XtZtyqDt0stjDu6VlGwM18bYIg9oCphGP5Tj/
NAQbf/VIV4aoNNRRA/Gtlt5WhH+NX4Ep355kQ3U+91MXMaPuzba4TkaGU7Xn9FFP
xQMrsUsI1LIDdzXP4JjbukKgvyoIl2J6UgRZ9CnweyzDeItmKRDuczeOJA4bwPar
rgHuNPeay2ksUlGnDd3GKC8CGCrMxzxqbCfnBCkBEU9MfaxJTrf8JQ51cUrxDKxa
E2Gct5UreRzDbOZ47MTPhDWTM2UwBsDUk9Wn6EvCqIN/7I21ChLjNberuYlfwPbA
Juer61Nve3ddg2mNjsQeMqefo/CWJLj7MIHCsuqWgKr5YeoxhRt81W9eRINJGAXX
qXkcMOHlgg7KsFKOswtS4Q114pggMNJhaHXBNVGDAF5B3/C083zrenVH6CLLdvd3
6FMb/2x2iN8eD26zr8sBiS9gCQSQudiSA2wMj19q+1/ZMCkETJ181lqvb+/jChz0
cAcXg7hOTxlBC/HHubVXObK59kBhtetd+MUK7BOJj2jRGWUvRPoc35HEasMxZTXL
hnSezajHomUdc5v1HxV6mgXDDP3GyNd83C0Bd+w6rTfvpNZSkaSjZa+aLlyB+FZL
Fe/uVcHRswExyAgzzsUW3ASCq9V2g7sDoqKn3/lpyY5Zo1OciwOTCn6IJm6aG6l5
1ZsAHezDIEBCGECZebzD8S7VoiHsZx2CPoObjAGyAOuJccgxG7MawqgFDbzsPFyI
xhhBMHtggolKDVSD8aHGcw+dtx6E1KB2j9Kb+JPmWPX+bQD8sfIuPgRLSI1A4o3t
CPf+ckR8bnSd2ICph4sBymeXoAsUtO1dBaenRDFlKSMkc1yOKdK1+W3jbLyvVj0c
8/UIppekDkDHx60rjQiSb9R2gJJdJzB+xJHMEJyD4xYMYX6nK88FWEgH9r0fFVzZ
vP+/dfcjZ8T9h+n6pCaXR2BJe4mNZlgbSJ/Y4cte07a8+5F8pmwPpVVfkHASoJzA
urxfNS8A2P4fJTi6hbe7PAqPHquFDBknGkX1yw6HMe/E8AIrYZJVfZ7JhjY+Wf3T
h464n0ONFvtKwGQVUw1MDB68HP7agcj7VDUV7EkmqeqP7bL1hzMmHkhRWqGWvRvB
nwDsWCOVXrytpbhhNM8ojXpRFzh1eDH9NtadFzzdJ6nwUAAiHJg17272jA7yHb9x
ZkoWaq4VdiC6M0Q1d4jXR3MbV29uKN1GGlDMeipGWL+/QRxW3DfZEWZEFZOl/icV
TNm7Fpquqay0YnXwB0hu1L34AiX0RtrYPLMNPo3mB7fmBBsle6Kstzs1cXHE7vQN
5ygyaWB52RQ5p4SuJU0m12Qj2h+Z4I1zbo+CnhGdUFaEAfQ67UMhygcdG99p42V5
k/0LG1uNJ8IyPchJLB/GsF+8W9srwyOQjdafIN31mtoZ4Mtm3Uu6d7gE6G0k5xJG
knyygOOvgEO+OyYKn9RiM9U6TcgTTvSDuZdl/ZRA1MjSR6lVW9HPHdUiJZsQcROI
hB3Upt7SC1zRDqQ3JkKWbkHJbsW9QnCxrM24H7PA1xlJd+qC8HfHYom4SPVZMNjC
WnLasgRkeldv4oqVOaXrzgB8sc1kFci4eNCuJtIVyuAKMEUIk4pzE+HkvMgze5dG
LL0hB1SDQuM60S/YOLu+IqqSNJ+ZrBwfYvPZf00Z54Hxf4mAXG+20fQujmgSJNER
BOo6+66W+TqPi3nWtf9TNVmRgN5I29h//Ti7618d8sCCj6CvutyHsGP9blZrDyTF
d9B76ssXH+ZczWHQcjdziDlwYPChHgiLNUBR35UNo0nXvkmcG4gWsvkxlbwo/N2q
1GkP+TH4l7YY/06vWj4FF1ve+/+T7aGCWVpKPdr10dKZKYs5LYAAktChbW8EcLaK
Yla7uo892OOrheW9dODH081vJEAd5ywDem4cZqbtcMZ3O4jh+HFLeMSkeZdLsf3U
3Bqra56z7nIoD9O4gJRs7wj35y79qr9a2lZfxagYCGWdnLBgZsD4Vf3Z4Lm/cDFO
DCeCCfxg1yVOsh4m84W595WhXM+A1Nickbf1U7naE1fW2wwxgamEBrz1mSrUwdnq
d+KcekUpxSMQXof9C739qRcF0AZjSoQixKZtnlmpC5C8vTr9t/tJEYwTNc0IWhNY
V9SfUJh7kizJdTaU2buyZ58IhjFYeoHkoqTQ+o6FWVjcDvqT9ptGdvvm0jnsIdbA
vLsdLLaCUdYk5y80NFBxz+cS0fLWd2P8B09Z+ZAfu4rzz38m5BifARReLDuZNqow
Q7me6/D4G8qrayugpWt/z7FewhHcoIwwU1t1D0QWltDL14UfuD/sRkfhxNx7sLA3
GL7Ghuo0iL1KcWPJ3iNiBIHkSKIxzZAIx+wTjcCRVdx+D2jmLLbFeAscJT2pUhJ9
LsbsdMQYMPF75mnxbe8+Kk1Tm+Y2NDNFQ1NmpmNFg58jUT8HJiG3suw/cXrtvBq7
E7TVKIp86cxTmzH3C+bvZ+1TJw0ymGh1AFcFfmnziKrnnVbmdLV5ez/eO7CDNE4o
HAJbDq1BfXhuz5JV4BgJx2Aarbp+F+gIpSTIcbjptLy1qp/xmSJ7x4GAKuw9yHtK
7zDYr4w1GMGDqoUQEi0YTuZhQpakLLBrbfgFay4HQd0p8qh/S7xg+1jSAqmTHBkJ
GksknYKQ8jneL7hT9mhaaqlxSeO7f2DGJM+mfa7vBjeDF14BL43P+Dj+ydo+mV98
n7JWvIXYygdESY5uWWlUWLodJTkWXRXCPz7PGszyfjuQ9mA4aRmt/IdIBmIKe9mi
G7+Ah9TuS0NwqHpZXx8xjOYaCXKXgE2Ol81oH1Sy5dSahrLAN4NWZILASpWQQa6D
eivcKI4aKD/q8Dqiqqkmkh9Xv/e61WedowJuTxq7acmCyibnx7qNtPLd6IdXDSFc
Zaolj0WEys4UPPr4ZodX/WezS3csj8Fd1X0u2vPl+xEHhiurkRdox5ztVecCNl+g
odZZhhpShWqXVKy2iPFOIV+ab24hlRKvaa6QvUxulMO7PbxleKsE0kCfq3dZ67oB
s08ILeqQy5o6YL4hAKKb0Co6Feid57h1EFvxoCgjbYnYtC5hQkmUjeRDll5lVuGi
dQpQ6hrkowK8InVK4d3aWeA+OMkIcg9qXQkg+jHTBX2clbzb2xG3Wx2zlamIXTBS
arKOEwUjggC/vIu042iBCgzyrI1cwRGuIvd3+/i3K0o35h0ThUP+cDcN+/gxqDaK
8UVrqBFMDnGRLhQ/04bpoBS03l6ZBJLK9CZGfqKS/cg0t2lZUZkJ0Qm2QBKmPwFy
ee2VQ4hr0xVB2Sq4/lAsh54QZZNQPq+f+9IX9qEOgycNZvzqHdUGNhcaQ+rch3yV
EYGGQeDJsKFEok0k6JzgYjttodvcESrnFf+e1CGDkw/GnO++obVeW6thGgHqILaD
AHreV1Po8sFl/djWXxaBBs6Jsl6/9VvINP7tKEuJhxWhnUF0IPKzg4ObuZrigKUT
qUcLkZoFe/0yYIKblFxmVxy0XV4NpWV3NadUL5bOTqvC63B84ZEaUiZCSWT6ZadE
pFZW/2DUHy5lOonD9MkAAH1aoJdbFmk8FtRfFQfttBt2a36qjGkSOs0sDuwl0iLq
Dt3Y8aCkfe0PieoCOhmYsHpkpl/nWX/grOTejSWLWA+wrpbZYQkd2WKEJrNQPM0e
TmEFWOqndKG7NTwQyD6USh8qNG8ZoBxOzUWbwkZJ8PfoN3DEVRLgL6II7MdiF2qL
WfBbmGzS85iFBJ6br/dqN60SzfgC/lAjLBMRQBd15WGIj21Olbe48DMXY2Du9J4O
BPMuOetO+ZImhJKULcphBrUNo7Fe/LuWZExKxCoigxrmGAj0xjYytQOxaUhUT7u2
/KI2wPuKf6H7eAVf4GMnuaqzexWwFpCyzxTOUm580OsW3F/8F4T7k8sp/FryZpAR
U8VSS3Fa2ZY0ZGfFJzSVIP63s5WwOw4ECvg1S6rZCgk6Nej96rmOqF+f/3M1gLEV
lwWKmESuFyaq2LrcJsDgUXxUTSllMmsmwiz7URuOYcEGMBbmP6iwoHH65rd9GlpZ
S24V41Bp5QeYahrzjAe4HuufI1QJHNwTVQwm1gMMZalpalhH66Yf+VNXztyUphd9
FMD20TeicsRjZGV6oqMsx0jD21qj8cNTmc6sIU6JxkOdJTmfvBS9THOZ7oqlpYN4
VTsAXVK+QEVt67TOstMOyaxYDz7HajAXevoBB9RgOJqXoN886X5q86R9GX2bC7iG
22+CIzyY2xC9mysmutzyCzg2c/OHU2c3P0Th4cYP4ALQawRgZr9yBbrPc8INDYi8
IBWK0nAyINvXxbiMVUWWaENrGh7OI/BkL1y/LrNsKgYaLqgtQzSsGGv8UyB1YzqD
MhBKt4tBLFuecTpa+fuA+YZab+JI05uCUrkRZdjU5EvXqxcof2Y+C3wyzS3suHkz
taJv+OmJ201avuZDN1wvwCCdqgHAuE3BJTsWwgSMOtutEwuozVVmGgKVe86WjF9j
raVc6SDLeLaA2vKGFaV9Vh/T+bP4Aty40IRWKfU6ZPCo0hT3tzfMfN/si8iFWadJ
zXA303Z8p5fZxTRWkM9KGPYp6W2WJDaSrDEHdtbtSBIyZsA626xvHobzVC+cPDSt
kw6EMXIR5sfAnzkrF6Tn53csE0z45avsPkVcDPpm0Pi0KWTZx5nk8XhUTpXmcqVM
/zOTy6lUtfDa6lGPBryFq58vqR4juhkvqS6+JnyKuAXfKr0J6bNAb5FDgWkGCQ3T
kbY3/flATb+igRSJdZMJnFXnTIOVlCyBBWOmTO8j8quDXzEZScFwJebkI6d/LBVt
4C/wMD78TS6fjLG6lXmW28Ri00Q4LJuLCzgjSSaaRwFC81TZRrLDwixhb+cRud7+
iw1wul+u7DePOeNxABqFTsL1vMKAVSCnGDYiGlC1Fs//Q5tMrecwBMaOAbw6JQ3w
Jc1JZvQbq/KNR9V6Kkf5zhaOt2m6N4Yn5FWHalYY1MB4+EPL6tLW5n3GQ3JEozef
c/wDOvn1PpkN0ekzXBqP7n0yqv8NUrLOQ6J8rxL21ogmhumqif4h515FSKH+ssb2
ftLhQ1Rcjw8VFQtkh2t96/pgfcOrwfHmlZO8Vsz/I5Gyso9AHZVy+C3ST4Um6CIG
ILxb6vzJUBp2aYhS4HUXfzn+H5yO/6Qtl/+v37DPOJbxiJEDhU+DCybN42lGIHZl
sEvvZdrNlrq8dR2hDjPzoHszT1PCfTyoNlDq5ZMHpT1VL7GXTMCHnzIbJ82pzqPU
Rv5pdQeOiKJ+AYr2is3q3z8ngFluTTd3w4VNjSU128fDlIyS8WGzZd7YoQVRHAq6
+x58n2GrN3pk/ah+HJplF1BuethIt5H37Y01xidQpl0Z6BEdZwHTKeAJpcTKriCb
AR3La8WoBsLDwL7zNZ2D3wLk9uAp+5BnV1l3jz6gbfAq/ocEmrzs0IblNJFHLaCp
Z7BOoS1i5Rb/UKaPXcml34I/2FAtzWwcAmdKUQkJOgh+RR+MEckGAStHwOeKWjO4
xWq3rBzu4xty6XIn9go3f76rbi+/KJ6YSJJf0rXC5zos+VyI1Wyb4DKsb5pVIB3j
whJ1PGkm81FBW1ju6k2cd3wDd/z7awimKp+O606cXJnWulTl22nd0Nu9f02Z2mh5
CDNVSdGGlV6CarBdeh7OsVVdEB+qzGUvVprSI1zRalCf5k23OA19cJQWuh898ulh
ilb+oqAA4Ckp+RcJCHYXeyVPp4dNiHrY2eZLV7w6u6LOV9SNyX/bnkFA2V9eSnLk
urQU18EemN89LMKhmmxLN8+Rik7ZKvHRHeDfnUJ7pbE/dDB1yUD3R1CaxJOJgNRE
K4qAXMa/IBojyXtmvwrdeIbqBroj3oydlaUlL0YhWZLr75TpRRuMjWBIpPyhgfnN
F6Lcd6ffviYMTTCiIclg5q3GaakpRU3c50OJWYp6uxfnk+WZ4vubRYoSG6DDbjR5
UtXdyUqAwvTxdiYLGUo23FCsBCaE/fZzl1DAJ3YpWv3or+jMAJGbS03aWAt1V2fK
68JdIg/rwnEk1Sk0yq09eSgVPKOCmUwCPTJHa97HvFM7S+M2+Yz9Nmw3mlDfz84u
6Q8+85ZkX+xuYgeZj/d2ZbsGaYBAaSI1umkty9MIdVef4ZiymXBX4qV3zK0DOpZx
a+CU7k8drtr18L+RXMYboO1JarpCf36xWlJaupHzg7kx7jdbOZr5UFCdHyI9nxuI
1dQAXMX2WdE2q08OfGQXbDZ4XtQnCpdH8IfMXFoNcgZ11NaFOGF4yxbzZiHzCSA3
XHVXE4NwsBdE+hnWl6mUhNrVjSzkTnVUW6/GjtmYIf3ZC9Vf7glglctJEgauEIsr
tO06LErFSa1E7M03WxUUlZaL3yM5DuWCYTGvWp2hZUTCfZaEpprGMD800VpPDmMf
/JN3HLW0UvAQclGsJ9HpPOMpK0tjrAmWC2YWHRt6rf9jAzbpHu7HNq5FCFGwZshU
D97LK0Buvpkbz4J6gAgKhl9yPeGFP+ibpqPt3RSeKm6iyGn+ygBYAF1K82PHYLTC
rodpFxpY8aF1OJRPepIVh6FXttDw9KF/wIVJ3eeWFFiMZTfVyQzyyHn5bOKpVdAa
WktWbXShs64Ial/6TfI2Cz7RWd293Bmq3/upbT10Ua8J+bCfjtFGL+3DCo6tLxux
l8jnIFv/b3IGBosvL+2FlWLZzAfZw8CMhh2XD/WKcVEbDadUMzBu1yJ3v/wiYsBL
m1QOkmdJDOgJWDL32W6abB1Pa8VdEY+oTjERR0lplbwfCr48TqpxX0lWTNN3Ffl2
QR9E/4L1/j5ugZuZz7/z1NLayD3xyZFBeGrDO9mgRrY8OVGd8Fq/0zYFk6Im3zei
4t8T0WqDT0wCqZvoVaaktiMXUJPReNIm5B7/hAV/tuzZ+7iYpkmxk6f8JLP1j1qs
+8UaLsD1rMO1cDDM8OB0yC+EtZvD0BtWzxbK4RCzo1M7tUTLDvzkKT3fRLbPfMEs
9IQIRhzCAneAKo4OfJMQ91pEPTkKgDS79c+oikrmjxVEjq6R0btBwoZsbbHqMGxQ
cmKmQUSjFRS7hJ2cE9Z4+wnHVSZXAMNbpASMeZRSNyaaUUtCSQMcgDcvFQl7dX7j
PT59rGFBTBWnPq9iHGAJQ/a7bg9RY/LIswnJJsXJmL2uTuj4hYQ8QUuNE0yAf9l6
Zy6qvr1iPnImXIQROITqvaHZD6V49qNLKH0UlCQGf3W+S0fvoBPYQ38WsIlNrN1L
4dpfiH9NYOOpcSMUXsUzw6BTNibkUWH++7y1gnSrfYDHNvdan24ajNTKRxf0W4SN
Ltu2IwSlrAMLtiEmrBT5I4+I12NndigrwB56uN96g8ByiXE8k0QCAmkbOzSTc82T
XQb2qW3kiXkLQWa8NZB0hlJptuA0S3ir+RYjrY6S71xWORvvmkDD9D5Om7hdGs08
BUbjkNGl5f3HWPT60fMh/opuWV2jL0apYfZ1sRD9UwvWtczoGoLXsZGgjU00e7KJ
rHKSZwRjDly1Bd3y6Bw1MdBgjbIIEjsXO3AToNnXmOzgopZtEX8tLQKqIL6KqqF4
mbpD4PB8t02N2+OhDLIV+uJVveHJfFPOFZKJjKMJiHcgHTdY/KiKD1Uw7cXWJ7nT
dZIcNiRBEwcrpoAbafQm6PRKyuI76CcWLnP0jURpNB2bDv70eVpevuNQiQ7sv9q7
RQksoYRX690nVNP5X5PcXJePGA1gVoDjtsxHcbS/P4vgd3PufLMHBOn1N7a403CF
ehH2curb5RSSbT9y2T9UEwQKlFIhywaARBsChPGfnxyFJuSxt3KoMhgKn/wo3gTa
VQj7XdW8P0gmlCDKVf5LI2xl2QesIglAhLbc0nO1HUs0AHG8Sx9P2t1yIIePcTlU
clO2N4EBfjk2u+EJI3Mc6KOr6XTZLbHr7ET+D+O2Ya8yvzFZ1LDFLOCp3glpehTQ
/P7xU/Z51tyHnncFBkPLAaSoVKKa0TLlN2hldWJDC/FEmDUUqFqhzp1XfbMnz1rv
HUrZTdDjYmsigE9PQAvotwNofpGA5JAvZrbNIYVlaW23LliVXVQXlSgEleV2Qjvr
8wq5v9kPUuwnrwhXAUc+7VMNdIwfm5HVyp+wDD4os6C2HLnldyN440KI5P5NTBy0
JvIjxujJWD3+/R90tyMV87zoFyKZqgO51zTxexOsoST5PQwsvvJyPsQ93Km+7FYW
C3GjHPaqMZgD55kY6FTbHWrSZWCV3N4WJjksmWvUIlVh9iEc6KPFw2D9dax4KQzX
S2w5ngXIKE+EgUT2JZoxIKjVfn40BU+wvgjIfbrQ8kpg+nxWeog7dqDY3XFesFQq
SvgwB7cD7XsJYwl1U/X3BiASoLAKT9Vpr4v3/XSm1bNjS9FQOyztP1JqIEzsZ8Y6
8mnMQuikCci/nvGg6zOhyqsdYnxZ2C13gKXwSe2/wxyKax3D7FWk0b+BcwMqI9Bs
biCSg4YGjN3xZkQwnCFcasn2x45pGrXCci5lPx4483gkJdrXJF3ZQ5cmIOuSspnB
guaYme5ydqPhU10g1HyOVqkhwOB5k1gexW+RBE2Gd+URPMKkkM40CgHcRbqZ0lQa
OK8jYcG3/e9sNtYPhTIabSQx2CC1CMk6hKmCwyKDBxKr6ST1Rso01RQj/MJOaLUc
rwtrq5BneuqjEW/hGhQZepEPC1NuYPhGBkt0ywLYJaEhRI20GWVQPl+ft4AmnJ8+
CkkjUJRW2zDcYChu4Ie+VQYsyUjjCAMCor2t5bz9+9/yVrsdNSzAIlPQZheZq5A8
0TZc+dYPtaSCpUOfbiNNeq4HOIpL0JXiVw1iV50fLPr7emikyey4YJfuDUS9P5D0
0UXmCaZ+TYjJEwFr8FXsqpT9BOochFfFud02XmlshyBiEV2CS+1bVrCMnCJGWb6t
gc0N7Yw2doS3AV3PsONgcVC8AJMdbmM+LW9+5llSTiBAs0iFBnUqTlPeDYiN235F
NSJ8WYDZP67Uq/ktz4vXdlZMjHGkhcPlETxUeIJm5te/fLMjb3FGgK95eANHeInf
2KuJR/oT9U/ncnIOS53EoNBeyQId+NShFSvbezOosZTN/G3DoSVBrQKoQd/79PTf
IVP/CeHkulTNmFqUO1k0uzgqMOE6POBlDA5v7yQHjVfQKKMkw5UzVEWK6+HPlPry
ek1Dq2GeeJSNKssAOpDRkmcYlJ5lVAaajf+WLAb8rGhXFd9/g8H3xs7eYIezIsPZ
xJCvT4giw2oiOmA0rGtfgRud38bdRBkDaULsTVOK/InKJVyGvrfbCbeacvlooA+6
pJ/zsgxEJY7Gb+HqLPt8DKIm3C45y7CEHRBF00+MEocPhp0xhtXeG70p0+EiMjt4
FpGc000Ps3mNcKevF+voEBOBmPejU5Bzf14TM/asTMTZ4yJztbbSxsfc7fS56Cjj
M2YSiSv0L1txOwojeaGQ6G+KHIPir9EdPiYo3ng1OdnlPzKrzWrNFgruYrRHdqKA
gRrZS8ESj8TJ/AvwtXDTKCfwrPxQypp9g0BYlUmi/E3eGZYODTU8lPU1mUVxuNUD
RSqnXQEmyNw/vTFRDEioJrX8iKfH8L4kcOa5jB4iLynYeSIG+btO0DSlEwiYhim2
D8eVZMg1VCASVtf6AUKOayPlngZ6HwHrKU4JGayXUyu52IyI8OBACzZzj9jgiUPg
iGson9z18Ab9O9lJBLREYIKhXuVNsoiL8RgykRLAEQMSvGPp57xknL6Nslypd9jA
DRESIYS8XYt797ndEvqLUNhheCWN7AfsOG69QSejC3btRv3ejJ787q+BUolSWwVO
Mf2xs/K/fp5ZNYMGe28Ajexi8bQSRAWC9sq5Q2h+7/UJc6wT2syCheGHLTuuJkq4
MevloM6P/5T4XyJ1yH5WufBuXxOfsQLO2EdcoFsjNUZKSkZHC+7zsoSvyEz6Qu/J
n2j2ZVW4NLi9tpP1E4Cn89tg+r+HGoibaLLoK4WmB1K1HHGkxOFuAI9mfU2jJLTe
2nj6yF8yms4MFsKzRhYUOZ8Gt6towjI/ze3WQLGqmOiHrsFWUGo8s1d5LE5XN1DW
wtgQjy5O2OHay87Kn8D7pkluj/rcYdoHyR+85Zyq7xMC/Fo8hhJpyhbNZOsc0Yfa
HUto1RzkXl6y8SMP8Jsdx847L7tw7HoD6FoOenICzTYfZAc+r/tbO4Qjvu6llLKt
qZ/27dv6lAL/oH2287IYL7xOVMtPckL6x21KJIyMvRE1o2O43ymuAw0ruLPk5SxV
vsa0GLC12gbIYba4n1fIuUrFEfVAtIWS++ETdoi7BzRtIEeNAK6dCOl/2fZQ3I4M
3yUJO5p5s0/p9oNbHgag/8bpsRzMOach0bXKp1pVrJk6BRZIzbNX3LeVjdvdrL6t
UUehSp4p0SOf/DZ5mVIRc2oHYynq3tQvlCIw5w1xOwBqsBXyippBZ0Av5lfRpRLC
lju7670gRSuU8a1Xi50SFUCvsmKa/ZyUKiaJMNg2Nc/ybVP8ER0Rt9izNTi1HIp6
WH8Y0AebVcIkflvQHLXSGsiaaZH7YDAhh0oBZEEUqwOKg+QHZEv62bJhAy7NhRjR
U0y7QsZnq+nWxwQ8HYjS745bVeyJYVCZ5DO8NyP1MeeZKWVi5UmpTjON47O+19f1
7GwgXaGEa7kyytf2Cz8SfwCE51fwaI/Ln6RtDf3o0Xkvbr8ywNeYxeZ9sD9Q+xG7
gdtCuJAxNL7h9ZbBoXTCTcLxs8wkqNUSvAcJN/4+Zy+Fvel42W8fnadzXI0pinOY
vtb4L1vEo0J3sM7C9gH5lMwaJgRNcZtXPVeQoAf/uOCQGEqQfAh8FG6PyKCRX+tW
QCYblj7H217UGnJoIYUqTFsJdej5mBG7vnfwWKM7kUWI4owjD1TqRS1lnPXTGWEn
dlZOytvLyTamPUTekT/fKSSPn+9aLHgjJeJdlw1aU3oVhZjcIViM/qCIsDOPCPS1
iX4MIyuu65TFIlGKgPyCwF250MNFMOjLhNowT+xztlxnpFXpAWjTUWIPJFaWfjue
smHaDGKi/VlXx5JZZ0j5Ui2mQpAnOTZ5VN94DCB5CYdbaGG2wtEauRO5sUUtq6jf
VpQdqHSaZCBcllRVgCNBBzx1isC+kNzuu6nh4roFctPvQsHYpC5iVuV5Fy9TpIQ3
gcXiHIpoCt/0Du5LxO71NEF9bVPVnPt4q0tYbc0J2so6lHw1REaazENSeMx8XF1m
g8H1eNQuAES3zyB5Yn7Fb5mYbpukKMr8cCSWYNiLufLM/Ai7YXvH5VYlr4WE6rgl
WEfUnovl9N0b+b76aH4PI9Px6SwJ+gWaACGTrYbjHNF4bae2zU1d7S1v90sRlhHi
v7u13kCryQTVKaN41JKMT2+0rI2/qktgW02p4bME/wgvvOCHFIlN5FWbI7hvQ+te
NZABBiqyn1pE3iwulmjovIXemTXeR9vSqIrAuX6lkIVjkPbH0vyXs7ZvHWDONzbS
UKOrQoonS/xOQBpvwTN75JhNNGhNanMrAcW55/vBJmMNtvHzH8L6fwuEiJ7VYhgw
HRbAEKNxKUp+mfvdMIzYdWyM8MCHU6UcSLdH8IRz4BI4EtjuIUW884/o6VsOoUXS
ek4NpvXVwRrysBrjTuTec60+q9teVXQspHb/ulMnVyKU+bMMmrfEGAg8tCQCJM1N
0oJaVluCbtTbsLPtBNTl4uuno8xF5+Tr4wVuGrFyhF1dDQywodNm51drIkixb+Sb
hdcQyURsG1CkfpuIqgouBxRrZ+wt3HuzN9UwIn94XVnU5UWOt5a3qagi8KqWg0oR
Cm9ekg22naQREaO7ZEEpek8IDnavKrqv+OnHlcIIJDtUFeAp+7T4C9AOjqLET/aP
3Vb3X3CxaRGFT7lOBxURvRjqViY4IuXUsgTM48cv+eFEFa/PofGUv7MUrx2FJvZ/
iRHO3W7rwk/RS/X0rNYN6j4qVIlsZGores2oy9tRo0qD4THcITrACvV2sy/uTED0
kf137TkVlnlDB0A80usblM66DwlTZb8prvJDGzthsg/TyRCPepVleGIg+xuBjM+N
hVCHb+etoWTZ6Jhs5DgJqjw/52wkR/SCi3blQ/sPf/rRf+7g8q67AA5Ri/LP0/gR
2NpEctNhs1yZOpj+gC3UQZ+CMG+l740OqEiG1JOWR1K2kW9aXQmce0o7Kd2r0TYf
0IontuzZfFx4H9710KBeQEBtdBxA3dEg5Eke9cswj72rHFmE46J8OYcjFU2zeW6F
K93KYGI9zCkjLLY9RRTJUkeLtDlJxuLSXI0kisqGgosFmfiAckRDscjb+XAJaYmv
m3HysvhdwjrMTrOwtzXDPdN5MB8Z++lyvRFF2zzP7GSjM+kn6nsxgJFI1g+l6xPR
TpL1SjOGCoPmWOc+MF7RUpnH7vTpsuqfj2hyJlWcEp+hcuT0h3bY74ICm1Qf5E2A
Cf7nx8ZVnYPOQxNV1HLPT2RDkFPRbBrxzUCFeBXA+cFIV5AyTrywN3GSuhNwdd7s
Qh7VrEapdTyeC4pohLr+autrVUhgtiYZfg5y1eFzejqU2SqqT8gV3rjV2E9szrVt
wCvSOLCnhnzhx4X+8azoBXX2MHNPgW+H2xZYSPzaFZ4pTIDhhcARJurwgBluxX9+
IA1hPln+c4jXNoqwTSh/bv2olKuWjnH/F/Anv5WRskGX4hJ+aGPo9+IdYurxZU2K
STZ8NPg6AUoFezEPQmZehh3rJxSK8ACyGmN1BelfyUHBj3A+qGAXsG2YadxClFAA
8NKxbIAwwbGY9PZICHwm3ek453KtltD0E6MBMcmgWfN41VVrxX9veDLBM10QThSL
9DbdkYpXk6j01NVl7Azl8VviMp3lpAC2jnubFG2g3lbBSOiRWnBQJ1XjEJLH/CWD
17P5WhbfA78fSC4p/aER7wbKd55ACoKZzg3qsPtf9sv1TVmxUtjyU/q5vxF/+Hsk
0vgwYV1dEZ5kYkOpy5HZVgN+YhUWOhnM/wj+xfN39AKZRPV++FXNlhIdmhOEh37Q
80d3tmD5agQn5yTpRVWON0IHcOObkYRlG6/fz1qwzOSJpMYTlL1o7Lx2UoD+vQu4
aTHhXmVLr185nQC0uGV2bKPZXr9MQOX+0OBZvDjnTIEylLDRul+u5WeUD5sZkIev
Gp0NYKlWtT4cuJOz8bsLyLtreHNNlezPtOwH39CrvIBFUtd/gV85ylt3tUrHMpH1
o5kMkFE6l25hMggAMUFzF4OCqbkM8Z4eLsMBbcxTt5MKR1ySEgRcRSPd56DqF0NE
DCQJc/H6p/71STSn08p5VA5KTUjMm/redmtpuYGANR1YqrZMzy3tPjXPCX+Zu/l4
TB9RrYsVKPFN2F00FhlATbXEXwybPYwv1f0tUQpgEaC9R8gX21kB4ABfSjr3hS3a
5i7FFIt/yv0ht+fPd+MVj6Qhzing0BnMt8Am7xZgERxaAl4PYcgGMKOxxDGjGqG/
cHsrCKYMQFhPT0rmHFvONFDB56nIIDehmtxiymaX5i2elan7z/8Fon6wIWpMbNht
IZUJZIL6OQfbJbIUZppKvwKN0xvgR7sTWVhKYecdn+pRdaD/ZrITaJkD5e/0udpg
apm4fBmj7Ld/3ybWinYssyxTnANg8YiosAOnp3PemhrXv3bn2qLbazhUvwyDM2QO
HdRipNpW/DjBxtD2oAuJj4mqPP6WlndPendvR4GarMCBh4SMqV+XoEHIUB4g0se9
IcDoG7Byubb+ErPxxpwtaEeJZ3ssox+Svyjt9vkOfylLiI9Dc2uHFdTLU0o3BjZg
CL2RHoFDXA3+wo3hDdZe+mG84bDh1bJvdGVumhN1SuAPSwMA2j7KF4h9R1onP4Uv
yl39oEAhdEDxoYWMxj0GxzZfnpD5MQj918HEuYoJJ/wW1HZyQx4YroUcN8p3xiPn
ul4dDApNl2bXKGrOXSyNeffNQ64bkFSYefchuGQ4vhLkMIMSGd5KsUPMTffe8sJW
CyK2IvWpkWrh7ozZETk1DBBn5U2b+qFw3l4CG+i2VYunYXxcanXYJuGOFGCmbvZK
ZNZcGOnvKgDheGcTQ2GmkbPohnl0bOxU+lIEjPLN2a4u5U+yW058d+A0IqeS86+J
5o0NsXmNbvDO/Xi4RzEaS6W11TQKcm2ovlxqSKN1BPJKGxO5I1ybgptwJzsgyHM7
u06QQIintD7m6ESGBPsKxLSBjzvHc29f6BmyImPfvMWVaqgqQoAz550Yx7PwwDhg
V0Fo7JcXmUMS3S63tg4kQVmmurrk66w2ZLqPvqHy0RfK7INquOVGhFbcxaCN5KBm
DmYZglTRKjkJ1ZPHKaPpdCLLIXLGippLGpB64wbNBCb5qcWS9slXJ2RxYAIv+p1j
b59ZxbpZlyaiB7nqhBVXZk3msdHtNTK2QuXO3wCp9vr99Xp+qeusXaj3teRh/W+h
gRzcH567NORnNJ2t+XDTW4MbCXHe/l9lueI6Iy6CDNc8Auqn5LY6VFPdZuZpDDUp
NO3ENpu8kGS4HJksPwsZ3DYU19qat7u1jxujZVBAoFAxboXS6uTIoPK8LJRFAtlA
yfIySjZnneuKnnYlKu803gKYCBnun+YUfjyP3Aq+4OePA4CJOc9ceyEn+/oCqPpn
jGWatZTu8smdVM4VSC2KgQYhJu1znZhQIZiFWlnb3upaOdgc0VnkVPyzg4tjUXTS
JAgbuWE4VA5qWdWvNpDfFRn3Z6TI2zNuVQYOpy59ibZaQV4SIbUC3YsPdFq9UZ2V
HSqY/2zIvpsVff2NoQta6T753fVXLS7/xQhsOVmCsDxgMXmcqEObQICjGsfqbChM
DJCbFB3nQ5FAIVrOFvZWCG/TdT8O+NroPgxg6sPoKi7+dku0bSrGX5hRXRtTCBae
7hQQ+d5fwzYy0rAynoXymknM4TLjIis2v2xXqAx45mZDG3yswiCQ5tksXZkELLNn
ZhrwJrvGhn4bwbIZ9eKBNd0MI42Tfc+zPRpORJaVDYPLzFhgH4RKuxAK8Mnzaedb
95X8TvPLt8BtPgsmuAxja6ejuvTB7XzMDukc6RMRLG5nd76CODy+cLSPr02LPMpF
O43l/mbP6d3HgKPOcUHtYu+Tsx7iwbo6BrPHegdG4PCE87xUAzydKuDhR27hI3ym
g6lUkCTOY5wFECufx3/A8Cg40QBRAu3501I8IoY1wiJWEAnt+OKX7mjXxiwHksJh
h5aWD2ExLonK96jd9QMTJf2P8PnG+GRTsK/esv1mjhjK2FGmPFr1wrXtMb1x4lmK
uCPVqQ1XhgtGN3kvy5aGbZBEJpDlXIfqAY5vyc6laqNaTGP4ptZUYGFyYL2BQRT3
ymhpPLkVndLNSbFrqA2RnuVffsUTLUs5wuJzCtJZClK4kzTYB43wpLwgGYuWK5bs
okEYkPHpOBOUoHOLREu71oEfzO5ozSCittZ92hTstQE5SMVyf4ziapI+R3fsyJeK
eVeeDbZG7fTSpDbbU6XrZpzYDeqUrf8Bb3ITjHrbJc/2rqUGpzXER/Z1T+EhduwK
rRzvbweKKe599cAPpDfjWPSCo+hJDWvHRfxU3J6JaOR3+LIegMKT15xtfTSmpCen
ZD+dTwc1IA9cr7rEypYY3lVlVi7nFC4l4tWf1WZ5SMQCis9/qxjONeOBAAvXVaaK
U1qEJ0nTQROXw0Xpicg+gyTv8zs63f7hPr6H5eEgwV4qe+/5jMWvhRU3J0HfBZeR
+4XOyK+cAV3HcIyeVbYSOr0HtTb9VUh/KqYXmno1O+8p4cOOhks8g+4WMEsGhBbl
kzo1qUPvng3Jn0tNjD6J8dgg5kN9JeUbfDnqhn8+MCiq4qH7f4JWr5HSGiFTp2q7
PGUO4z8Hql/WF7I6HbCEmNa0oLqyfL4D9968N58OE7+ArjRFjJFqy2w4BtCsoSQk
QYAcmbIpcxvx/BCz8k9V0yW2XLLwBG0jXA0nadmPlGMKxcrH3FZOPR3d22LMoh3z
P7DK+sdbH31nH4z3r2T1qePHkra0rS8xu7ARdCiybg1sW53MMKPg5RbgeSflOn4z
2ege3dhx/QeqvJyvCjbW4LZJDfen+wzQNRrTF20Akqt40cm/Viu2eSfhXB9d6b6V
j9/E//9TzTX7nc/6xAyXS4ozHrVyOk+s4ecspPhFqVsON4oRWgfok/6Ku/N8raoS
BX7dHw2gbKd0weIq4Y6aRBTQVecl9W7/E3l9tSq0qNVOzhjJc7l0v4XM79t9OZjZ
QW9Fad+xvd8WKL1iv3ZhDOBzM4aqEHuTdfnavidxj7Bk5le0y3maboc060t+iOdf
ySHAu6ORJPkOLZOdqqfxBUslICfFZ9lLf9uxE2XBi1G0GQq/d40JM9VI+VGo4+D8
BmFhjpLuMhycSQa9Ezj+LfwTIzESNqxbK7ME9i6dguKtBpDpdc/6SmQwyuX9bsF/
9+IcK39+1dkj/8CUmXGqOv/r4xBauMt5/HuFcYz/Yy2CsMLxLJeU5dBzp6rIoLnj
mOrq6MuqXZIbhuIRprj3szvBQLFo5MyhRMO632mX7VCpLYVvzoR1VW3gVEfJzt+G
x6u0SfUKmO//6+O10G3E+Q36wJ1bYHBRi4smtK/DIolc/s8oQGHnoHIqtVlvMO3b
OKWgmnPT+zzo7ZEwEbdN4BE/y7xbDI+0il7mdmeOglEnnyUxdAJxxZ+DNlbnIjLL
BckTNbvUk+Ao+zTnPbrE31Nfsqq1O6TLEqlMf4g2CNMT8uFtVHnBI7aMgR8w+Zrz
x2ghzKVWzWFBFm0F9C0gkZlH2CtNydgZ03+BpcPu4g8OFrH7rn9syPJm/MbJl+p1
UKdg8Lvspf46maNtT8pL6f6jkXLvNYomttQlqH7P1vQ0Eg236+lyZwMthBuLNB+u
1jCaSb4cVWFriKUBf1m7zWWbSesT5/vh+DqcsSOgVRIExhOG9tBl6uYUyRUVl8ma
lxMt75Xt1m/9M+9xxYGOa+Zz/drfyFvdFr88jcS/Mxybi6dDqRYt7ihfB1REYiBg
lqWmmvdkxrvNJhgaBdTG4wW2uU13hauID+ac983NTfWxHAC/oHX6ViZ9GiuGiTBc
BD4o2bw67jIvsDLtMaOk2T4YsnlEMDxMMzaus3Gn5Bdqiwp47PT3JyQrQS0XPT9f
lAgPXQ1/zA1U40f5gh31Hwogv1pHb2+BHGRj4PKN11sEtmDMtQsNjZDz6N/ytUgu
rzhQ+ug4ss1+GdDGBBTPgqPq5uJy9pDLLv5OX+9tYiL6Tfxx06RFWvh1TfmPYw5F
FD+hxVMxgmKt88IEwMgJzvX+V8CjVaA7UjQxs+2N9FB3pqGGjs14Aln1AF9XLhzP
YoTdkUFX3x/npweLUrXP66VwRKkJ3H6UyMh8X+0N6nvAibvkWMktBhYgAOM53Z0G
kb3a5mMm/tXqqhbt8Uzt+azq7BI3sYxicw8G/MtaPOeXeVpR3cfM6+OJC8WknTiq
VD8N+2aWK3yRb0vDJm3AYeDPtti2d+YodMdDQK/7j0+ZdwsuTFeBuS+oZuJ6xC9B
yu+/yvu/UZMavS6mKlDGxLNhNv0wFJQc84V3qXIRtP5h6dXMIZIsby6GHrZl1IiH
xtCJTMJkvYvuRamUxX75M2C9U0josBBCOWFT0Ty8DcAx6VtQcEeo4Ast8bo/4oM+
fHA0o1kQTMzi1RzfJoo4TMV1MKd9/8XArH1JzWZyA9lojq7cMdu1LTqfqX6G7X/I
d0miu5CcglEq9Lw6146NL+uvKUZ+3av4gFxGXLinJE3jcYWmFMUKFQ6CAm/FbhCy
vGj8eMWgPmVYcQq6hoDqN66Wg/UBOjajQ1YpmcAsfNUetTq12EGTy3+U51CJTU7Q
ZEDHOPzUCHC+KvzpGQKmyiIk9G1bqEjJHlPLES/x//JUgMOlIGdSUpCGTYI7FRCc
AbKDM7l7Gd4aFkLaOOH5LZcMBiaDoq8BXvB1E4zz22kyQjK+flVgvI+mVGaIYhqm
P3g014G0TeGvUlaEE3voFgREweDnZb6X9a8zKeD8diqUWwAWKMMw0op1gW0nMlWi
aBEnKAXkttwM+lKgY7MBgLsjxJt1xce6YReY+ouIfUdqTf5tMPY29PE0bNZ4UjTm
BLRimhL/FNtic8OmJsYsRyzhMIJBq8Jp3Ri1q1njgiRCv+NWi6oh02IPlxLZyjs1
aFsQPENkB72to+FJ+vbCpchmyFJwNucWNoK3hremvePbA/zDPW61/C23heS4pzgK
b/dgISy8TVuO0x5ekF+hxpzwCyZ55J84F51QuUMlwSA7Ax1TwtpcJqbwIyYh2hZ7
3/4jBmiiFXG4HAydIIcKrypsUNtJQL4mwxiEhUj19cABOQR2b+i+rHgAjFD2ZfS5
mmUeDZno+gdPQoKS0ES/16nuzdbiIL7qVbdE+qioVRl/z5NFd1Hbe+RBDfDOBlDT
roUKFDrEYpz/Dg/K0rYLNx4IUzut8LsFgq0Iseu3XfNRnVcZvjOXR4aD3Z+MhtN2
9FMNz0f7wIqq1fZnV72s9lYaTMi7ZpZAXBqQfa/yrSCucoyuhDL4TR40v2mYH4d/
pYPb9xLvrHR6fM0LLX9ijaiXT35SsBsTVu0N+M3TWqvQRcXmnhPdwUxXwystRhK4
aQ6upVVbu7E9KIdjQwXyS7fhz0EZDSn/gjLWlG+IZItSzRg4LOa5g/XoV+K9M36L
l7g9IoWEVOovV9VUZvm2B+H5Ev1I1eTmu/AFTRz5IEKT48HuC/oRueQf8Jw3PClt
SIf5QLnI8eovtkMi9TY9D0nEp8uwJbGAlf3I2EOJklaYeTf3lgoMgGGvcg/vS4T8
g+pQNa4FXY4CjDyej4sgnkqByA/EX2WulFXLuHWuIuZyUu54n8TOFkvFzM5UKH0c
Pap6FISxyvy035uJWF/Dr7h4bm0eWYvIkFUniJqUtDDwg1FYjjkPnqilYw0fHVq1
Kotc495lec8l6uVRzpofKPl31YezVen3QwecL87aHH1c2Fm4dfzBGlg2e3/cx7bN
P5b2rc8rXOv4d6Byu36Tjw/vY0GyDjzILRiGFRFfpp971yjGZIBy/qJeQktmxBHe
Wilk/40DaD4REQBBoPDVGZxZBAzMAt0QSNJt5g2Go6ip+cgkaoEDG5aBRt/53MO/
08td19ET2SAgZziOKLjH3Mh0bbPakQJf45tnZLnu7cASONLJY21j8efkdfF1RwRa
oJJuUWpy6AxIDdrj85cfhOfmsaiDtTs5AjHBXDYiEsVHTDYrJhbY/RFIyFsScJe5
m5S5K4sYukvR6mVb5zh9aSXpaITp8DUhMkocCgkdrw6vq1SbBqHCiYHgVc0Rl1u8
jAbgVxtGxFIh2fd7a24aC42VomPNazWANDKIx/PSuq6PSrKncpcuyuAfnG4joj8d
hnq6qxSopFpupJedIu46qzY9715C9P+f8+ADV70nBqVVoaAQJSMco7tUPk3NDhQB
UTd5YqpSCbPls/uD3v9Ni91dD/tkCUHebBKLuS8fmatwKoJOsiG+9/PLOwAePQQs
KsylDwZawXwVC1xpLBsYjCw90/vAuxblV7uYYXEQczQkBChDvOQs1aPvhMMyZFCp
UEAZg957RGcanpUwxQyZk1D9f800wpEohqtwKFTe9O7Xwz1e8ZCXrTT9nil/JYqp
DNcU52YV3D8AqmRQG7kPakDL24eos01DiS1PpJZ6mYwRcw0aXiAdsTl5KC4wDyfJ
qc2czMCz2OhJwH/VJuVDsj5nJmE/KYgrkuGCiymNIhQLCDCTGSPV6/fsiayP6dCF
WtkkXKzNZGOobUa3bhkNmqdAW4m7k+b8Pm4JgpeHsnkq/NZQHwXaMJpfbpUqgppG
ig19IIRtQHQqyjIebU2vGGv8Y5MVNG3bpxDZEmgyDIciGovQMdxC9OyOtLBUIPbr
Uj7acGynvIs5fr1gJ6H+THF7z89pnyysW5k0QN8MDP8/HDxn4grZve1H8cX3lANg
4BRE1Z6MNCNSB00I5ml6ai/PshU0cSfJ0MYXIe/CwEmfBWPVTMf+sXPa/yOe4L8Z
V9rzY0MHQ/SBpvML1aoEOC2EJ8vGL5UX42rGN5KWn0tHWDEq/uuMqhGfezY0A2XK
xuIA6ahRyqqjkSf6CLzM1BaMTpeBR/hMocdURdZZtl5opa0ScMuJXSaO7ypeWjVt
LT5wcg+7f+x+lwveACp+aZzAsbkajVwPs4YqDhFNylfvDp0m7PDYoDC4em1cA2Pi
2dqovX8Tha6Y2w/APLd5KXvfWlhamI8aqLIewyACaMsf/uh7hOAmNL3B83JT6wII
YB77wGIUGaHOEJrHWiKX4iEkDeIjwpHKx9l9Ne4uAxy5Q3iBDiKaCHZkm5z/UuT7
nMBQof1UoR2T8tPaBS7/QspXSjew9rF1sFJwHlJiiaALwPNWJWisosEc1q3uu9c1
Q8vdemg/f3CGoiKNHzA97nMvHtBihPXTxfGFr1yf2PaZmkpgFpaTUsh5moy90xyh
heOLxGBrG/bWJLWWhWPpop9BweVeRubV9ly/dirfbShG1VC7Bo01Z1sNCsT3JWui
LmiXju3G4j4j/MU7lmUCuCArsVHrwXmKi39TXzYcUMNwHuVpRSewZRkN38Nl+8pT
X4D+66kNJYmSXHpP7aZFq+b5pWK55rzuecDFWuK2OD6Q+XTENCsWT0lx2gi0eKNT
zYUEIZoJCHoZuo5+oX/sZbOYzjxcM5kTn25oLMRbx7vzLLvL1vV5vfnCFvJ46eLP
y2drpnLXbnP/2mZjW/6GJcNgK7CQiU1f3ajctF5B6SVx2tp5kHYUgem3/XWKMX4V
WNm4fV4GDB9FCaLrST5uLe1MP/92X9iQ1r26Kc2FGTqW/+QSa/l8d2QSBR0eUpz0
6vz+mAb5Iovf2mWGAeNbZbYrp34Sy0Lkp6oywVS8VAa/b3hOhpd4bCwchlPPU2P5
x1LCiyHJg4TIpBu5rzNz4awzsrxk4jJCUXrZVrb919Wah/Cg2Dy1RfQU/pwrKFa5
jucjPyCSgGXHMKkKkLp0pbAXmFP1wRRwD+BNlk/hKjGgmKO1PEYE5hLP6DssK4Ld
1wm0Y5L0dtl52FBUKVcP3aJTN4+7GeOyh4Y8o1wdyqLQB3yNcT2bMeUajuw/EtRS
0fFpZpjmaS2atBxa7HNuThjDj6iZaX6/rEsxoaazN9hj5A3aZemgWeaTilQgsLwK
Vox6JY77h1Q0JWc2sE8fJdg+eZWk2hmOii8NZMLK0LybKxetGMxP2OobezU2ijxP
HFzwB6KTcuJmY49aojG2//cMebTOfr4ihLURaUHUD6i50vsapwrFUg26iSUAV04M
X8f2M/+8xBDA6ajQFMYkPxxaIVnNWxe4tdgQoHcDoQJqnpdF7Ituzb9BkkkpS+cU
NboyICj0a+7t6L4Y+ChkgPDf8GWkGsbHTngZTB949Ezuwa6DbjKxnseMHYe2Ppl8
xFFiYoNAGH1DvOYqNBY7/A4HAEm89YvtgGRkLfxCnSLcP2gCDuPLJh6aVp0dIEEI
18ZRawd/xLfe4n5mC1sji13eJlEaFX2qgMW334xKsMKBpJXmgTslgq8SlUChpBLd
K2sh9JThicGZz7FlGgRbFq22djaSqhXeRSRptwKwaEK/IzVisGpy//FebaOYk0Be
MuWLnA0rluB4aqc+6znzaN81pNgzpQJW0BaEqD83boXxGOFPc0LUwImIlaQ6maas
uG61KfU2NTjRMrn+tgLtjpUzWcXJJqDP30//LhHS3i9J/KiVE6eSHlLX+5QuG9L0
bUpawsb+0IXKEk4y9BOHOv1FmTXK3Ave93QGO/2tNtIcS3gmRfPs+6XpUMOybVjy
K2mtAFUDQKKvoeLY5BcHI9Fx+Y5k1zTq9Vb1RLyArNUKu9UI4QFTjsDUFlT54K/4
R+G3+MpRbHawO9EOx9ErWXsz268EkTrh9Qo++BcedQ/OAcfqhvynKpzyCCIVlMTp
jqKiMSJmbCc8px6N8AjkUL6BfKir22EcT3HtHa8zmjNxL2M2d5XWk4Y2flk/NUUv
0QdtDW1X/avrnkPmI/ZHAqJt9BTuFO6Xy8HZM7VfYkNRvD84LF6rJ8zCmFxQm/SB
AA4T/3kVJaZPASKnkeSzmY4rOMWhZNo/MguC6v28y8h+qP3mGoawGLWAfE5M9kU0
tmA07as9TYQbKGB/t/bRT1HIgF//q/8koyyRT6fE2cMzQhKwbbQ5CujGxhESuhas
XGpgesy9Lg53t5z7KCn2Ina6JvwB7Mt0g7C6yw1SueCY3FK78sE6dp/oNNZvsVX3
VuV54/yQ0NgCBQI1wCsurJWv3QqaVp99kMvrPFm92hd1AD+WOENc/DFUKI2LP2xn
THK06kacA9qM4TDeaboHYUmCisw3UXr+O9XpKZqWYvBJRcDEL6ByaV8BE2zPfQ4v
pTpqz36tp0wsPUWFNlIDsQT/UquyRogyqyKtcneRKklG1lifGYbWkpULdIb3APVd
3Y8zV0bUgOaOAiJtbGAI1Pa3HHazarEvXVU3A8DdfbN3PSMKlN1ff1uCsFeLnPox
YN7ydV5i/A3AfUgOD81bjSrjcgqKy2V+JAL3UAVAooM0haEfftwumf/p5bvIrlRE
fuAV+Nmv4dUHoKvImfPQ7UFSc0FAvOA+X6dkvt5TAkJ9Qrr2ENXJJr6MrqB/eDnx
A7tIS6TWCi7fiv+gxHe2FGS7//U/wmgmT5YzG7i/LrkRwnQXmcxbduRxwdNDXQMm
XGTQ56zZUOAYKJ0nKvef/E/qliNtHfUW4NVqtdqWfGtVOKqsRqXsfxuVv1mgW7mW
5n2dEhleIXK90jLCQyZshLva6P9nuNP/M+AS8sm5QBt1INIkj11mO6wCVTEn0o0Z
c0kJZpMKFf0MPZpxd7jyUkosUsDb5DRauPDNesKl953OlKjq5Ixdc61dhh638YQ/
6xUW3Aw5xJ2nC1YT9bQUUqdIRd4PGaArlJOqVZEBXfQ52x6vrU/o0aTKmdd7+W3b
NCwC/LbrBxOnrXd9Gv3HTvpeopb2eauDEJspHZbXjD2YZr+OyDyxexHWbVKAnaK+
EHsxBAWo877jWRjze9AXtwXKXu0UrPQzcVz45bVQQtvZsOBvrD2qogVheKp2mujO
h+hcsM1WhY6AqDXc5kj6uHRXQjbKHjmM8jJkLjBJ2gWPJ+pG2VVg1sDfqk5wxSd1
B6yYV4c867CZNn6Dpo+JB6K8909e8mmxKueEnoYSIZUI1iljZ7J8MsZItRxThP2y
YlgD2HPHzjId5dXnGYyevjJV+2moSfJLmoIbB+gA0QGeC8TPbAncyDAeBcllhSCC
5Vh4uPqRDTqgEpmxfXFQQAezlT3EFoHaxh+5y9fUgMJxTCYBOOCry+LY2gQNYHCK
5BjWTEK9FRl2NpXWjUcGwylF/2HM6ZhXkfEkfOkLkO99ym6Pipik5Zom5S+XpBkF
8P8cLsj2s6Z8XbmZ1bzNgfP9KwygxqqkIiPbu3x+WTxoMT3kq+wpz60GabI6WjOa
24tacLaw4aqFT3ViOzBqyeWP9IYI2PqDhswlZUasrINtAyukIFoKmVDn3LtDxn4w
2q/jqnrYV8pv4jMNkWr7+8asDmoOOne2bRfs5NuUIyH1YszD5CmU5QDH3zZ+iYb9
8ISNgAyJverhPOS7/n/p2AffVEhZQ90lsFfQ7q1JtbmjNtmc5Z4YCOdY1eqbnFfb
In1KUCkm4boQrLcdYKkeQp5smotdlvJbR+253wgCZ9Rsj59Cj4nF0X0W5O/DbwrS
0rXIENxtLuylDG8H0nOvKMIBVr6Az8RBx7DJ6CkklJqHUUgQbwfYNszDu+XDBEpK
Od0pWRmlSwQe23BPxEW/oAJU7W0/Xti0VftYx8+m5FUGtoqmUq0A5WzIs3gz9ZA6
x4muEiCM5jRH6tD5PEDqRhrwSh492aNSoINqxkaFOwq9hwKg0YM1JUgpObb688s8
GE78sqHAwi/6j1jqHZolTh2t5STbLxQ8+42QooKz5M+LF5od2cCLSDyRDeAZauIw
dR1VHNzWPDqP985pTP2sf4ViTy4qyA+XWDjA+GCcBICqa00to2bMwIniw8Qy4wKU
K8k+3RJN1tBYslxzjZ72Op0/hRbzAXKDbc4XbnSIuwvFBVFAUkOJQ+45PRYZRyVC
Ccou6qeHp02LyaIfgbCbBEn71FwiFOvtjhYAf/DbNW59wyNRRoc+ZnfS8SWgHuwb
VMjrG1hY3+flmWcWUnt5djWqLml8hqd12JsuQw0odT0GQov5ObmKxE3RWyqqnWQk
xFqMuxU9svNwCJyB4p4rGoaZPruU/GGP+I1s4p0qPg8mNMR3xvAhPmHzhplquKop
ZcUN53DIGTgY6qJwmGQlazEPqKWYuYJFtH1yFpTYqmK6uySWuSs3+yIQOedSkCvN
8VFtaePDpT8chRmNgUhgm0MBHvBEM4y3wpnIaa8B0s+zpmBkWF3AirtfKwf5DdeC
jVD7+tQjdIgZq8aMxDGGTf7cwSqEtNDcSQ7egoZMWgn4BzM0XF1Cm5qDn4+hC+Pp
MfQaByjNOMzuYd4P5LZeuwG6xaxDZW3qxrwN8GpvTLV6LjJodn8/5ohmC9ADz9f/
53awT36m8rY/t40HwuVJEsze80370KgdSb1Yfb9r+IU7UTmrhWvJa8PS3cVF2a7I
dqEjgPrPxLE9U8srPZKBHIjOeSvgY+DhKex+Wi2EHnWoZY16C5hVjPJfk2/dnPDG
tGvPUo+nu+CpluQnk3TEcju5YeUODNd/kYR1qWF47pNUzuiYdH6KxRWNI94Ffj8W
6wgGUWvLA8V4AdElSoAlRtA59WbOaanNsW0hE5MUC1yIMuC+SMWs3/txW9pIRQJE
macfJZ0gOwch4a6nmbSnRkUKlkLHUlUykdeN5cFb9BpOtwsQTEPvMgu0CfkwTvSV
v8h9dYZP13Sgk0+B2YSqSCRsmZHFzfqGKukF17t/cI9fjXOXjC8MYsSiDIFapRa6
Nd18yu/+KBf5zWhtvDdlshgnsMMUs1UDqGn7fgeHtNt+Hs2g3GmNMTWsclFXhVmc
Fx80W/rCpza3K0UG18/Tt0zS4toNUN+/xBHcEceAi3ZmGCnr+O/fpyygmnMhJQsf
Zt3ifAZ2dj81qofW/SrELXWaUUGQK+7EkeIhVq00fmlBQbZIMxFBmhx9a2sgWFi8
GFr5IP0nL+CAUfTctnEtFru4BkbfEq8Dlfd0U0nMfkiSaqqv/Q5GgxEyprqZBchl
FAKz4DMm8n4fKBvYrEWd0hh4rVLLlu9RwDZ8KZoDBMM96Mj58hXxFJP1egIXsquB
Ur3vjoyUUaUm+I0f4WiFzCp6LevyQvE38+aznx6x13BLvhdIMjv88pLpMCEKDUtN
Of1YKe0Oa88+UCO0Gj+SQnGsPTueHXvi+2BeQnmYzlvNI5WaQdHXh1Mge7qNeP4I
ZSuAJDyeM80cYvVt06M8s5j1O8uYSN0SgC1oeqC+lWi0qQDzOe6wnlfej81hwi02
6Ao44ErDsDeFDeiDFWxoGtB88844rnCUyZSGKRcfW++YqdljafoO6QluitSKuiAs
7hcYsLvepCijVOHNq2vWhvWvH6B0Si8HbADNIFJhXmgb78FxO4ZdE0i7TPnf4TAP
DxdpLh6mQ8rrOQYTnbQUTI9TgcUMY0M5HM7t2i/jbh1ODVDv+QiW+E4EgXNYQR8B
VGuime3gR3WBHWsnAlYdaaPLrH3TNrorhtOEIMR9uqWVI0ziBoSjFSYhxwSApwDm
mxk4kTsVTNAgRJV9WJr8xJP2YJZY0wl0nKjsJTz7O4n+8d5DYLL6ga2hR+Xdr3o9
A6RDmA/U7scXmf/nbJvYlgnX7TTKItxv/AZYTAcxlywYwsvuAkjtTVWqtevliter
1MoHQ0jeUXABfvkR6ozWsKC3WgwY9qMKORMindXmbRBrpw1NP4sErNDhUda9iuDF
8D34WhZX/zEFs7HAcv4Tc8/9GslfeKigZmfib3e/AUPKlmdCoGwaT4cktmf/7HBU
eGYivMWU9p6Jro9G9M7BNVS5+WmHuYQ8mWi4kAntmMIWhsek90jQP3k7gd0Y8BYT
2Kygd7ICkFyL9DQor4sfQBmoX+RLr1ZVY5hb3D5xpbGrYreu9R0g/9kPm/sUC+uk
0ShhYe099eXOl9lGS5hNuBUBKAw4Gdw6RoJW01oNzE+6WGiormklJxAfGIskO6lk
4SvlnDM341x2FjDdSqL8bF+Uo3nvxQnsGTjcRDBP4DSwquNHoXU72D3DqRtUxk5s
+iu1vhtnhMaojDZ4wYPWH291hdnD0TKrQAVNewReB6NrBTlv0fqCikOQge/AWTFz
3KxarwzBr+9mItCcdebgtflSd3L8BfHAHG9KT/7c73u/MXed6q5Vo6IpU9aThfWk
xPGH9EJru6XozeqMshd4BIqOD6p5nx7l1/EcJr9OlhNt6yet8Cd9WbR2hIeyjbpE
aOBrK6Lw2Tf+viMuLZa55eEGHnQiI79vp5ng+W0h16SlTH5ZdQUGhOkitLvv1fpP
JCEkj5+wPqlPU2I5SqXjRcKaFXwwRGxBq2b+jYD1K4BCK87rmPpliXB4qFuCVZSi
KyJnZcJthBY5Zh2mCYHCRplBTNFpYcWbmot5yWz1a3M00XSLiM8ooHsdofMR3cRu
g843cm5NH/I+uT+c1GUTTcz6i4CR5hQu0Derfae2GFryDxvIQPnLL9/GPJZu8fpR
ohL3pgEUEKrRavqcogIN9i6VB1ubuykNZnuKlObYF3Sq6egYvna2ak4LcXYkmiYH
1Yg0FckyXUnM1aMPTJbsMM4KFdynW9G7dE3pdkwxNW5/mM/a5xKhgQhCNWYlbg/F
ZGuGqRNuONS/SUW5iNIyvHmROYMNLaQbZc3cobGuxDY3vMiepQSbT2V5PzbYP8/d
nmKZQyLr2967dL911/Xj3iVDHlgUdePi1IZnnnH+6c0GBOKzgAmXNkUcTr3C2e2v
83o3WakxYo3QFqKAR71FSBSnDs24RvYq8bdvWQzsUZt+cdiw/OJgh80DlNeIgBRs
ZdrIPb9YEl00YUCecEWDJFOiG472y0Wqr1i7FGSQ9dTPx+di0W3V0NWccVQv3lxP
LXuInp1OdL4ln3/gvaSZlLtYoK/9pnLxbBNi8q5iEVU1PV8Zi5efskZbzW7sjCl2
i9QPek706VR7oMAVOqiG9RUx29ZhxMua+DDsRANyLGY9uS0222GWXI8P5hRZyYXI
TEnJ9ziX/0GtAAMaaRajvD+XZzDNubvL4s6nYzpiz5jX8yeq5TQLEY6Aik5Mt3e6
ZUatodfrDg8QAhwsCJThQZxt1ZTJEFR4dAsSB7Urwm3r4nncqQfJGGo0NmOAkCJV
vensGYCHienBiWzFJj8h7vA2olR1rTFWlsOl74M9dLTR9HY+zeN+nXieypBg9siv
B4GEuuVE92ipe3uuDc9kwLP4w06oEIew/CgCtGcIkRZTyvx9LqET5wIy0rQpsRqL
L4hwuWsxvzyen6KJcuD9SHR4VwrG4egohB+DC7/HnwUSWk3N1m/7FZnkDvgxQdb2
98ZD2HQZ3CkG8K8Wl2RRZJOCBRMIlxD8gdcjpZBWgO+WFD3y1nGYylDNPTiZykhC
Zg7ssTTdRgmMk3nPAsOsSNAuQ9YKgKp8aVDS8uuzCkeTZAk7i47K8N74qV7zV6O5
3PeBC346CaTezF0ZjNZSZso0/6oMpKSUU2tFdWt4TOhxL/iLnHmOrAgRo5g3MGgD
HfxG6lR8ej2VNBdBsVlbEuU0pY1V2W5TD+zxAlHRE0axB0U2yU+UoPigxZlaFA7f
exXRyS0ETnxWMOf3aQ63WIwLcUUnhyy8KVRMU2l+0cYxljk8gXbeKyG4YZnfqLKT
Js+4Pwj9cYTKOVp59j7Df82Kszmnau/WHJ855tbMq6EFj0j9Fy1nUDEGznsufNN5
84a81pbqAKPEMaE0869VdZCEF1EToIZDCP4XcRf7vnD8cOp5lkMwAMQp6bqvfwdJ
3kGPEpbz4ZEVSP4RPyTPJoSbcYX1sSenVO+7heF19KiezXtWRi9K6xV1jlxiKIFF
uzs07Ubk3Yo8HTUj9QTgvQhGci7N0ADqXS9ZQvu67h2RgYXuZD5u8oEcYIM5wUu/
Ly+C8JJ2P6vq43xIKi9h+R8dMQAvXTsLwPT6t/rcwy/7b3TTzZ0C2cOa3v6uMfyJ
8xCNf6XTSffYMe2/cCfk6OUqquGG0t9MXgv0+TS6mBOQC/ikqZgATbLP7T/6/Vs3
gN5f/geJVzxo13ra/htbgerhvEmRfn2b14QAgP3hzIxBcoJQCiymVw9LycwhCMZY
n+kVCEUrL0jSltsfZAzAG+1JUDd4vAfESdGlqE0+glaKiMUWKgskfux7Dunx+iKu
39fu+U13A+AbkBx8l6X+ZrRBxvjwdKmMJFrRakz0noCtnRgfe7Aqs6tgOd0bf9i0
88bqbPu9MvpvVHwaeVw5OP1F2KqGU14MHjUP+l8W6wxjwd4BhkluH4btWoP2wYNW
I6BRAYFmflTmvAY9NNO9bwtffXS8hPiQ+1XqgV2m4LBlLu/MqBimrpOF3Q8os0E6
gIYaMhgPoX5GZg5p4ObzRS6Egk73T7IuRhOWkciE2meK7XkBGpkHm3JUUOG+GxT9
+HqpKoNdPHFMW/BcO793ZYfhI5s+aRwtjPnZ1jA1oOdv6cmZ9BMFfjDMz9ymfSRy
ZgfiyM/tQBPx7bHY5d3B99Qw7J5M0YMKbFGm7FITLtIEIv8hk9QziPpWoAC8lepo
oUYmqcLOGEzPwUsUIRx7Bm86w6dJH/JPHksXIwPVUbFs6C0nAKPzZ+n/aY5Qnvkk
AtC8Rtbe5XWkFXu0nYjl8zZimd4iAc+G2JqooCOC2evHYT00dCxVYm4nVM2LorT2
KBp0XCBrHj4KSgFf9+dskYB7cGWmUITQaApjXQJhy9OEIMhXfhvzavMtTQCLZjRq
ebv9EzlA8nWjJpQQE2GjN7FV0auub3Y8mruRoXoxhkvB/mtMVDLX4JH1kKlJnKAn
TLNStLYII8XlOE6bNn3Vhgu41ZxBF2adxV1asbvuuq5dneaKXMP1mlddEbZekI1B
/FerU+ktpaU5NkkCdReXJGvVFU1cQCqQnGU6x2zkZObopodx4EBP3zUykRuaWl2Q
pVBO7LOYI+DUqofb0bUakQO4PIT07zxhyOG64MycC7sa2Zkn3lyPuQwlHyK6GOWk
XGMaho+p4xIrp/tUV7gF25nYfBluDRQTFzFJBA5gChN51ViTnz1lJwzlkBs5tqmG
iQ9UcmfgZ4vtBSrmPaiOl/g8sDtCGkhY/ZkdZh4dW6xeG9v6fySaupRxS+4aRRww
4+pAB2YWTPJJkOwgWgGcTBu4pnFr9b33scAOiVPNzgr4YyBhw8SaBpr6UVCcaQTE
zYkhbZnwAULImIH73j1kMPyZodK1OZ4EbxQqAcnSyLxh0az4uYAq+Rx8UqCaK7qB
L8anYa+Jwz2QAfraaNo52Ve7lPc7OsCT9Sk/9nq49JMxHJtp5jv9wY0e+QdhItUR
pAmbvHsUqbZnE/EsmTkL6RUknwlLw8/tdH3mLQE5kJo+/R2DqpOgUURr83Cf75SD
QbPJRCWi6OwWHartuoB+ow3vSQ74x142yHyn+vDmcGCgSJ3W1EMgOVSxKxWvxIVi
Yz+E0yQqfw8Rl6p7GFtqyXmzKGNxq1PE5Mxk+giTqeWVwIp02t7jLQO/fZNKmdhF
UJiaX8XEkc+vGSyPXkqrjq3fKcmI6O/FkAGhGU22+tU77HTDlTeiV+B/+9eRq6BF
tUtav6Grdpgi4tZqdjw5YAp8QNK9cVa2M/zVH/I9BVTyVFZwtXue1OkTdDU1K17Y
Jl1UMTI2hSq5ptFGSfL67UFMtiDBEhGCTkHWz7KbqXs4iWmiTXem5jwC5OSmUXg5
ecMzkh8aKnuIHuZkdxaCvUgISVDio7qkM3IOVbMYfunB0pn5dxjdW0yytWkD3DEE
rJCBTjg4iLGAnaY/DX7nHHYaEHUpk0srtUTJwuEf/8d99qea8+YKx177JEYVuONG
ryeOy8ru7M5zVLF+9Xm9znzogUTDvsD4ZWPPOAKPyDtlIWAXBPS6U+cVzt1ks4eW
3i448DXKW7lPX8SZj/0enwKQSVxdinGSOLmG13uUaFFrdKB/b8urHWHh6u/Vz120
z1rejW55/xBf9b6PjgA6AGshVQzeaDdadPuzF4nDfel/QiIus92hhiovad5mRW4m
fCSB0dN13ML+mnSID+PVOILJnkBmqlT9/6tcZJ9UW2rFZrgmn4GHky/Tc6AZgF0I
CfRYzrWgOysEAjzj6XDXbnkP4c88IyAtvFgGCS/OOv9Kq9BZJlCyy7ZM8PjwzSFO
n3k7YtV2CDa82vW2WPhCytcb3so+CqB8NkuZT4vC2N5PSnPaT6wWDbwdvmxakmi2
dFmlX6kDWLjS1nvMyot/Zi5mNNHS0UKggSxVjFT4WFAUIGvBX2Yqn0qJXHoVnqr0
qn8ID7bfBuFxAzyuVlh79NnUszhNzaQZDUzC81Jso7NjHwRCbXzfZgZt/jDKFAAW
RwuRx7kuEXQOR4JBFp+oLDvzki6X3qarA3b8IgtrurU//fVWXJvI3mYDm0n8ZWBe
i3m87tMpbdQ0492U3xpfj8EMrKVltIkn1txXpv14twlTlomk9m75OSTVTTp5ZncN
s0uf/nBERXd5QWzJAwTpm+HZ7aCjcKxpK8Vxxz897ERjZkPA+S5hfhzwyQ05MXzR
cMIYj3SV5t6RxkgSuoffZHx+uy2WRUNcp4KVXUPm7Z3r1YoifDyRfAnEkxs0Cknq
9TFyBKWvbWhb+l6591wdmttwknDUTxToCrXr2BEEnFRL5TS1lczdsuVHoAJKeUni
SZThvLvlDB2D1pUbD6TgCy7KkwD7CirtZRjEPBONsPs1LH6KJzr6MsgYx2xBwxUN
g8KBozQ2S0XDmRCcXzI0946ec2Eb40//oTap1559q/IRUdQEcm/EOGy2kjFijHMc
HO2LWOzsOK2zbfWs8HijRcluljv5q5Z6K5qRwqp8LBu+5k3YgqkkmMGZE4Xo0RXu
HoXtsDdmnZn8jKJuFx6nRH/iaU6MI55TOdNx90ZQDa8oo71/rwTq9Y4wtes9lqXN
NstuT/WGdGn9muv8FR2RP7Tv7HWjLHRBwcuJ6O6TKHhe9UYVrA3wFtQ0vpeMyIxv
hgcAaq9qZdsZUvmTRvhuAeqK3ZhMRlgOOUgH8JYXKmAC8ETvSOzSoGtXl0eO4Iga
GwMo/KgHGfk+cy/o3At9F4tATefVSrUF618b1U9yQ+Rij8HmEL/p7MRNMIRa3Z8O
u/YUFPYoeiz+w10YF9yxFcSTEE4dVaB/kkw7s6Q7Nt4hOdYh0L77wn79XRIK6SgW
DCnw30fLbXqaz0lKZAQbnO7VJDeHsT+RISVJYBy6q/ldp1qdJNJc+HRxbWzgQ+RW
LnE0vdub18dM22EAnsqxbHoI0wF2Fr3Up6zs9GbEC4BRCOVaVzY/kiHaL+M0fqIe
xfvnBAFSvMHm43bARwTE8zUUV3ZYg3lE8xI9d+n789w/9JThH8hYA0Qayb0cptgx
hx4Q1RxCwUg3O+apzA8JdxTVom2ty0DRQpFJYF+lJ1QqaDSgcgpa5K3Qct05iSku
jgnmE/x0UBSvQP/6Oujtj1Gjgv0++hMVcizyCQRt3FjuhU2s/jsYZQutqWJMJ/WJ
oZwcVUfL//l/SocEwO2+MucsfifRK6DwWlMJNS8v6ImM3Zl2iOfiBa+TiL39NBtZ
9DlmM+JsC5E5jcbUnqur7O8voZQgTPxs2m58NCjO7oCdTr4fc7obleamPwDc4fgP
JMb7ySFv0qhcqWUhSya1AwC2R6bufkPRP5oywaGXibbMDsPF5DVToq3nC7Ev7nxL
FjAG+Q8oJA27cfDiHe8ZAGQe+9nkEynhELgpibTs+srmxpO6VQqXk62bQTs19dQg
YEJcOv6d0tKXVvcWb1v0T2CydXoW8B3cNrzzJG2R+U+XwLme3Ed7E4Z97KZL7eWu
qUSQG8EoaQDgeEH/MpxyKvwOPAQ4v8npGLFSfIRuxzg3Lt8cDCYmz6CAciI70+qD
rpWZrjnBeHCqYOPKGgE/7N1suv1vdqviNK2Ih42hv/Jm4qQi6nx3rePlYjmdVAul
+zM3U8Bq+InPf4lQf82h7YF1/52qvFMZxSbugdF/RakQIFSVRYqQQGRc+muYLv/6
N4Ly+BvLKFH69ZFOgPCzN0qicXXoclDg3CDchnMnQUMYgi3LJ8IrN0XMAxjqOTW1
y3zmfyFrxX7TFL1GaFNwhnu0r+nrFH5BpNaNVyiwi8OI8zRW42gooQ5syex8VOEo
EgYh1X60csks7KkW2Oc9qJxl7Bxe6WXIYMOcuqY8hWDsADFesSXyVKW2eoHDEw5N
34pbqLAyVYgWOXiUXJfEj/TDIsZKIHyZleZjGk4nEs3qXU1QLCK+b4PG+cYwxoND
bLF295VhInSoiXUeGg8cAug/j/OzXhlxtY3pxlr40dqJkJPgz+2KGGHu8X3nb621
d+Iy/JJPXTRG03Lx/f2sMle9V3MEB/cD7MQT79BpcKRvp3Y9OFKw+98xyrczA7KV
UbgkVD2iBFsx/X2k5eby9yDDP8CReTfOAg+z6yWgSvWd4AGudIXxPanWMsviAeSZ
HcBfCMLugMN3V7DYm3+q6sUDwfClaka7XqmO7gW/V1wWEE5InFHkUgqEkdiajGUi
tR0rWjvfMGtALVi8l06mTKZTzJ9gxUEZvSZ3dQlj8kruq7dWrtGobVPvPQpGojGV
ifHNxE1DNhh59Sg4opSF0NVq/x3WuXI+pNuQEjD6Lt2oGSy3fn08byMznwnguAZr
Emek+MaJMkGPof7AVq8iyn4dio9XyTpN4SnWAOV3rktPBzM5R2dYz54YzeFb0Vvf
WiNcc66FqOGG3Hwaf0OlwlnMGGGjxkTf1MlCnlUjDqFTfNVGS4QcroHBmxuuQhZj
TJQVZTjLpmcV6DtEYmIDr7f40IS59mMQKyj58qh2YoRtnGZ/iyAL8WPQsvAgSk2A
kpAP2tSW1h4dhfs8VDuYL3zcZm2zzcQiGq8DFiVQEShsRmcyBXJ6B2EitVZO/Wzx
5IPNIzZRPVlQ8kRsI8c0XveC5rBmRWDAvrI0FR5Oi/+1pt0TOgKJWx95sEpKrjEK
ZasfnMjb4o4e2JiuPjoQuHN9d40yZdzsNwwHH+rFMg4/InUY2PdF95DuhhYteq6C
HDPUIs8wJAzJKix4+kgwXyEcIzH+ylN2D/Fcz63lK5A+Cbt25czSDspDbMRGGp0w
xW5Qec/FHHvbEztzkrgt3VkAREVbw0hAfbemZxKLw8njy/RMbxrD8AixwzMKL4qc
aR7g1IAArh9jg1GjyV44mBzevLCcJ9mai11yAo+1ZbaYhK/Rcrw/xTbK0UYkMggY
hNAo7LirTfw3kt5sio0P2jSDk78JBF4nI6dzTVpsR4JoP7ODEeHnpXTJxIxGGgK4
igXNIYUlHsE2DVPnPlFdKW5hdZmgfcuSjElbRJAUqyrVtYpKhjpo9A8F42zDLBYh
pqlCvJYrFm1XZOaJW74h77LMn0VKotv4usC+sKQCNIygF6gLsqp0LC91+RN3cwwe
YymWKkJ8XEgnFauqgOhznbAbgpdQujZXLOk75Dx4WLS3N9dnpX5OCz62IS68+1I/
fgSjIlde08hYPfc1a3gc5PAhzPWkuGIU/vtNegy+vf63FhcMSG/b62dmGk8JX+/K
midVvT0h8cRqUBT3gljcS0/QSUxExUVYTRn6Z7G/X/MM4D4CVvck0hMAN0wrfCut
gGG6uh5zYx4S5CvrBIJ1f5UWJ6Q8aQmSEAoNcH09rNZOxzqr4+CJOh9cVgoOwvhl
0rnGfXt7g7ald7ka7w/9G/YHARbnX8swPdvl2OI3ESKTprwvUvA5gNsBFVoHmbOD
/swAki32T6RMeBq/iCc+pNFJMM4DFWD7h8K4nTmdBqv4RmVWrg9b9jBheugaZPo8
LXemY/VgvwRmSFOgWh3GJ3ObPV1zjMoXO2eF92cFuFDfiz7nGLHkw7tHAPfPenSF
1B6ZQPvjNAq2s2qNXeA+Nnp5VxGP80TpuMcKrOp7yJVHPGQcGOyGNY7qxaxXtCkn
wZY5d/fFRhbPFvQH98QVoFzf8XCnQsvFk6EMPSqxs1mC0AUry3z1jiYatr192Uke
3KdNJWXneQxSUTTBTks2CpZBgXTgXSwXXsfc13SABwkiFi97R1TGfM3FCYMg4vt2
U0WLAvlkAr2He6eFiTIqePm6S0OTPTP6Rjave3oMLTVweypAUQXacmhEzy5elKhV
MQbOjtyW1C7mMjYM3nzBTt0pd9a4Bx5OQtgaYs6nOjf1xwG/M8wgD/Zvr5kh+cvl
Wp1wzZo0BlwmUqWQ4CheVmH3qaNY8UVCRhoo/gWu1v2F0f2LeaBF6yE9cTmhx1qz
zICQanHjhEb3V0yTfkhA2Qt0qahjJ2KoI5uI0x63kk4sB87KHVlaLvGnhC0G5QyS
j5qf6b8Z1KJPR8fRE2+l+GTrmWK34pTcDJVHzMxZmSnmBlVp/jnw+L1O5BuYocmg
ID6Z/97UuTiyqTZixg6nWGQdOlZy3DRSQoeF5+DiFivzErxnsHwsUISwMYX9y0og
+SaE3+HhwUQtBOUqgy/Nide+5PIZ9NrzrLozcmqqKSDWvcRvwYZkj8nMFPhZGt/F
hOK/+LJv/sctN/6DnKu/x3VFmy2YZeZC22q5XcIr9pq+1bXXJE75dbi7qgT4H0Sf
Kh95UUcPSqGSv63p8VTCkCAY3RhjOyKDYioyklgseikgjkR136GHseZLtdJ/GU6d
G2+3AxpeOB3XauwAtn4Vmqa60iqP9Gh4WN/2t3ktrOKbKFC4O19W7xnP8iKny4f0
rMtfuRsd0pvSqbD1gn6DnyTMv6PTHr1rtnInjj5irrGUq7/kYD2qKnoR8jFPlamt
Fu9czRdlk3A+9fCJ3CFF1SjR+1UfL74APZytUNH7XL++3jjQdKUN+Qi7/A8Agbws
a46oTE4CCjUUJw+xUD183Ck5qf8PdQGRmg7fUaYIIe7U6sXNVzFPOk7KbIrq/qx3
l6pABrwKBoGaMcQt9P1N3PO2swZWh9uQXcKPf1UWiF0etPqDbRhnyqHwQcZHeL96
3CLPYYVdDmIjLbM1MCAjjagK2xsGMw8pdm1toKdttBDoo+AnUwCYOBUGqOeTGYER
UIF7aBYLQd/9UI6EBCilQsRcFx/eteBBJ4teMCLadje8rAXOVoRhLke5w0U8sLhk
OxyK3tLAlJHxmU2y1kALPVuOhR3SLF0UC8v1rrCa6jrxskwT2tnxjb/nT8M7sprH
xsiuDDvvYpMR2baUk6NVfEiGViPhSeSpw++MXO2j4r/Voj6o3BROgV4I+HOx2XSC
5hVjghxfZXXJQEFuSDlI7BAs3u3YIcSqpbxe27M0UIN5TuhbItAzdBxjjPrlfyIN
Ejzu4lP+E+aYRP/NC/zyE6b+AGj8nXoZG3kSwXo15KkdF8yVnBx0MrEkKdr6W71a
jLctfs4dQgti60gJcfcZo+dgsHjFlbpj0jRsk60OaR8o4VV4qLbV3W57neURSHzm
zRf8U8aZn3hXTPLfKfnZ49xFxT9d7TEwfEDjwSxE5jGV7r8Po3NHCSNAq40/y/fS
h5AHG91zHtphMJwqq1W4amXv08Qldkgx5vE/O4xkJvJXIedmACNYUx6tQQdNHzfv
6x8KUo3HvN7VKTfHc8/PX1VAba7Aw2p3NKr6zzxwAkwpczBpMn/3DaoQinJk/DaU
7Nq+q6vHn8Oog+xX840uK5wv/2FNHZyhnYx9IT+UPt0g7Q0XIpcYb7epUJhi0ugi
0BlzlRoAgn5leONB5HmfopQKRbCsueFSCYkhrANWAfj0hzVhdAtwXsn6hi5fan0b
rw1i53w1YjzDwzA7Gmk0u4dADeTVCFiX4z9pV9Y8Apmgj+kdsZsOGMDWRcPUdYdj
atBR+rHBonbD8QHDiiqsAEBweZe5DhUVXZD+Br9FImgWMemB6aR72+WcLILk6rpX
EnOHJ7aeWOChGh7YW/+pXR3qA9prrq++OqtZgaTUxJjALmkosuYB03UCcGq3TvuF
ncNyaUguDU59FSXPqTIknYzbGUo2Y+Dd4ULDCi3zotGOzlAvBGQwGyOXCztXAadI
HP/4VE5oSv1nYhi/2mNCFH03KZMwvMzao4dgi/IwrgohVg1sQaRmXdUESEIc8s0i
Ng8mcMMjmV7eK/5rp41KaNtw4m/WwgJMqZ4WNtZE4QfeWB16ShHlAfvsLxT9XtUI
JAfCfyk2Aytkpy5DWINtW3CsauCoG9AxyDsh4GFdQXnPfXAhyTJbZAHY3BTFgVGv
m2JSvYWbiZbgIF34Kwq+qQhgSUflhdrPAW0kBWDF6ItF94Q+TCDiXWCSjsh+5Nle
ISqe6BLqx36kmTirwOnZ1aMeCBuYrRqDrBmmjD2SxMD6mpGJI/H11O9ajfXYtZa3
bVhKLyoDsmqds1541oMZ70D1h70vQVS8vqICHgHJqx+KUWDWxRyAQ8DKoBOlLbtt
21MLdl9MJ+cThhCEJlMGm8nkoJU/U0e2Hhw8u9aOuLmZCcWeSmIF8f+vkmedlzUu
XPzMKB0smsr8Pxi7Gq1LM5FgFUCeL8XB2dV0XMUHPm3lzFMpyLlYVQFB1nr7eJ/h
H+J2fTIA5P6lWC+QfYrAww+mhK9oH4p9gZG1afxhZ5VUbkKiMQ5Y7DEkktb65QHi
7e+9xgShXkV7IWco73ic8OmiD2joxW2whWwv3PnhVP873vezh01gLvKREhA5MB+D
8xJ35GCebTnRqgJE2d5d89jKEOMo+OV5Ln27TfDK1ovmJ3Q2Z1N/h6iBqxI3Jvw5
NWdOB/TL4h/6Px85xkJ7np9XWKzCdKJyRhAXbnaYzVABgngQE6c4t9q4qK+odrCS
hkCD+mcUHwEIxrg/roWjR/lqqW9R8QJ6fof2IXwx/r8V7zMDYTCJXGeTdh4M7I2Y
2WAyGPiTCewELoHvvVCCasmw4L3gl7l8gtL6r6mimGzy775Xc+OKoZ9dg1nEeSf7
nseWms3YQM26UEPELhwganocZI0tEDSfngmm2FNOaI3eBughoNioQmoDFUJRVzYd
TBA65hLwImh6aS5dwregD02FeDjxrpeET9tJnFxJafJbNkxjjMSKvzRQyp8kFWRT
AEBFHs21IBY981iPaLBXCETVOAAfTQzz7gfhOj7G6Fst4nspr2pc3pkbiHZah9g2
45NUxcUl/sdjEbn5nZC9a8zzhCRx1Dz6W8kFUohu9WZvSFsdrEMMvoH7y+7JqcWD
LcTY7JWfbArdrCgLQvtRQrxmt+ITBR/XZYGkYhv+nhKUq+uqe8bnXKuz7O7PRwa0
+sEzVoUBLvY2s97LcvoGL63q4YLUdCGS0ZF/bf7f2iwmNCZCCHOnFP0mwiQaBNpT
od+o7dwcikTS3CpB97PJ5GzUvxXb/0/xxwPyfvIfXocTdZIh1VDkNHhOjQmWAEi2
POXdCW5r4duoW4Y2RLpPZhVlzvL8gzZcr6YzXGxgk+jkWmpcWbGbkjUL+lNkWDlv
aOp9/VtgW/VWu4h4rBZ3OJ2X5vo/D9OnQYyw2T6prozjkJe35zM2q8pMWR3nfNd1
QpugCfdS2dInOMrhYg6DElb3t7IB3iCG5jJdKl8C0MdW4P5Zc25340Xs3aR2YeRm
2W21akNq8Lfn7Dl31veBJnEV0VwZOvspD3abvoFwbObbjqyigOpGiJ6MXkeCVrDy
Wq6Z51jbOD4d6zVobN6lJt5MlGwcgauk2Uvm8Lnnc6ndhynk42M2O13Re6TSDP2/
8gJE42DWyUY1/AJuUmfOejuSTf38j4ohhajIb9SIzJjPKIgbyzPHt8YOL0nMp5bq
r2cOxZB095cyA6+egw6yaE+iIpb4hQqnlXt94ZBJCO2K0tYsfzP+5g1XK7QpjyTE
C7UAZe8aIBTiRoa6A6CqX0WBF7ujEUVJV4kY9xa778TTFlhy7XeInAGdZSz3Xnrl
HF6WY1rjDt20WsswtpTMF0kPwkNyjiTLoBIf/r6FY+FRf3TuAt1dxiXgneuJUwyf
ybUzytI06L1UHLtaPioifHBaEG0G1CS836zNT10q2LVPM6HjjG/InJZWt4EbjzO4
MTdCK/EVcUu9EDbYhCR7Qfofi/c7xNbd1pG5qD8fHLBP50qCgb4tyR6glhi7Ttah
vl6Ld5jAxCL08JFr4IhV8hktyrjarYiS1mGllRjKZRj7BJVcJ3MpiqVb3+I3utv4
bvOlNv1fhhaEzbvN9ixRv38Ka5lDEBHP7WmlFKtTi4n/a57FwRxBbud/+jepKSpM
HoF9z9dZQhLENA5WU7EaWnbs6sbDFsiWrWDQQKv+eXHz113TTHb3d++4kDPpVDfQ
f3oMPnJQxBVzOdE+Mw8RFtAxRDXvsuHYD3jc+8nGaJtP1LXqTX3LfYUpBxLhQCZY
3968pkHYxaEQDAiDN7/R3/Ym4HmY/LjaK6hy4r7F+UFGOiQBq/7eMtGF8MIveRF7
bkr8FWIIEhZWmqUTF8/Py31jpzN0gA18y7EWm5uUWKBehr7HlOV88CU5DOQPZAmR
T0LcsjtzFKfqlNEs2lIkzJrWa53cC3oWUkiiMpXEYIgX0YgMQXAqBbX3QpMp7aDI
9wM3ZmFn/2nptbpB9k46cD4didoQkVLRgjIaqdQWqtV4a2TV0Ymytpmvh9baY9DS
+Wjim3rRlsA9VZScTGLNko2Sb60w+DKAF2o9BoyYUh/zenQCNTY0JEuf7DMdOcC8
Kel1TNd3resqK27p7VydSlES9KJq9+FMUB+fS0x1UDNE5Po4189nl5U33i3yTo6W
gh5sZWITbsmhZ+Tp+3Fzg9HDs7y3EcvhGOumLUpn2GBG5DQaBlndzcaz8esk8yU2
RetZWTq1AkyaP8nPdsSYt+YHJz3epWzMnmOX1Q2yTkAvRmMlwBYu0m81lH0yyMeX
iYJ92MFeaiLSkpcAMATyLPv0zUIgzJjUsAOljSLTsiYAr9hURFnS8GhMLfWX4nHR
yMRZjCbz4hLns/gBTikSr99JeEo6ZlRg9Mj1iqDnqKnX/24ip1dl9oa0D2D1NVkE
Jfyz2M8LXpjQQ9Z44ocfdt1cGFY5KcviMLz6tlLNiBzbDWAC1kCHesCArQEPw99q
K/ABICpvp1kL+r9tyxAsIp2R6xb2NzjOcnfefkfvTQMyhxzV4a+ndOaNuLOlVSrZ
HUwEOUM5U2/tR8WBI0OKIUdI+mzfDmG6BcY+bznypu5caoT0vinBJSYw6+bB0HHi
5sFHHKQrhoT4w3TGDbVxfS62h/ZDMIWrKAtTdeTPo0+zCRK+3oB0w3xXohU4X++0
ghZ2Yf9/Z2gSPfBETHUmpAr1BxMdNkh657XhLIS30dfP6S3g0dLENh6vJdO8jwRq
uYIt83Mq+Ycm9s/sxlYVBnsuaebgKE7LEUNNQwiG2b7n8p5NJ81Sx9+sGu+5ghzK
K+v0TORA6ffNmSYSiLLWndDzutOGxDsYIodSxa9hXttc+aCrCL3WquvJgxc/EIzz
JCI/gP/QFzWk7yy51bYgQ31VkkGE9RsPPUY34s28VTtkM4fzuR3EeHQR/QZsQB8x
r6w1Q3pY9kCcimYVr/Lt9MPHZgG3jaQOoxr5OsdhYS7KrvUZ8A51Lo+sBR0XyZZ1
/77BZ3dm21FIGZBs4DvCC1Lm9O5WIBRh4KNdrL99y0hfa86BAMB7bykvkMk9RhzH
gP1rz3JCFGeTwWB5jAK+WNsljXkLdRj9pztBrEi0Gc44wkrjFKfOKasrwWJ8kNO7
UVfIfoLRX2TWJkrA4FiAZQ4XZPa8HiMc4yuuNEHSmdhIMvrZhcQEz3HHgrUOStp2
P7HJy5VZB2yG0nGEbdtztSPyKh7aoqtExzw5ckBvp+7dt3FFl2h6u3NyRHxaR1Qa
mKOFRI8xqAR6xjpfIuElbuY9CWDMAKcdMXpTbAtH3P672TJ58DHzriL93WjD5TT9
10Iq/USNhsslQ6k3fLJ+9/GB/C7Z4MkSxL9Nv1iFRZFBrRqcqdcgJD/6cBkOqD+q
xTz1OJDxZOJKDVL8dxRUxlZqBQTSeD9Vz7g+PrG+eXfVbEoXj8z+4pSPOgpD6Ck7
HyQqTSCM4lZS/ZwsXBc4FSOiNdOqtTjiEeM0MLLemVBO7wHysibHvpufEeKN7OC9
iqflRjfwlZNZomXZ5UgCj7fbcwzcsraAURXdCnMIrIvrjFE6GiV4w9xSF90dhPPX
nmHNRVsriZonF4rXXN4Rr7HOr4s9Ad+btS8nz7tW/VCi3TCT9kbhj9R4EEDN/GhL
Ju311DET+BKv5rG5BqR/kzAGQqVdmtjOmUNEVg00fnu/o54Rev/sgQbTpaODFsqT
ixA9ONvVhuuUAMLLDzuBcs7BS1zQHb35Grjo2T4/HMsHFi9OLuAmTWu/8h07x+3/
nQfIbHYd1paK7AxAmJfhNy6a4cmRSF2B2f8y2Jgnkh30lYivWAZAlpfBKeUz+gbW
ge89GypeNC6BxmLsAAZkFINDk5BgdV1RvX9RRykulDD7fqPzOXuGQZSS6CDRHI2u
yB4avwR0c5NP1kSo+COntDYQaUtq3HZkVN0D1UJSiJb6CEO+BG7TCxB0pKXvdZVp
ZHOdp/C8+OhTrqBVT1XbGeq97P4DFFzu4DUZ6I5cSSAA5/47Z/lErpltFnBaC8rH
eBIJpgoinuy2wh23SztWnJwjo0nWegM6cPqc99i4sYWVX3NIJt0otv/2AB+9tgSl
3W9S6e+IxPdTyPJkPKMdrtfZWuFJs+gnA3lp5T1e+RIeEEC9OXKr6zsfr1Z67aPi
EycK2l76EL8MKzUENQefn+rggyl77zKDp3ORb3w24NNhm4azuu6EBpOpb5Ic8uUz
tmn3JSVA3mmrjBtjL34rh6QGQb/eU61tMdlZuY5RgEmewFIxISBCly44mPDYOM+D
z+wn4w5zyu0Ry2ugJWfdjwwq4+ykxBcYdEMEczQ9ztiKZ1PvWJhcMbwYI9TiAIAH
lu5kF1lorXoFNTqEcpwOsSVEEVC/i8TVBA+Ej0z+yMUseg+GuivziSq32EgfplpH
xiZb/REDyZBoA1hLhhfpci52ih7AwYE9NCMNRkmMuw0IUu7GJP9c3Z9UEv2QnUoD
c1WYQyA9H3dt7JcjAQ2aGozwpEpfQC1420QsFpzEx82JIYtBrq/Y6gzxX0JZhrN5
+UWif+4Cv45FPMLSpELbbbDnxg7lHcmPo1hyvbtQUCSyM5q5NTcDTEATnkGYOtI/
XlwZjCHFjqvfi3UieTyY95Dtc4MNkE451BiwkP6ybp+uGV19FJQG5sWRrmur8HR3
/BuwzHpmfUh5Xdoju8PEclO874X1xlzheFyv0wqXCRr3CYyCXbO/Zi+AmtxBnOqk
2LZRoxiUlJlTf2WNJlxyF33FBtW7MGB8KO5jKXswn8UkVOaIOlWSfzgRvyou1f2z
JSEQD/d/NbQYhJ8fRN2v+IaHLSUBf8b/pYCqmV8cHxZG6TzVas8kPasqgujujO4v
Z1R/hrfQA0RLCvMyUxEGCrx6wzN3am/pzjMgLz9o2DUpYzrl4+nx/kfWJ0GHyU45
6fJN8/Z278uC1+NWIcFieeg7To9brQI8ny8pgw4X4t/RULhwWqvafl6J7CjsHBrY
fLDtxilnt4fTyixI6sUaOUYJ9q7HuK1N5Q6k9rZBUx8U2QfWgu0+22LRxPYfQTjk
31FU8u2UhH0xbnmssjo/S+c0Hcb+B0bd0RCswkOGnHIBRIT9Deh8SCYMitJMcnsq
pfx0TOCZxP8hzbeFgXaeH3Fop7wJXfFvBWxmrHlkI2k8+bEZZyt2u9j68nNeA80Z
Bg2MYH2BdpawxWr+7zWPh1aXDiUHK4+/2DHej+0807SpIL1/iPjwBWpy9iDIGMoS
tySM5e+3anOqes0mUnlvXuRci2efH8waz7LL8Vo7XZHnUkJXowAzUrWzwi9l5TQf
8MROSasPEBLcnnri1kw3sqSDcWsP2CUogPduNsE16CusUu/994QQbMOA1KF4Ukmu
N1tpo4GnaPVuyPka56daiFr+5huqaE+HKH2RJ3YddhNtO3zJg3xn3Ga/KbL88YGf
+8X5NC5Oig6J7rIt9Jqm7B9RwU9JgB36hX9WjT4/5CkG5bLUi7fHAsxNL6krUbNY
K3eKEskr+R2rE+ZNZXr445twIaNc+Zy4ZYBFK5xFeoD78RsmYXVkY11h6oMOCSRc
CsmCcANHlq5dycQhO5j1xglcZpJBPNLYMDof5B+bvuwqZ6goApAFgfG4Prelto+N
+MWX6I3+uvkU8vsdJ9f775puTvZImHWRF5G73HdzJhyoupn0aIJo9UTH5TpBnhGP
fx8UCcGzsmG5mEDBaiQnZJ8rzthN6O3HbimX8hPv9oVeUUnvhOCXx9jQp0rTDU6M
tnbDUGvMGlzl0m7piqQi2P/gmVoTS3L9aHDkwGHvZ0VvtF5nIgsVT2hLx2KywPbC
vvfT5gQKk7XAp5R9qjUudRdLv39ZIpHt3y2vNy1I4YFNR8HOwnNh4TrGJVsVAKzq
AguFlx+j43RhHOEB/UvFHL+njhwLEDN2/1lVtmql7yquAJqT4qcIk4Inbd5723Yg
ewmO0MbMQGoeuPoGt7T/Ykxuw6wCgLnweipsEjxH6BqFH8gFMBAMpphVfRLGN+kh
NK3y2J0BYfAnGxKgctJBsLXQeFyUqs0LoSCtCEZnWtxXHCekkXljyNWNXQ7WeNwb
11fJkXro1zaV5cq+nhGoqy9pFwOtPoY5nMv/irllzKiOsIeN8TVSlW9nGTjwl8MS
inrT1YwRVld+VtRBYV5if0Tz4iGWQYji4yOnUG6sVfb+yO6IUfp6QNdkh3TJygcQ
3Wdc4aEgzabfqoMU8giCyqeW99YRReY3y83ZzOoGO7PqPwY0xWg4zqiBAiYni2U/
cnU3uRlCS0zSNPPNa+bc5STIEn8tQ3ZsqxGJrI69cOm7+eUYVAYNwup1wS6fu5ia
0y1C2Yz8P0xyP0Xu3cQNbfn9yMk60M6hSNneiD/fVXear5kJU0IMGSpqmyYEP9KO
M9SBWxXrN0ZS+wcRokFLdyK3Aem4lBjSEEGwO9mr4RkjGxZYtaafvmBHOLrO/Aeh
rrlSLgJERfOicapNBzFTMu6qM6j3C4dkbEJOzCg0UL2qCHcuwweTlKRAhmHBhgNj
lrwpPl0VOgeMUEtZlTzjcSXy2sLj4bVEf7uLTzpcuYiOtLZxTgsNT5ce1yk62v/O
8cF62stQIGSPfAgPjPLbaDQjGtp2SyIjwc7bbLW/q9cXbuxTNzsGRhUpaEyYqnSl
XLhnOLpmecZRse/WNKj8BuHevOazHkce745vr/QcmnxtlHrGuNWhal5Xdb8HDwhv
JDrc7DJR/8gNs2BG8DKDJWtd+lmuhT/CxFaxpfWzOlj2hfyloawAm6jjvUlv9WUg
uaErWwP9Pea2u28lkSjTjSAof6oJ11x8wVxODrNJ+eHpjLYTGWWFugoWR0WIwtVO
P4CUSp4HB82Qxa6CUfIR8rJkT2RCge18m888etCPdyHKUo4Hz04oj9rE1mwWzjwU
Md8XtsEO8bmVclHyraOwBOskX42KUWdEdr33CGekVxXy1KPwBzAvDpJFetgtrf5c
8CV8u4WyHBusVIxrzjPgnSlW8IZVi4bJDa25nwdIgBXlAoBREz/YyYTqwHXrAAqv
zSbaV0OXLOzrifFO9knyOFx/vDLnKyXLalogaQmFhQW7wnaiLnpM7Bl//N8wVb/b
IB/FnYhm4AMvB3d2Y3bzweu8urguQPFaaqCQRJPMWcGszGgCS1j0G/vDYu5U5bUo
i5AVZ5Zfi+5zWAY61DlIKk1fR1/pWzyYe+9hQOPZZrzJs2Wofo4ITAl0q7+ACaaI
Zs4PL00LQL4CPCFIKqNHpwmAE5ZjrSsmcS1hHLZax0ECBQPTIXjSngDh6KD0LrHC
THEhKRUG9Qxmlamw7pyA9yBpcQZN1E7WG4nCSgt/E9CCay5lzWMlgB3j3EvK7kbA
5auUEaCI+DNjPABYT+ZIfBxgP866UoIf7blHB818VWTDf4FpJjl34BGWTtawsqme
1EAgVzXvpxmx8RthtOIQHuhfdwPoVk36GPceU46vBpxcTvNac+dWh9QLqdlYM/lY
GJ6UVmDyWAY6pv64IFCVoBK4PE6fEzqSHQ/OjIE1QLKLWrcJ+TiD6zNCr068VBBP
e+DRlXa3mdUuqpwhaIcMJq1rIGLSg3f9TtozveCIxRmSd1qsvUMRSLTFH5UK0YCN
BlXYOVw2JX+h/WK3iDz3hnKXjQKeU6illwHoZ54kA3bdsH50JnCruE02vTQWFHe4
d6a8a87HULlMkuGjFGWPJu/Iq4wTL4iTgMUdTrPTLrjWVZs8X0cf39o6tPkIV41n
29evQRMRfpJMNtOMA3Zh413sAMMzXaOa5G88+3zHixFs/jAfpmcEyr1Ysmy3yiaq
MWjoLZ9HuYk8iBlvfYX+YsZglSNIB+5rvDZ6L4EkehahC57afoGAQOoncAiyfrQt
QgnvUaiTbym0gu+MA7MDdVSovihn4TvorbiTg8ETx1d3avXvXtkEzjTSb7sIB8pd
DQel9WFvOvfq6zxkp/Deqim93FkwykcVJDUOjqzyVEPUdZOnseI2CID8MAAfgKfr
Oq95ZLUmTfOokAhWSvsBRva1t/C0Dbu1PgUmKFJY6t7h/KhnFsnY3UlU3+Kcjdjv
jABnMfKC39oM3v5J2v3/b+wuT1DONF+CXL3Ixr/JuSZP4/9AIO1g512klGyeiedv
T101+CbkZ5CfZ65YlNJ/eAcZfsNmWlKJPyT3zG1wEsBWScZrkpuuERRQPeMC4hWt
7NH7aQzTi5QRQwhoFzkp+yhCjah1VqiiJQlcW5xU+bPGKXPKLWR4oy19rB5OW9KP
Gf7ycgg5+oBa0jdsc0l3gTr9U3No1RP+KUuDxdUS5pRFLfYV6fW+7pSB/6M5atxV
JumOtPJPAoTKa48I/2nTHytOi53rNB5gNgLRTjhE1Lv2LoqoYY5oBmZDNcN9k/xw
vKgkdydOb6jbqpDeyTMzSHPpyc6ECMeAAjct5N8SdSL12XMO+zDeHdHcCKxTmDp4
D5E+91uajCCFG6QlWJdhN9BhGdx9zBkkVaiYTm5g2y6WaMqJSs06E2C7zi6o8LEY
U9zQL5MDRqlf4XYOUulPuGBb+JUjkLA+8pFr7FzRETTwGs92ltjke+qWsaQOZ4Hn
n47wqoOdf9Tc8U8IMGXGO1isqgoWgf+A9/PsxCkZXIEw+kvRGBZsQwAf0fgcZ+tN
Rb7OIKXLoTkavugZjsbUr/MBHBFeKFFrw8tc1hoi2QHuowmOO5oyhm7Q/a21Iqbv
T/LJdpsXceW7uBGm/A/iF7T6sTezbEXSL+LCtZuP9i0r0No5+8XwZVl8gXC5JwW+
9t3wVqpZ8B2b/suETC4ZEu2T3zSuYbSz2R2gX+VMLloAhVirf8Dgm3RsVsjiwpHi
ROvsW62nh8Oyci07tSkQmKFvq+6WZl0A+ZSnrRSHQj9Hv1dMO3SFDgqbMDNdVKee
WixEHuNGS/1BU78f27b3icSvpu2mldONJvRy/KiezJbIqhXaLB+sIh//ifxe+DSS
KhqkBG7dtDYq1foUvWEHY3wUHloVI5Bp5c24qwdei+/OS/3qcQXsbjzQfptUZQuV
1U61q9TdLwxYiUjB4zQ87IwQsB/84rNom9eTNPyOzXDUQWNvdB41VJMSyY7HtiR1
98gRWIoEZxNBL0QBCBmiMKA1nYNOOFAo+Rqu2gJWL0nRJ37xqIoYKj0/R2i3Tz4A
MXCiFnZsGci0y/XbrUZM2zmaeGQvs/TAC5fUWbmxDcxs9uzJI4FHabbXdyDdvqQ2
bGJRoEz5uA2cuw8fwSY7xH3sczx82+xMmR+v5yvPtFz02BMVWWuqx8R3P6/q4Fl8
y9xp2wSPxygvOJxS0f243JWlbLYr1L8VqXWlz1qmsXAY5bonX7lv/ztwdPLNz9nt
d/kQt0ku540CgbzUw3F6U4XzDmk51uLIH/vm3wfV79hqLHD2Ng4BPg/JPRVY3X6S
awOtiVG7ibJEEiprGaXqjFyXZlqGpV/9BuuYjKrtDD5MAAdcOvvAe60KmKW7KUx8
hYFjeyYFbrQCMRXRIsoY6j+frM+EXdvLbJHXDZZ/YO73Xg0Cp0pHWQR0wZPelGQA
tFMktUaD6QW3owdfu9UjIlc0p/6stWQVcBzuBmLhHbEPJZK+tuMIJR3oSXuKCTV8
xgKDumPBWQOUaPzKxOqsvPsDvUjjXEUvvRr3BrQKwa6j2zTIFMLpwC6LHDCAV3Aj
TpwcVtza6oO9KN8qTRlpyoDN2VMkhZaaK+NJ/nLXwxPmltoVOrghPxeEOcbXenPx
Eb16nPFI/sXgmzSrjBIb766Tkp3Fjg2aEvaUhfsSvY8H9rn2dy1tJj9Yu/wryv3j
zoNyNGZjhMKj/D1dNXldNVMhZYOV1qJ3UYxYeSSP9ysrd9IkIou4U538Ihgg4FwJ
DHk3HvOjB0Arjulo8fEpKK2lon3W7EAT2lAB1ikw/3v/XaMytK+sMfwyjmJkDU+E
5KhaMJiTt8aa7id2o31NK/W6pSwYMvT0xWtEX5J1T0Qr7qEim3Fr0MKUfoB6h3XZ
eXHiW2kg0ZNXcn3c8+YVcsDvcbqCOC0+0BFAAI08qHWPVadmVyy7H1R857zJ9fO5
56ndi1drYx0E6QYwUM7HWG0eD8lUb1FfqikzKvj3B/7+LLkKPpK4SrJp3y2q0oBq
chuXV0taKF2mhBlfPoGCypndO85lVknZCXpzmLnz3kRMm1CaU2LjeBP7C/AKBQQq
WtOsAMb0vM7e6ThmG7MYROlfVqrh8/UFQqSJY2JUW/jCNrYZcHs7egn3+8PcOpdT
sNZ20YZTOVLS18ZF6TmpmSchWcPnvVzlt9JwMsA6VzX1pfHBG3HXMrV1vt+sXWa8
0qQBr/EUPrvyhLXFf8oUJ5NAL/8HIpY3wdMnSMr+XWqfEyh/qG+SdS9miyeq74NV
LWJLnOrNz+JgCFE8Ex6vMIzItGV2TLfN4jLwkNtiOt6+1loxYL2jLr4oMaxdZFLA
AHosgXkP2yF5YGvQOtq186o6tvh3bcMEoMa4Ng731b3YHiu2DXgMJTM5ww+TRN5p
b5KK0nxBK1fKc77O8BhoN6o3dmVEAryPEcumflaTlr5sXkdfTbHs8Tql5gCuwMD5
xU4VTBd5teQZgIcR6m5Byojtcf//CD++05Bi1Gur1DKR6JpRKdyJ9Yz6jpBiPikn
ai/Bb0u+WUMTn7QL6E/NGqO1+clUP+QTaOSk8gG10I4pmuHJJHbuKYqNwQZb2ysU
grD5hLFAKM2iUr53BZ9kHJ7Ql90BbiHvUo19HDybFQFA/534guUS9YeP8yLfMlze
UG0gHzzelO+u1ISfjVPhyVGLxfHa3DI/Mm+ccUO2fpvMTmQ5zlX1HH2z8R0eR1Aw
3oC7Lis1AamxxuozXSTSBrAaoSGuYnlpEcg8bbn/hJwIsHSsPFCV1o6uavOQgSn+
V4An7qZ7HO2pHSCZNhiWYcLcQrxOA2K7LMIOXd1Ph/BXTstQY4nMNiObaI/Uxhzw
bwR3WJXQmrNVSdyjLlExv9QJrNiASfYuhEsrOkQy6nIIgqwGQRAd3lBY/UNK1q8C
VjT7iKtnXYSkTZIp9pMe57+Tfolq9O7ki1SCM5a9zmPsQexgrWGvJAjHOunDkO1u
cEwHLk1vJWNQf+lOS4A9+E2YHl4dDLmo8zCQEEgOrsPgabcFIJjbp4n8p2lE13LE
nULxgMgoc+rQz/0kxMkdyqc2/TTR13LZPfyPYb7lOrCMA7p6L78qUU0cmT7SyJx8
6G1j7+kQESziKYu5z7omSst+F47dG1Xt8+KYFzifz1oyBjny4I57T+4yKZ6KoBNV
TkMMbtFGDYoudhpEOeo922+GSEexSaQIthMWhEiT/xvA0eAqyW2nDQm5wgJbqbh7
xv0bxIrTc2IdWClfwOHrds3mBcQqBRCDkSL92RSMBrplexdH7zNPNqim9HiOyRyi
tcoSKzMt1g0HXD3khSXKM0mFbFtVXlm5tLdow9s0AllJ+HGsbSWRvO986J+BhMaK
ABkFYT0GJg6PvvGnXNt5+KbJca439Q/n14bErKe19fIoMr+uoX3XB4BedYWPn/50
TOW7pOl9ta0RjDDuEpkK5cxF8X2YzwVVojv+8EwwwPeJdHP9nRGgxC1nxoY6ftRH
H0lUdiUVQ+FxDmBn8ceUZklw3KKwvmYdBBVNF2frgTjCU9TLNqzM9jbm1/Vri8Qi
FBrOb6CkYzg+fHHll+yfYJc2oa1YxveGfNwcCARWO8h9H9ZwBwQ6AfL2ZF8GScbM
Dud6D2L0nklPDLSMVjJeffcL7Ly9DxrduniHEnFBLuLlwSqt50DCdYfMl5fVdFby
brNxCKgX2adndxPZFHaW2eEaWTMvNf9tJTLQK8Dq5JNz4QrrBsRvrWOlO2uF/VKJ
OI1/OnsqTuWZLsLerc9wYeTAvt1xlIGcwkE4+shAlIHN5TSM3cGdr4pCVWXbKXIy
5rTrk7waaOM7k5ibsVLCkXeaD84jY5G5/Chy4K9Wb12tYtSO6NN/8AF71eUrwiZf
zFfnwqZ+Q9W1Ni5yUqqLUVGSkKIxxiXJtRElBv0l4alUBPb9p6bKCtgtOcKHi9aA
7D7yfEyox0TWVm5Gd/0JA6cGagkN19qmI8DFQ9Ro5w78m4yKNS+xj73JV0OMx5IH
5mYhE4tUsq0OdF/JJWgkaAvbsnAUyaZ7CjbfE4FECIBNHvPdJYHhOhPPAyUV/s9e
qY+SGnZDML1P/TDUy6+Z7qAbHyzHkNCyqRZ5T0SGgFzHCju64pF1AOy1rSyE7k/l
LBfU36HFPbgcMzqGJsFfXGLBD7bQzR8qjPASbk+xvepMQeC6ApFrMLzV90zvuSXn
KAcDsTjL3uOf6xIv1aqlvZGTyhK/C7xHIeZZGFVA541Z4DnPDlS1p4gk+lxTF/wI
/uAySXbOsbVdlt/u+hp5e6XPP/s8PsYf/Wf7PmlQ2h6VZaxQetHqBqkR+2YkZsha
F8Ok6ObHEYLh6yX5y/myCvqkFo4GBXghBdwCil+dpBsCpRdwBEZhKPtX3hXL7xlE
WLg/fOyCC8WKI3j2jBUIVg70MDYCDrJ0NkV7hExBQflYYkSGxNjWmJREpGdyS25Y
obcrLW6EEJIUDrjpygGGjsur65zZ0NrwX7yR4YNz1d2C/EdidZv4Wlb9ECwaqDzK
m0UReeoQR+B4yXoCTjMOICdQsNu9IKs0RG4p4u+kjsmWoq2tx/8+6EOTkCE3Bryc
AKzWFUHZLq9XnHNsd2w6FiYYlJOZXxmgzwxFCRtwmz4ye5euKTZL7rqk0AXlIoJ7
87xuXjZZAiGFP8MaIZfudF4/n1eq0gvLq8DH6F/wof0HKQF+mDNBmjbIvFDBWTRQ
gGJ5reRMRzzMkGj8TFqBz1meYznGvJdY3auD/cICXRs0veTrixYnad5W05cMnB8i
A8lUeoyHT/u4j5QI1lkRcymjbLqthO9CSJR94omITXXTJgC7KXyMjfRnIT64cBhN
7l2wk4Zn3v+/ehYICj1oVJQ5bUQGJqy70eKZTu5grM5IPFcUWK0KVDihCXJXhYlT
DNHzBi97Cz1ahrhzWIW/W0DVpPp0rPVYcLrGiMt3BDNPcYRbK1HirOHVuptSWmQr
+xKVWrpI+CfZkDWN59AEJ8t6MCy9rGCJ0Q9HlRqKf2zFEPr6mMNM7a2nOZK3A0OT
d97NngTY7AAHaxrEeCTOsq4egOXmTftFGpN4Bta2OfV2mhOc8jDd2EmPV0o/s/3b
sT8M0W9O6RDTjXqph6YuEm6197HSZ4EPMLM+6t6Wp/E9waoN9VtWHwqAghkkIL26
ovRVpTtAAmfuZS9X8Md2a4tERHC+Sae9UtzZ0hQE/lInv4qnDyCheFeo77JxrSVQ
d2PYLct8YSOXxU0swjxcqDfcuMvkj4ynRkxibARe0mNEPI9aIeaG8SFrfe9jC777
00waP7FoPCdv2ScAKqZqSiN+OjeBoT+JHNV8yX5BEdMaXWAAIrw5MsaaN00bzGla
SWAhUNfuXsqUhMF5yoV1Sr4ZSzwwnjsfq2o3KWdxYAW2hXLHEw/XbCgWfh56QXYk
eNBsS9LJfmsdp5/XitfwrasU6xWmRunnxuYdw97ZUSNcK1q+W9H48w3At57tcr1Q
M9cweCmzsnukZ5AhHVK76L1QrW8mPhvplkHTS7K/w0cRcQtgq/oI81V23f0asj1V
QbOQv/KbA5+ubn2idU0fQj5sKwMsTC+OpH/BH9H00xaOHI4diBvfqqY3EU41ioWF
E5wOobk96pDWi1ozvzD6ss88Hk3NM4ewsM/A7o83TznyPmEaZEX6PXK0aYM/uDvf
l47OwFJCajUe3Y5A/7e4ETb/d8C6J6XpK+Lkd31Jh1rzm72ohoSKjB/9vVCR8dYf
ipi5RpiLNeP3s7WKt5QuZ3381TBsTSYcFwSBrCGAhVdak+BMoUImdmhY8Kg1ufeK
NKT4guF6zm6+g1ufyHB8dgQDSR1vkiKfOCyEbPgKgXMq0lpcAMyj65V2qbwMItTZ
lfYm/PbxuQC68acNcGFWzTZ+SPZzdeY9z52iOkG3sBwwcjlUHvE+ypjgCyDoRLMv
IW8bMy3zibUerYcU/21au+ibjCyze5RtrEKyQWNjniQMpZRxdW9UykpypiXjUtNh
llDmzp+FHWDLXDze238sHKKPL7Uoik74CIH1k2hDFnFCrZg/02jpMxDLffdkaLV0
W4attdW9rtWITQnBe2qpX7K+R5KUozG+q0KEz3rHdx74H4X9E6DjO6oDP0+iiZm7
0MePtWM5QjU2XXyMWX1cV953TA0s6ClcCqGoZ4G0Y1Hia7LjodYpaB03WUiC/05H
dGQ6cU/jNqnImGh6RC667xGbcQAYRRsaALRQR1d7PlSjrnwtbg7eASxRr+gaLPYn
2qTfCCLPnIScpHeV/c8jXXxV22R66cv3kpQv+/dyPoKzERParAuPYj7+58qjg7XN
Bn6+8uEPeUvrhw2atkberj8ArfVrArNYbYVpA9OfGXMnQ2TZcSkMWFFwy+JMbKeG
1ysO+TkBB63sl4qHcD09ZINnGmdLeHDSIadOsmk7/WVeRn7wAgQ6rBGbsGxJdMgY
T7veOdZLUtZ5MHENDKGtQ2vDP0p/afO/ZJlfrigkkoBLDgWpuyVccXAB+c5uN37T
XuahtYRIHPg3T7+IwLEOym42UIUBmASdal08U0DYveD8sQ6fxISrtm4TDdjEODOM
g9oo7anIM/zsgNcHbpvj8sRql59gABxgro6QzdE6mtsXkUrPPMva33iC9IuNfJrm
J+b6CUxcP+O987/r6T3HHSGxbQsUIZEXQePe1bhapRv1UynTxR2SVmNXPklmgZSq
MsHv0DsLadJBlfpMun1FfhpwRidQtRXWJ2A9iMDiC4eOZE9OTZWyYJ/JxEqf4DK3
FvOaY0zaz7fhl/560T5Jyu1H46ZWR/BobyD6o8tOT+30Z9GzR6cstRDbgt/Zei0O
ff/9v6XDfEOCIb0RVXYYsjqX2XWzWA5t8S2y9dkKJV9+sS7WqTr8dwKrICDjCkoS
r+b4dlMO0Uo3j1FieNm17Q+rnZGpfz/l5ANe1va4cMh/IrAGfshteYFW9vkA452h
ob2yVmpuDrcW0pCWPRJt7TAB4zaE8zRL/NiqTIkOar7oRPC20fbLqXXNR+46Dxy0
cwRL8XzL41EpvbGY4DK47pilr9BgMLdjAqpzFOhjDzLt2NAw3xtRt1QRkoanQq8/
TtRmFQ7SQX36Qf/z9p4Gerjbnf+Nl+TPLDXFEPvab4o0leBRlXUa6Z1W854lWNip
kDHurME4ZGpIaJfmcN+JEN96pTmmdp4q47Nng+xeYCCe3zSAz9T1/MNYJAF1xn/9
4kAnUR6m+JlvWSpQ+diAoShwL5p2/bMELiTcnQEeIcGP3am6TL5swQBirJ/nSjEY
JyfWefwgn/tQ2O+pq17byAYJPJqNZ9NaIe/ZpfD0b1agGdEPDJI+20AMjDoEYdNT
4f4HGS/vVTatMQLfVzenpX/HouJQgUyfG8WJjXe/7tuqdsUb3LGQ62HD5HdvMnrw
CasNjedJjPmChvA3XnQNSChLRzLK/f8qtV9dLdM+VK3jjfX2UJuR1JkZU8QZdOuS
Vc7Ekazu8W1zHDS0k5j/rpiO6RtaXU/br6RnSIesLaEVnoj2R/CfY1+9/uARXF9U
8Slwat8+fGCCa1Nodkd+O2KMSQ+q09KlZXklPQSS2bqe9Axrvc8c0bbeeRCo0DK8
rG1fdjcPiI4jrckEYnTCxUpJFFM66LdErOS3t53P0zBNHE+1agXs9lMxoBdASsAn
GttXw4CDctXGUE1UBgInLMnv5F7n4IhNA9tb0ln+NXs5AKeyk6bmfe2GRA9e/ABv
QGdag127pOcoJ8NuVPVfDafT/N4sllMC2AoMdm41BeSs5PcdZ4ykC8HaCTYLidKX
Mth53E1wG2fX+atuB3QrJP9enioey3dOLZFw8HeLRfwcSDWJoYmDB5YzZfFE1cSg
pAfcIPbaSJ8VLarD561V2gS+LA7A/NuvX50hOetstwqI/dnIbWul6visXOJR5hS5
sQFuJhVSCh8zbUozyTcTOyntxT0lPpkyfXMF/NQxFFs5bL0/LEOY9H6My7OeRU9Q
TY6NV2sovd2nnpRzt/MxdgHxG/0ITV6YG0AbEUSYp4IJ+4CbwHUGFGNae7tcDMYE
gaTj2k6gF52ofbSzJzhBhIRgjNFWnzFXiEIJ2dmiNBvZiJExPEd22mR2cnfjAu/q
SPbCoGSgqBZe19Z792Zof92h+iRy5nfYaMSV7XMYmsKvwWZY8Dzuh1amNt60MleR
eH/0p5rafA/nscKNndSYq3EmmmcUpHGM9QbXI2aowaFgXT7g6xTrEfQPspJSMmFZ
KiYYxVzC6mB48A/EG0a3LEvPdyJQ/b79Yp11wZkY1hu61sRx8ufsdBBbkEbY51n+
cALr54Qfz3QDtsQKwZU2zPwhXpvRgXGs7+wu1Ltdwgh+sJHOJBN216ZO5RwTTjTd
Mght42ESrkZhN9qbzE0ix9cCNNBKCYSjL366H8pZlb5LIBQkKHsc1nXI339zpWJu
CfKJ5LMUZgyaBvMXd2iWouDffJGp0Idbrf8HoyAzGi83Z4v8VII7OkVmySb1KJwR
Gi+MnPV99LN13KFWTX9Na6eBV0Uap1YKTLaieFhT4C+JeWXFYfZcLB59CLIk1UTo
JXrujliQgEh/2yMNmwa07LujNSddxmUsiisglIDKzQb6oMhUfMSWyZ2tNIbYfLpQ
DK0FacaGMdtTsgX5mP+92l7Za7BI5JgI6C5akMQm4Hh3xDUCfF3TjoIImgHHGIcZ
Vy4a2mTofzg5V4lPa5+2M4akYDXIiadoLsUMexK/nsmyV/7OZRiLpoBvscdGqIi1
AxjE70h3NAvTtq9HU9zaCZVnIGR63lIXqdhIyqkUMDNNETRfXc5q9uECEAfe+Red
j7BKYRzaC4HP+VY0soiXsl+DUbijglqOSYPrRo8u5X8h9REQafRu2UeEvHnJWe1B
0tt1ziyMc0khanOTdv9ajcT9YA2+ICvcBMx2Kc0RbCFSO5otS7o0VrVLsBxZSrE/
HhCWwZyvW46zLBv1tileyuAVaZ4w0JU1ZSvjf8mMbEEXZIBm96bohgnkTKuwUhe4
ZtE8slWZMPV13pCOMACelbUoP8M8AYJFvbUWy0Ui7zRFX+BivUpYwJeCeX9XyEsd
GpcyjwxCVKQvyzqGZ7tdUaCKzOyzWqgsS43aLKvbl2OlBeU80IZ2XsDRkIkvXhWm
rIREUXLkaXQFUsQtVDvD1oWDzRkhnpBJ0tI9zHxv7SJoHxC7Ew9yxsPQ/CQXoWC5
0tlHa5BuVhzQd89dsl2kxg/aUJVSCIIC9vqjBLIzBmHfcspbuG9Z7QiN/1zfwmpu
elIZ5i1Sfqi0e1LGXKpOm8WRm3La1mXDNYmm6TgmGi/ApTSmnPSqARoYKyYsH94x
NffvxYtTATNhkDQ8JZ6ElDdilifOBswzuLfGOvhY0VFZSkCiOjnFIzk3VEj6EoKq
Klk+PNMtsbJOoSKHr1MwLSwfQBAcavNTwG6z4YcUUXoIxlKCxZKg8wEajK2vYzLW
os4M/fNxPQqwJOWURbhzVXlOD1+9DeysdAhTzdpmaa8M0t77aYuGD3HKqT9JsenW
kmlZSx2m+MgShiTUT2PBV2Cp3GHtkRhW+nqp7QVVlG4zAFJc0Vzd442F6F3+9KDC
jva28nvZTj23uqxejbR/AJ4vjVBRdmKHEF7nWopj395IRmIlFaGvXL20kjea+JMP
k2KgQS8KgUEPVUPVLgXSAYJQbEOSbohgEtSyx3rQp1ZuCM/jp9KcuIY8SN6XBrkg
FtNvyCYP58a8gLRnntcORbo2Gyx7syPxkdl/w0HCA8RmRtFxd/5Z6KFL8auxFcH+
63h0p5RWjFmnBIZTgRgfRYKGqjpFl2IgcacNVRRrYm/71NYhbZWI5m/TiNnEKkbY
XiyWXvjCy4A5XkB44/zvDjOkAZSzFuTdfoh1QlvTDOenuErptOQBxhlFI31rwwEr
phDz52FHvdmKejZMAjndzuv1nhRi057YHdCbrbsGSOIXN5wSSmXw10VtkWMizv8B
eSiuntrpJslM8g5xjXsapxrOFPfowXD6CtWi8wCbjgdg/+CcKYB89ZB2ruhVs4CV
tPb5gEG3dzAY2QvWwJiUHHdM4vR6lML+VA02Me42E+R8URSZzRJyeD6Q+hbh0SQI
NzgY0GKmElaKqwrUBx/NgFBDGLaw049SFoQKylWsXX2v8Tbkc/2oxMI9dhXpljxI
iwaRru7FeWpeQwh9iDIw0KuNSNqYkOuHiuA4vWiTgj4qkj7LbpkDUUcAbMIUvzv/
uRBRjmCjc6IAk85HSwrPN4MtekyFDoZlFuTIu0Oau+7B2eVYPFbMHqFekhEwJK/C
2ZVFz+MbO0Nfi4u727Nu/gbf6SSQiMswrcN0qRgpbUNf+IWE+346vO2l/fh7VWd7
MjUqPJXunXe+DbztkPBzPxSheC5sC/pCPXleidMWcZ9+KsrRxTRdI1uc+EcjkMK4
wzLcQUAv4jCBDrSbwKKDlcVIUBfXyLe4+hzsYrkchMmJzcWwrU4BJXsKT179i25s
V0pYL3sEVDQgwTKJpj3vyT5oZyMysuKzGl38kEQ8nKtwiisxBwfUiCxsvvF3f/04
84q0zcJymnwVDdlsa8e0c/Nwjjylaa2eCzotFwJJV5j8Ulno56SaDaOgnKVFYvZg
gdzysy8+ySZKt3VqfQa6baR9dExOH3v7AoJ8+HqnYtIbn8OjzkOOL7F8MRSN5fdm
jOtVgQg7BbexHrTFD0m+cw3Aqlp2xGQEq5anjO3kHTNeTjbTaj+ddFe38g7ZGZYO
kDPjz6H3h4KzR25phUj9DzXa/7FppNSTOHVSMSmxb+mzL0gmwTxBX3zf1vwICYxW
plWg11/ouKjaePsbBBFZAHWzMKG2hZCUjORFheXyoS3iTTdJ+8DLsKvQ39zphC40
BDZ/Lg7Ft1tD3PIKDKSlTAlEwECzHgj9G3SIyWukh5affJgOMcszfFLzlEUdf8Ww
4wdsbt9ypPa+nJ0Eejmku+1WZjV6OqhO9T+gs+IpnigQ0oT9P+9kAL8iCT8rVkmZ
dhuYeBk5534R1OtENxwKJgABkXxltmjXVbdk2vaBTkCS7TFU9fPx2cukJYJHcjT1
lOQYBv4Bqy9CRBcGDv9Qxc+EH7Uf3IY6y0PxTRkcRhROJTTaiwGK4A5gttmF1tIO
sU26ys7VhxbLqMkmamuJbA+gZibW3Unl+8tnDqby1XzS7YfXxDUYYyLSV3VaWJzN
1Hr3F6GSt++jtFOKxk1OmPSyGV6bJzcwrnGbmfYit6p9D9BQCX8H7fIsRX1SBhcX
SZdSe+I1GZG3/9EIkhPcWN4/gwRkeNwOa48xoBX3B24C9LnZ2nKvEKRAhOE8/yWG
pCpDPcRiejXDELVBrmBTnp6rZ8sa5lfwNqV0PBNR7eJzfSsTopt14kLY2CK9d36x
olbOFjZ0lHhUwuV/eOqfdVw5FlaoxmZcrKhUDfcTpWGLMydyrzhSpqLP8JwnJYIh
e7yI5Q9I6O+jnVpc8413nXMES4/m+FenDt6qMUAJV0O1KIeSNT7+8GySgaA6Zc87
pAT4sWU/5u4J0IE7E1cOcc+Rc+s9zXMkX+RdICqEYW8vBXyDPAEAHOJWH3INhZ2T
FomSesB80RvWvyzBticFcph1RFGTIoZupLrRLc1DVaGpN1GyxGtkHNmVigynyxKH
rTFAUKHQtnrluZAI8a6+r8ThihSyHQJnO5Jcb9ebd+pBlFeIpYkOjpnPCiLP6Zkt
+OfIciW9QbXzb54uv9TmnZ/8pAkDy3TaWzmVTYO/QqtnGWbkoCDdB5GrfxNHSToi
XMtyR8+ZeCMJBur3wl76hgI4jtwSaf27/mgs+WCqF0bo7kJjqOgrSlaZgEpbA3bH
C5Aghn3mDaf48drG+a7LAQSVkoULiAb5phnkvpJOKsmVVtwamCBUQWbhB3wISKyz
5JP4ATtHaW+Y4gg6SH7s3vea7g4KQkUuNRbnzD86o7sDecQY8QpDpOUQLY3QprsP
QK9CyBn+p+BrlkowF55RwQLDUmNDMeqx7XZs+tBxmUjmM5pDj+oPRr8LW7/y3BkD
UduWvhSWGMQDPWHstOlXtJ1eFtghRnSa7p2l/4KTIDXi9I8HvB2rLcnSlBkxQkr+
WgQqnbRIVjrjngzD2kkXvLOxibAJRRGltCPYNVmDO/Y4ro8FYzOITG0AGAvMTtWk
NXnByoa1dwqzGKVQPFWhvvaAaKnQfASVtAtOM6EK1a7YYPIyX83y2CJV7SZm2hqz
pLHD4T1f0+NX3AZ+r9QMPQ84nKCHCfKdnJw26Mr+srs+nvqIgXpSgVKsWICXUVfy
WNWfspPhaFrXQs6PKa++cpkDUzLvZufeBr7kLd0+KLv18ts3hY7B8glAOg3L5MvE
nOXhRetUr8IWYsUrTCwgV2p9ROuxXiOqKuLa1EtC9g3cFYIa5aPZA67h0nN4oUAk
NWvrrHm49ePkaa7m+ufPC6HKPfhJIiMyy8U3/L/yS7CDRIAqV7mCgTBNj6VIJ/uC
V8G6KxZd6hxUNu4ZA8KYw5F2ZvHw2nSU/1irc9Ma51noq3dG3inCNwYP0fn8pjxm
GakNqMRaCL6UOF6lg8ZwVaQBLriWOh1QyBHUbzEEXjDdMRMAqiTuiOh2NvJL/lh4
2+F9+JzJo2MMcYbsAjxcqOvCMQTpxu3CkqHbSnpbZ6swYstxRwLEvVKl+PIlF0yG
Nz77VCD7QzA14BJJrCCMRBhd94lVh/r1J8UAk8d15/vQKsNmOg4wuNbgLOmENGCD
IaI7slcROwpaqbxhs8awAcIxiUcCGvuGHjaxoeEpkxyTyU+OEeI0FV2TdNjPzvGj
cvrH/abmAhlBBG0cjlsKLhITEDu0QFJuoNKcf+Ho5Y21WfpyKKcTlVc1bffVOwEV
/wCsZ2hN+sIW9skYoF2JmEm9ikeAWzXPbdiwymRSRX+iEiDpw/uGU3E22rTPmmcP
gRe4hFskmpagz/grEiBeyFWhFlTyAlECPc0FxQ7jdUE349ITXBeU0jOji3EWXkSY
6vfGh8RpOQgW027ZCFiPhUpJpdNZ0ctxHnrELj1OwA85YYe0E/8iLKsp5FYysH3R
pN2qO1XBR0jwv02ITY4sO824dmR06vN4TyUORN+SPVA22Bz7nsvmn766FuNkGBrp
1jy+6c62NT+TYg3LkKndgJXD+9Mh02Cqa9J+/3A/8SVv78n70QwnejD6hsK0i9un
tubY93q49ig6Wlf/tsid5Ebc/29Dw3AdOA8XMK3vClSpy690YjTxkTzAVL6PYUmC
/U4QkLtfDd6S/WDRZ8OGc3JizWcyjhO5GdaX55jfM3OV47xdBz5phSRXLi2c9QA8
piyWJht8CfbzX8EIHZr8UrOXzfvha2iSAnOI+O5cD1aUnMDQX4VGBBoy6K7Y5beB
WUZVsRr5JxbHjfOZKhGodvZYvF3VxNlMnQVDpWPBwedzf7Hz4tyB82jAH4pqPAHm
WfxYddB2oN+G1OuYA3uWL9mLE5l0s2sPvp6tW7ZnYCMdqQpSYtwpYKzV8vAShWQN
M6dHs/nTJwhAQhI5mBjRl7CMJSVACQJx2BHtb4/PuWSDwqRa9hmHxtolUpfB5PtR
2fnnanVbFKYrhLHZPU6hEwM101JkeEtJMkBjTWKFIy6+ig0R5TfRh4GjoYIXbfZV
sjD1fUHMtrljTPK4Tk0UqV3ROkniM45SE1MUT0TeDT5rfz6o+1gxmONZBj6X2Qe6
gsvxKhA0yM74F5k06ZMxeFTBuR4kk+NQS1tInO0wO/Dho+y2eYK9VrLEmh8ECPPI
GYSsi/FMxpuDL4q/TYieIQNDbbTWOBngvBrLmfx/qQrAifIliFLBVfFAhOy8qTgw
Su+EJs5jfX5eoAipaqbDLXOkoxnGT1By07ewh7qM2PhojsdurzIvIW8OiGTUdL8X
y5drZe2atPR1NumnAQUw7F4xZjfENENTodNhYlq5gZ0Of+VzFDm5Cp5xNsutx34d
t/Ijct3crbZX8Cz+1QxOvtD5yCRuZ9iMqYwFsGe+Xg91Aa9IrgvLDb5yJcuT/oqk
oztP15nXuBYQRSKWYfllq2jkfiH2kPpJHyc8SQdDOoFVFvo/Z41bv89AiB50MM57
sKSBKQHe316fea8vsReWj7SLcZePIbQbOTKnoPXWvHv9vZhpcT8cWi6HWGFGaFhe
fr3/IQdwWOylJc+qTnKVpwN/LgkAVAmv1cnupkKxenXUrloFfe68QD8ehZApx54E
W32AH5V+PnSs7Ry74uQiQQZq3vtGiS80q/Dx0J9dI8QnlPtxAf6s05YCLDhURlW0
1fLrXVql6nLtIJWA/ite5urAj9HG4CcJF5WKY0sEF48CBzc9vbcFnnYALOGw+Pre
EaGVGdfNmLZPVbK8GeCzalkXITkgAOjA7otqoMkiULkQ+HcC7b1mB0QDLPLBfryb
dpBTdc6F+zRq0krciTS50SSiZs3vf17hdPQCPDvWQBn5RwipiVul92gQ6cxC/Kki
/a6NlUR+QoH/KhgqNHEEVFB0goL89juG9vP58KFa9SmYs3YLkebQDCwdSmoN7Blx
rt/y8c4c+fhtIBDVq3GAtxyS3oaCgRzkQl4xT6Nb1+6w1IznXvXylivVi+Wdaupk
hQlNji3zObMuiWsqc6xbNGDtXxScbkUkgiXWtjYKIDFuml0atVpoHMjafRZ48pmb
F6MwvJe7ezvRBsk0n8k/H5GRvxcMWy9/EjxeWYObSx1OBDjo1/6B87Lksy5WSBn3
JZo2tYqNv4qM9cISl3jlJ6XMXoG2kq8k9hzPk5bWO9l2sLTsGBqF/zAY1n1AtZpG
M6QPOGsYsQDwQ+ic41oV5fCuaj1FtST3XvQOIdoIG/OyPnPuAXzwYM1EbKhaDmcR
VDNyAmEJOyxW7g7eTW3Oq5iPWNwdZpNGa8J/TGfN2yuhoP7LPmD4swKYik37+OfQ
jrqiNMsBgj7uWuKdc1CQoj7S6uWeYD1mHcb2DyE4U9iijUoXLzrnf0h1/ps+rv3+
X7yMGZIDsbsfkoMRkg4tsmLQmJ3qmppgG1YKhTO5BGzwRv+2/holxOD1DHrZrhC9
/NIbYY5bqjPqWD4hCeYCt5xiwzWwLShoReEwUFVuUy+htz72kjTv0ba+CBrSQ4mc
arljkjQCxTocie+lFxA3ohfysFEVjcja0448p7lhCRbWB/j95u5Z/qq0XRCovMH8
gYuYIqHQMH//8TbV95+py77HKdJcRp5D6RPVOt+HbwzRw9fatvl26djMXlFULSGS
+4GiFrAUQ/KXTf/hWTmfOmFh6ujLpfKAlZQQM6aMx3hy8z2C8rng2CNXAp0n5vxy
Yb+0BH+/14PPjZ3eeDb9DzMebZ+zD7t3rzgjUtX2CEoNyeqQoJAkbA0EzIGyq5hR
mr14PY+rrC6FmULNt5bJhILWXr3GSw88Lbavhppkjdy/0PgkbqjDul4kt4ujpaOm
LX19Z7Xuf0bG3jHQuo5OyZLiy3swuG5n4yvvKvHI6sOAptzpBDjUlR5xPm40trbC
SnF2wGqmx1LtRkP/+hBoHhmlvT02MLe/v5ihxExEMSEiOJgZ8H5LILUS0UKevtg/
jeaPpvmQbF4oyyjFHWteuKAj3hRHL3CPEzljYWrSQGvLYS/GXPFC9YwzXIhyj/TK
hE57AVepvW1dM21am0JzfUMJA9zAcwwLIZcXsQ5hkc06rrmDvDkmJViKtls/cWgX
vEbSj3J0TzUygzHjT/dJ3PUR7YbV4OOhUZE2v/hcsXGpoK15HoW2h21k4tB8oDrM
snxCL9a5GxXStAredKrGYIvtyxB157uA/D7w0yZLa/NtTfjsjscftRJ3mKlM6hEE
HLm2K2V9Qhs3ve0Ig49k0zEovuX4NPijIgXwLA9BE0T3hwDkxtG+HalE9BdQwzSX
aNqQYkaP2IAGkdqtI3sTHloyLJac8pUodVwUvNNnKa07FTM9eV+PD6M0ilZ2jXT2
4VzjH06MZEhHT5PgceIPBIbJRsHkJjZmL229R+RMJ0C054z+vUFmRW4olsQEBkHc
Fvi5r5bocJ58UDTws8ZjzJkD+IvYMUcU9PfyWPwgRuZ+inkUnCbRt5eyHH0XOLI0
AauulW/P9/o+uo+fVsVPbkKEi6EQoD9YRp1i1jcLTbQLVFnSjmq7cqQ0Je/Ud+Od
6j9oHlyDWWBRdBRPwmn/c3m2ToXxCmAZv+yr9VUMvg/sC3FWgkZeyMLNbbDopvoq
u5oUGDr1cvFLV4OSxCaj27DxWw+aShj6u3weURWZxtBm4PRhEfTcdNrqFqDT4oeB
mQeADd6SPgp6DUV/EHW+GsRbfnMylu0BxLRIWp95eZe7oB+huzw77QGkh0THab1B
b5YeSZmmJZG8joTpYfreEEtnU0mwxDAr8YDaYa0vgONuyHJVgJXsrvBKYUuziItT
AXd7a8kAbTLSmZ6fTi3f41fz8OudQ0CXItj+ayZpkC0xPW5NMgxqp8hiusrJD3D/
46lQJgUWMvneGiqbiaIf4OvAs3Xh0W+XyNmwJFqiXWaK4ve8LOVRNZ6GLUvOF9mY
gb3usKUO0cgt4Bsg5tmYmjW8MOj3z9qqzzHV/cDenwsVdai1ImRc7EcDqKR48Ps7
aK8zTrnbs10Tg5Xf1WTIIbvY2iHrDmOV4rWb74qQugXm3qmsg9zl5XHhP2L584vg
CA47lO1R7MEtdIsKJUNKf44C/BEvbRxai3Q2MWFQweEn31NrZEcfOIMcCtRdbjOL
wMRJVOUAxpBmKn/jDX9qs51WD+3JdM2D7KXLNv2MjGyUuEhd0bDV1g71rFWqigoU
uhQh/yg53dMg+JaSueOoLuylJBVqaCwc0cYSyy2Hgc2X7m5yt8Pk0jZiNFzvpZth
7x9LTmNE2EE8UAJpwI62xVxkmRsU+PvBTWeHU3euNaVrmB7Do4GnKepm2mE0pPK4
8j0uTd1KDb7JUlN4n/Qef2tdC/FlVHYxvhoQkfYVwyZ6pyPbjerHMuNons0vXvg1
sChwXd3RSveQfK6cwe8xHECt5C+Gxh5jsd+MfQUCvlTWiRAC62/yI1VAnrTQiPjT
vnuZQtKbDnZIasgtk5i34xe6gdAk+bbmHZBuQRZ/hyW5DvpBPLqz4IS/I4VaGBWQ
rTm3L8Qbeudy401FK2qT+Q0OBhLof7t5k81ppudurg1QvkntDOiqhjucBsUGEx3n
b2NTLKgYLQAGUy71M64srqyNRBB+HCfuBCgN8iKQ4BauDQHzfOYgGA5Ro4CHnTZA
OCDHAuluwmh2z87NeDdqgzDaTEA5tOfOY1Sg/fzia4yL3PD2B+j3i3iJF+5yQDZF
hLpeXPD+2WrqroDtSGJNMpMqGlUJutKv0rxy5FAY3gTLYRqoM0T3xinM3lFke+XY
nQzgkDU7SMDmZdFTnMO6DZ3pKIYsGyIrupGZCm9a6HZEO+JWyyMJiscgpCORA6QG
aQ3oxl7dtagprPxHb/bOqML+INheaJsENXlXRep2PRjCyyz4mV1DWbI3SJEe9uKQ
xQkfi9HSqQ9umjz3wZrZYz3sDSZzf6FjcKgSgtqOh0XwSG84H+yaO1DFQC5gdBeY
w4NKHTUgVMqen0Gnv5ZfKKTfx+VfhZgFhgYUT60MguMiChqNaDCmsyzKmopU/sx3
UKY1HmDQzWhAWWW7U1i+iybcEkUyDc3TIkd5uh65gXIOQUueHYwd1A8YhIMEHAXf
1F7PNiu7ZcEel3a+c2ddC2m4ZOlYLvXKf92rD+WQlgLHRiaqsuc6ksPtMn05gkpE
UFZt3Z9HQ4/efhIC00wOqpLgocc0YMrm068HeRavHbIw6n3XCEYxkJCi+YW8gND1
I6p1dCsfQMh/put7+//xv6mk+uJ5YZ4R5E0I/4twOiNJQMF5cowgtcyPsQXgKyDu
ziC47289OcmCk/EFtOgl4mfntvMBYLGsmf0V7UpTbbFp9TafwY8Yd14uUk0yfyVj
fr0/b6W+PkvJeXWzpY7rrhAEpa8iDGNSjvy95HKZdN95xlqlmDHMWXQDh+Xfl/0i
Wt7ZaAXc+ZOgPmAxqic7kRk+Pvs7xDQVQbDrz1DHafaKpUjJ+uo4JYGv43B1j64s
qLcYywn4vKM5DC91rFDNHE6665njmGJ0XmB9xGGV0nqsEBDpScRUjHfgTe9oyEAs
vqCY8G2BhKK8LnJLPN0URCUW0/67J93HtUoV7DSt6A0Q5YzgldFCuxc9MMWtb7hy
8cg5X0l4AZ80tBMm/+N5Mck9A5gZVKuv1HnsKKCR6F/3Hi4tZlVYqD5ceQ6+hFwI
CWL07H8TUeBuvoZd9t/x4cevOYle7dbg8ncjhx6uVUDPNVA3plQ79WnWP06p+WNe
rxD15e4N5sXKzArPZACKnFrM5whK8JCwRMtqIW+4FpIJ76x5Uwi0EcCBQsMnxZjO
bl9YZb7/24PDHkYvmkMusFi7Bwa9r3tpMY+okeO0XJIxG9dGA5j7xzhuOvsV6Yud
brsBiXX2PcNZX6v1eMaA4H715cerZgpLvuMM/9wmcnPSmlZbdYBNF7e3aEe44qOR
ob2IfnFfvnXbR6/2XtF4NPf4D/ZNagOPZoSPLAWLb+BFdSjTraBb45yvLmBnd+Vp
2gtdz4fjq1TLdGtJ6QvRlzwiGI/BGZcrHtieBZQ4vNBKsvX9OWJC6M/bE7+/R6sK
NrtrG+7URZu72mLuwVIxms0RMffXRT5A4h6phvDZWRxCceWo6lUSiR0mollyJYoq
PPPuG69EEF8EnbQRhlq7h6eNHMGHm40nfgr65+QbmfSBF0RuqUPRuXOl4kGzVNaE
5GyWf4urp2VAsT+TAjVszRV+Mfk7kNk8TiZQH6j5ry/IAGb6DpmwkE7CuCgOvRBV
kvOWh9nfHPJoHz2kAMfnrpMHyHCcMH9/vBlGtERlNKpyOsJ6BsU2loJijjnQr0OM
t3wP4ixdFT9Z3siWsodsdD2JAQG/HFnZLxss2qmB1w8wn4gEFIxfFlxC6R71K0Di
X8lz6jJryE5E5wEyjFY6Vr3KjXk2nPelyiO6F9zSPHvazDI3VVt2YSEfyIKr8ZUb
cgREEfc1L66UEFFjEWSuXHeHJhy9o7aEkIqqwXY/FNFh/PxfF0FekFDNZCmUWFLA
sgrmpJbdHn/JcGXP0he1qafzVt/VFcE3TQsquiKNxUfAxGR4kqV3ZqBsnPl9dDUv
yPjm6N+qH02P+2rrG57J/UtuAPgzX6nlsjwGOw+gq0ZLzAQdv7wwQMOLtUCE+e7Y
GVKrfJ88JirCHP+eSW0Cpnxxqmy2tV9szz1soUC9kMySlhfdhT1zf3matSeiwdPg
WRY+vDanihD6GuDL0h0j4aDBX9EY4LaRVuhnva9j2ns/yLmifbWDJrFUyOBKb0n8
kQk5HPmDwoFVne9PqTPwo6NRebJJytKIJWlTFwtmT+7w54kdkaGP47FRPmjIx1UE
9AnO5rlnJsGLYaaxvRu4huZCx1S5AGcvlqdwBaresusaX8qsheyfG5sTSz72BtAH
N5VEDQjuZ2qa1oYr86l/foz0MPLQ3v/wD5exyn4FnaanhFEin4g2V1hnIpJ6vWsD
3AERwo4BXshM1rNEIuYs2hWErEdQKA1Z5Ae9M0Xhi/FOX8jZR9GG1n1oYTCavLpQ
E38firKmgCoYjWDat0jT7I2zNiXoaEfqhfPu5yhfwYNeDRH4gCwn5qqgyJkj1j6U
/YYCFDQISN8XhqR6c2TOJIAMrD2Yy8rgbsuIVL2CusnURvbRx+36zcjAYMY13yHa
ju4PksAfw1QBzZSeRcTh9ImAgSYwtuojkpLnBj66DVQe4E7wsL+pr3T2NIjjg+GA
sDrJsAOSG4GbelkwQdhkv3um6NdDxJHMpQiLo+MOG/n0RARjwX/f96PDZeh4lbzG
pptxe/KbeD9Wz7MasRnK50sGaWb808gp738ZjnX4/vHzZpmNpghJsSBzQgAtrkCR
TuYF7x093amgJbYcsh1QPaUXVFbKvX3Re2BoaVcvhmc+dyF4z3KyrDKgo43ET7EH
ccuKhJgxLh3pNdwUltvuc9Gv+BlaCvxkiCp72S7soPUqaGago4AmDYAkhrILeSu0
oKuzJgZpilwblaeyZ5yZa8FtGZq9S5cP8qgDBxphSGjapk3cTcG80PqRlMLrWbiH
AbcXQVCyw8mC2kCu8FHtdJGiED5bzehjBrNllXkXhHMS48aSrLX1R05MmvYL9sRt
i7H2DvQVCDdToMV0FC4gECW/9fydp4anSianxOI/923bpRBR+JmRfAePP1yhqr2C
qu4eH5hRjt1ZxF01sMiicMwWeLTddx2plG9NlRz/nguS40+cix6biM6lFybwynBf
NtZB5A0xYTuhauqTMGPHfMhE9R+TfBijbzv3JKLCmMNc+LCJZI9qcY0FN6bHSimM
6Anggp9pSfglMWq06FR9h2v8jombKlMot0oX5ydO3Neb9xWDoi3z+gw81UjjlmYU
R3ayREwwBcL/7hVzeZVNPGaPVCp9BXehgbXHFo4Biuy7NztO11tAzkYW0ZAuMFmJ
e1MjM0vfAND8Llr98x8toE9+Yw7oI5O3LMGgLWoV+RkPeOeLC2NXEeKdtnOOO7Xw
50uQGvu28u7cXlzeOTPdiREDRUmwW0wJtc6UJVLQRu1LhLEFAc0uQIOGvJ6XoYpC
kjv0cjCOCLIthNLx4ZX0YLv+isn/UcRPYkN262bvohf9B5ssAij6VvyVesBBXR7o
L8Fi7lhMZTocfQXWxs1LwVH77f+E9BboUpQgYZsotBku/mvtom/dtx6OlzSivGDs
gTfSj9O6nWcsKOjfLqOmzLC2GwEWvZq75Ch7PeeoKcI0la3tP6BDF8/ZaEUktxyT
YnsmJC8fjvVtfRD32bwslvSWSpcyYq2OMsSzSnIvjOxY6VsaF6SkUQ+WEHjRlW83
TUatsC1qk143hZ8H014xBjOwDn0/jbBTI1DN9raLPrH0SVgjpvW3bOLO7BNbJjam
FtPo5JBylAT9xxNZL+h0Li4OICt+vWGQzl+AOt1S/xq1sbPMuKAnAEAFWpjTO9Rx
me35Gl8Q4v/crRLu0hmQsL0pMAJOFghvn28rulvGCmRbvmWkBssCRiVyBvIJjO6f
lXMm3nyBQWahcf46+UXq61X4WwBjTObXrJmTBEQE5GUPQLeMuvIlLZgAXUR9DWCB
dAGQ/HFxTtCp9Un6/ogGW4DwY1nwNvEbarLJy7FV9CLC+j27erjFPuWbKLhYjRSz
7NCf5c7i6vhGOFEtG86PmbaT/0HeQeRAv3fwSM/W861kcZ86/QRooUCVPDk4U5Sm
hPF58uLlEF32szBair3SOmSyylHs6lsNvsc2VX3Xd9RVp3EssGDaCKWckb3fOvm2
cvH67OkP9oneyFmMP8s7OBMngAli1oou9jiluH1BcntsmNGghc6K6Oq8z4L76OLX
liNMk/0/AlDPVV4UAIGm9Gh9HpSCKiif1XR1bXhHRix2YNZ8blTT4vc0SFtKD1rk
AWIyEvrXxRJdC3u6SyA91LOvJ7Q4yJfLx5OmAwnbe/NIFUqQ28s4YfQxHTyM5mgh
kCow3PPrK0hTolGHukbvSDzXMDElx8Z7IGrK32GkYL9w/EcYo7i46ex8TuEeKgXJ
LE5yTEqRmjq3d66ecLbHX1KObh9pfI1VFkRfn7zz6aveW1Jw0oJ0hUNUi+aTI9HP
Z31M5VQEwQRE71HHaQ+txX3wGooJkfV85SAmlIqGhT0Gk5WgrS3DDc4/Zzf31MXG
VaX/YqNsQA9xA2OQpEU2eD97idpXRkI+9sqbxXTSekiTW3VnD04UUmH9aN+io6Sy
aaZ+ABoZ0ZCVIyDF1z4nJc8HCB4eVrOk6bhTWsSi7+DrQfrkLpVNhNgan2ubbhjY
D4TK2tUJpFw1j8/6KEhJwurSPuQpEIid5TVLdJ5uNHIxAUW7t8UJ6KI7UjBmMiFT
9PRJgBipoPPp4w/zxO6qvyp/C701A2+3hzMvZ/ILxV1XTkqBEQ91Q1riTrxS/MU5
fbtxr3bWBD6QP2vRAZRCywkFmxTIq4je7tZlu4hun8zsbMgyeId4LhwKOsZus+pi
UZ5gc0pyDawGTB9B+37y3I/4sv2poXC03iGGFbJ5qa9QWqqVez5JeETOksf7cipY
//V+eLCcqJuNNg4ItDHKvEpK4HEg6+ORX7ZlThotO9vvqBLobLGMlcVCwyNvnpOV
EubqyriX9OfuzVrf8HAM6beSIpVXdR3zdDuhPiMCrAGpQ+RkFHe9qWWkzkI3Ut9n
hzjJeyuQb4a1imYOQaDG6YO6xmc7VBTxQMCZWYR3LLN2t8BnRBBMtgf1e5deP563
3L/UpaQiKnRNH6Jd0zzqeBvo/YVbFNBdGwgIMOCO8lyVyhjKkVyVWAmuUv0LaziN
VFGbjTZBTejiFljAhZRaFnS4d7IQzUT4Z6/oFpgVNWmILbMXtAF0L/Po/0jvmcyU
aQH1Ij8m7I1J3ULa2jEmHwmiGLH+FywP1TPTqMnGWPg1T/I6suNtyiNnvGwZ100f
eCyRGgDt2Kc4FAScRYQNe0TpTOeGfUMMl0g92fdYJ2Q8z4qNokj/XTROCKys2+7X
OnfvJ3xVdl/JT+XhCqxMIqaDcb6+HwpLcGKS0jHBgvEtuSW71loZ/JzyQy2VdZFP
RcRiybpqIPsdeCSHt1SkhweLHt2DcyGldJvuHLSpAceyQaID4HCbJ5bxtOu0pMLU
xzj6oqBznRuxwsZxzeEiM4XIlmiFxkkmXXQus/t4Loklxui73KI8wU2dm9cLsJC8
AfiiTFPqaHgqEcNUKUjTdnGMMdQjvK8X7GYuA6jUR+93MvQWljUSZMBf0Ame+5ln
JzvhFqDVgeqkrbmM9NHw7IQpQhvY6stqqPe7dUMxI5u6hgRrDpP4YOlNF3UkMklu
PQYNc3DXujqwOrKRK69k8WWnGCi6OHhXRu2V5+sUC39W7m9Co0s/7NmDpdsBBKSu
4+O8nPWbeYRY3hqj66SJlCqrrZz3x9V48hs1YX2YyPNQ4Lq8IiezYmK8QDXlP0u2
MbZUa2pR8Aror+2lzAuMSyUNWsw3axjZfOmROAOMIDSriMQZXHIyeQtvsiwO850e
hnwfo/lIuHvGy//IgBhsejk+huD2Sx+BpWz7vBM/SzhO73rwKM9FIIoC2Iih/6OW
Bfmc3yFe9VKUaOvBaqRhCIVotd9bSENRFv2V3tXMp0IID9o9JN5y0Y/H6mg1AXBb
6+7KYgD+NTkoKhwBBqiBa5VVvRH4vxeSx/PB382ZZjFUVsLEf8vZugnwIVfNQPmr
ajakTTb6hO4DvNKd/wNJeg6ydSnfkOzqRUiuFagul+U/e6e2qENoVG5iFfQ/zs/l
D04AVlVEAoPl/x4/3I+1YvJ5VZ5kt4CufX9RbEUMTNFymWp7ojx6APJFiuLKgL3B
7bQPizkUQpxG+jmAph94pkY74FfeqrlOebh3J2ZPh6dVkayJ+tIPqIiJt1dnKH3v
rIjUPSOK+Z9VLLRCi106ff3BlnJXUrVGC+Xc6SFVK2QD+wKfQVj4UGMLDJMM/6+6
7V/Goyt0mbacpN/bWWLGkEdsjd22dFeXw10sYro5rg57UE/TpBsy1IS1ziU4y6Y7
cWJ5hyGjdHDwDjUGTs+YzGm2z1TIXbHnayofDr53tBSK4C6Bv/Hn9cc4qiyooR31
qGiCKqck3l1EEy5ZcAB8KseMlzijwPZr4VnASFhnreYQFPmhpkGK0Zolyzm+GtWZ
uQYovNsJySjawboxrmbLGxLDcFaVVpsLm1cgVKyD/FWzjtc0TJBUzJkXOypbARq6
bdcUGPceyPZNwvtoXEYfPRvoAtaFJkunRa5127LFutkI6lwE+FUrypyGgOqFE7CR
NqbiZmVfM31yfN4GCp85Dp92l/cdWD1QZ8n6Sr+w5dgT87o4rFSmJcWW3K22cLJG
2aUXZFwykwTa8u4oy7WKL82GWz//FADjXtW7We5/6g2ONtiMnbasQeXWkKWbisNe
y8+CXY4Zf51+55zkf74uD4mqAZ0nvSaVXpm0ErS9va9+6oFAHo2Nrqb5mMEcSfJQ
lD7G5fCGp+58dmHc3QsqmM2FFkl+G5b/PcTXFekjN/0nr1SkQkn7nI3i/DbjBsx2
MOMzNgwSxxNnSwrfEnStP37dk6KlYFoGaCx2C+mbFrjm56LSnOq4LokcB1HIIIbZ
fBst6OGtGImtY6TJA+LKgn1vIw0ph31DWnt99wymeB6wZblrWOAMhPLCS5KqZ9l0
UUIG3vtGhwgupRhQB9I0ycrHUrqs2vGGvTHHmwPqcSw9wiwmuaAFka2N5g8ZtRJ3
SNG2rwWvS27hVWAy/nLUALcfRa0xg/FK1TNfvXRwKBw4RtuOBzc/YJPQ1nIVx3bo
NAeyJi9NA0/wmaoFttdUnfJZpGX6bVaKW9vUqxhIfHFoVqd7ogWXf9Z3Sb3+TD78
zsRoobeLHj5BbEkv5nNautXQa7R8zCefMbvLbUum6/Qyvj/LVdExjaWw5hDLhiEj
bi77mhYzbYWSOeksiolV9irDqSklA9ZB1kyxDuRW6yG7FNfLnYGei6TcRZT9RAmJ
2/WfsIdY0ZHyyn73IwIeDPpqE8S4j9zxWYV40w5mXQGxXt8Leb/ZaMTGmR64v7eT
zFnTeBqkW3m4xEbpTfHzqo3Sqy8aAistbngZAjtIT/J3C7ea7xF6GQY4X2Uv6ojj
FNX+j6+9QgCZ9Z4lsI4quVAQgIgF+Ruv8WqhUs4cheZJgOnycnkYZYZNM6R8+ZLk
oCSnZk0bWYvcsbqKYNQb5TTgv3tmgCLXm50eRi2z0d1eSocvfli9cpcsMSJgvnl5
jvhswp/AhM98oKfHDN0qhdc0ppN1BomPEtc9IGHyjsS2Wm1QnsvKKmkQKNVkHwPE
ul9bdy5obOYFDz5QuduI5CRScDIk63jez0eH4uUyjiDoSW6SmSoQ/F/O9C9X5Zlf
2N0SgU4oMI5714LqKcFoa0gsCOu1i7NxSCC2MPf00Vpe2kIFhRsG1vwQSS215YYh
gP5+xukU3wgTc9AUIHa974GG73sBs9J52UrCbT5SStXh4WmXrMwLe9IFZEpRvnAk
eNfZ/wPtA2TbZ0ScrpTodNkNRpJEEmTWsWb0s8mDd1fTMKf19Zcfyg/Tzag7nP5W
5+kWp/xdUbwEfOC1V2C00EX5QUNP3ij6lVc2HuOo0M3Lk3SNJHK7bwThWgykD1jP
ltPhRgr8/cJogVbGh0lSN+WYlE2pBE4rpETwRmdji2gdUZYFbQ/YaRy9p8PZGIuu
VWVf80Ca8LnfYFQKhLGi7Dyerc16oZgjbobwb3jEazhNEkTLywck5HChT/f2/Mqe
ZK731bl9O7qHPBOX0efIL2ECPh3sgvWzb63/Zr6Oiw69nLAaJnEQBpw4BkXOun0y
rdqsk2fxngU/LudSQ1xRUwfMq7X+UqtmGWfEksZ5HLARiP3E5r/4uERecxGCLljQ
K7TaezRsnHlaCVVhnbqRxD7PLg949T7a/Jqt+WmRZR5XyEOJf3TmZ56083/s8iGd
H+9fb/Qrq2EC8nmkntLkfxpHTi+6L2c+Hj2QZNYqmuaaXC9eLTbSf7pEVpduLzEu
rghglOZQ3C0xKiZGbndFbLo9VmRLWKrrEqqqtxDhGx7yE6q27tWmzwvmQJWtA/9t
ITBRVs3dyCxODpwkz3oCOsw4SIjPJ1ihlMuyGj6X4FqlM8VNR2yIxP7AI2GL3x3H
dbkj+8uJTql5WwHKrQ/sRinn2VNkl6eps30ZvNdyPYZoA/c8ITmjjCyu2WKj6i0O
XxhPI5QbPul80H/DjFmDO2xmkgkSUXiA1asyaPGXwqpSz/eox51ZS9mEhyJ7KfCj
FH5hckXsz3JQA6VQ24HUQwMBpi9I3qNdSxRj3vMvDAReMgqyrbDmavKQofNtOL3D
Eq3hvJjFtWyMU3hZRgfouB5/Hvkz0AUe2+Nd4h1YQeLMrDldMgsswBYxDFv/0gTc
Vg4CdESr3MGtuAId3ycXOG79l/ZMPc8+2gdYmn9/5f3tQm1w1ureQR9/EQdOvpQ3
jHlg3Q2tKjVxjFP5Yd7ekh5FGMn2xXQnSbpVIu8Us0z47FgZLyBW8NNT91DprtHP
JvHJ7/zjP0dehmnQrqsS6ZMsZS0c2DnE3iWiyYs7gyVtfe8FoP3NIkOgRyicctdX
Q8RcopFG/cV2AKLEfUe0Xo/Y8yPYdRn24khG5hL8x3jBMvOdgvxFlIYuICa/CZdL
r19wBbDzXJn0LnrZFPQWt6tDBvQuBJIs3gYDDSiSmLrplwOTv2w+7hWM9F7A0Tmw
3puP1sh8Zt51yxPoxwLtbMoL0hLBPM+yaMtb1+TDXICHLSeSq+RT58WWHCvWF5h8
/rs7izf8oE9miB2f/sFe4FEDSeCoe9kaB8p765gv95x1RSJfPs5AkVkvp0zMS+y0
YWg0SLhb01Ky0IkWkZdmVDg99kpIsPnPptm5vpfDKf1VAxKzJ58qswh/XumvcDkw
rue4Y58UTekwvkF9JH1BC8A6yNTaws2x9zgDu4yNlcr7VqEyqVNJokZaCqXFBm3V
g39iMda4QAJ8lY1FLHaiALE9TLk82wqaGHCW0RyWHJCGbWDTAZ6HcYICfYbz9/ec
HCR+2z2O2TW+F1KbhlVCTw30OjmqlNrh60nibV31PEWdmUD21do1CgyM7Stkv3lx
mpMPmBamjsUcZ3NlHXYwsbxmoynvFlKhGy3e2JIfbdmQDcbijxDC1knZp8/G3uTm
HmlhQ27lwDGCRUo/W7qa3HjbgoEcU+8rA1A9kuijqHNsbY3ywR3yLLLTPm60NGWC
tGq1nPgCXoOK64JqciETi5rHIkXLMuRJ5s21VlZOTQpjCTexZBcGEoW0S/Ko7CA9
liUYIrJLMwHpyYxGc26L1ymdsLTLRjIfOI/+7YpIJHpdIDwswckTZyCarbxPqJCE
c5JrC4Goe2XA+RWYRmI4+K2ApQ8ZqBsuJCCvZ0xqLIS3RIuEgQmIg6s42BXqXisQ
K97b+/7oIgzrb47c3+hD1QxC6zmKirWamj8IOkeWPlLRr4vxOyekY3LQG//ZNCgn
RwF9VVHNRAY6GZvF21tTlttdQ/QJTl3v9V+X3tg91u44oeKWA/Q3uAuQ9sNMn7Br
fdpZVsO9ofimw5Ou2BCDzqKugnouC5B4XuPo0ghbR0KgIr8EU05xfSFeR4CuIC7N
je9GekELQG9kfhsoWZkn7OlH9HMAhzoxkRZVq+zt2pAtEAD75eq1NaqYe2AGrI+H
Hqfa6/bJtyobZqDshyO+nudsuy9rxwSjNvlZgUcofI9xlj4fOrtTYDi/YUB+m1wE
rt12dg5XIcFuD+nOB5UTj5LS+PQiLm8OfokXxzQ4wKoiIZvY+s4hcDaO5GnfRD3h
7Gvjin40xXNILpFWfvt+gXScJV2U9uDfA2SYKabgDlkMV5JY/VxOZlwOqFI7zpZ4
c7Z4djGMsziMQN8xpTivvXTnmt/74NFFVTYmzsDPMyyS0DuIvJ+PvRICemJmylN7
uqaSxsvsvbiXovGyWR8BfbWtVmzzM/L8OLdpmo4UteSwrDXh5Yry5yFonsMvVmjC
lXQJV/E8a6A7FAa0O2QNE9NSXlC6vuZYkQylMmRankfXSlAMRURDXpdMQ78edC0u
b4sPRXxsw8HCUPUKLempm/s6UGlT1RrIUIYMLFhZJFKBfpmWo1UtCcuLz3eZSw0f
lRxI7VHGNc/UBS+uGa9PgVaXHTMQ62dztYbyZkidS0+c4lRVH8Ujbt0FuAMTMoY6
34KFi1Zu3nQHAJWfXtx4K16XIOpsfkF29u8nS+dV0QurTiSXP2vk1s/EnyOo3cx9
WD9JfrXXRpZiBYrpU9QU1SXnbinrkecPFOunzLvWJ62bS0nKvshRcBAHBJTF9Qdx
hOj/5XPEHkKkajpj8U/2MMnynTlnqK9vf5eMBz8SSTWCAZpy/GwQVZWpcPFn972f
JoNc0ePW6hn+pxzmb2Af6vSKQBuQX8m9WtBb4DyTAoxjcvArb17fKlDKxDBiWoKw
fOR7FjIUQ1Kvx7lexJs1N8k7fW6w9yeRy+8gp67BeK6VcMvW04Tia1ViQCkSdLTe
JFIrOV8yWXmMdsfZ6z0MkcrZjaMDKyqAsd3Sr92SwwilNBouQz070PjTZN2sYyJt
hZlfgptByMfqI8SzphRbbEDUUjVoHVlIDZxWGw2DDB5OJ97xHyrRaQPFRMwwqaQ/
14F0jyBnDwkSJQ4ZzWYT4E76YCKoEifaj4zLUK/0faw25rwrrm71WQEin0D1OU3R
L4iYLAHJ9WaKiFU5aLEoX43Kc1u9kg146Ab9QKIlCdkCpoH2tVnPNXQV999/qY/S
zjamxl8dFBx6vrrDDrKWwN+kjBUIofHCLcw/I7N5NfKCmPCRi5XpCs6vh1oV4Oiz
HfRmbjmmfLNjbhXvVZax3Tgx/mRSQVvs+KH+/fuTZWqbMvQ5+7jmP2+/Lb9uPqE6
9pTKf8nylFdUN/PVlLdOuCpHC+mmlOxzkvba5reB/TzXA1SsTWDDfSSjlvwP0+1Q
foA2bcFvStzlAnCMiJDbtaM1ijCrLDlTOh3yELtUNcnjDPi6PENV42bfq4ghOBwc
1KQ+yUXWOQTtvG6tk+QjAHPNv8Gud0sUJbSXVJM2ENkQ9Lb4a/cmUcwrdRsoaukl
owt+kEDxGidDzLYHHtiTGJz67PUb/wQUN1raxRbznB883n1UVNXuOGijGPx1aCwb
5QgusmoMt++IBAZoxDknmJw0Z5vx4libo3WS/xTA+F4RS4IB/JeocD3FZxx1Hxoo
APTeuZ7tZEwiyM/Yn9utwmlGy6QF/oxGT1KLd3AobXu2hTXWHugnjLVnDXussDRJ
BvWBM4wTADvRfCBz49TBtuWwXOjfnaenmwDIsoSUJdt1rdrhEI3CuRxaFzrTBEzj
FRXlkdooFFNiVFa2M0MmhjJE2qVgR70HIM/fsQzpiGc2HelJM7f4wWjRcCqEEA7H
k3Mo6hGa1O+c1lnXSitAVeDrIlpRgWTy6CTL1gsZpQcnoFTGUhYw+BwHPjPe+P1B
cd47GlX1RAHmUbRru2SHYordIwB7dKwivkwf4AvwJ4LT5WVrkDyujnCAvzVZwZp0
n9Oxpi9RBakXbrCiYM3/qNsocywLj7MJ3sKJvebRD7zeyGcpInCJxpU8TKLyC93X
wzuSu7Ae2hDPLyHYWf4a+SqyZEurGlOhu0sh6xPAo2NStPazYtT8b3ACcDoSDMIi
kvh2yMd1U6bA7XdWmsE+0suhRJ4BHqbLG1QuBH/7tGtxJjHHBm/b+kxzlhdRKA2r
yqhB7QrbIiEzGg3J0UCPTaKF8l9i01V/ryIMHGOHqNzaorNa0r9PsSkxMFP2OCaq
hy4YGttyK3fDneGAxHxkxiUmDMCvHQWpEajDAOikaHuc0Dl8aqHpcvam7OQ240uZ
dZqJqfS7eMLtBq3EupG4aim7KGQk12zRJdSqR643SWgM/gvv0shT4eGdhMDJzz37
qbgbclXKG0ky+E3azxa25pA/D3XsirPf1FdMaB6Lags8E7sbKtMl0GOtHLm++cDx
DEBjcTZg/pq2w17XUNvq4gZz7rKVfqvGbS8KJ1xBopF9pFlrvSrFUeddnU5AM34I
15Mz5CkgZJLaGbPw5INBRf+uFHhF1Zf6WPgvypIcRxCNFwvuJqZdTQlUuvhXtdn2
8bd+WGYwY+118U1yMGB8OQ7a78Gq242ETqP2C+xBxOWVMRJsIJt0Pv5uDnCDhoC/
TpmdWmyQWCVlsRLiM5boL+mLOY9tgvSmdv9EzaPDf7DR0HnPFLMah1KIJNZukiiW
3tbUkiM6GZI148KgnkOgm0eGVfWgGrVI0rLN/4uy3Qenf+rEityLJFhRK4Ne4c/w
hatOIHfchVBHYfhmTBoZRsW206LzXd3Mnv5PSuDgkZOq6MNXlft67ntACCNRKOD+
XuXKlXgI0SH8Jj79+k6vJR6CSFRCa8zSprIEXcOB6Fc5mdwf1DdCO4lPlHlxy+15
Dui/g+pLlkNNaM8UfuJKyfBJKokgWdakR2eBsmBgXvGO+QMAcuVxwY3iN1ZB7I6a
LfQhfVyiGGBtaaG3tjSfMXUR4Vtv9/5K0RD8IIJIAegDPVl5DzdCvRYttDWnP5Sz
hLjJB9aCmM9tCHgytGLd8sBXFZfToMZWCWnWphT7pGodpAKFWj8owtXBR6fi1Nh6
dp8raq/XHAzqH0qVjxlVB8KKG1sKcLtImBdyB5GLc1YeiML48dQoDxQm5uLyJVJw
ZschaG+HqjTn1sBuCW55F9iq35SY7duty+sc6r+dCGALqaNE4cH4+ep+Q6eZzZXy
8C4jgqty1ZYQzP9AX8AyYCYfCDWNvIp5d571sWsTG2YDh35jTT3QCRwc3FW6VT9B
MRrcg6EHBIxWMMU6fb/7bWxABRLlQ5LDUWt6inua07vXei9qi1q2jo9RP3bo418+
tHkBpg1VAh1E1e1nIwuWiGvfAkcAnD5CKDGXM3u8DJYcXkSp+gqK5pO7rO0BGasb
ycpxSQLQwCwGS2Pwic5ris47fCLdqllUaEAIJ7Kr0znw84g6pSwULCsVyTxkhEBS
K1+AkT/Kc7OJ8O/66hXEt2tpd3XTPJ3bSmigqyu/7zo9vzwf2qo1OBx3hOh5dEUg
VrRzbe04NwI1mBdqt2oXHIJa1kVaKTAqXRcDYGNK9zetVownP+zP3pSujCigKGo7
5O98hBNJttUeLw+UO+QHFA/GjMIucU884dikvcpGvXSKw9SHKXehaFo6/AU/ll7a
hf5oqV/dxF3tSzXVo5U4zO3fTDKPypIw6bnG2Aud8hZrbq9lMxlrKYCEwzJT+j7w
w3UrMpdNgHsGxw3GC7eU02Q/xIIOkDYF13im2yQfnmHlk7vlNA5Qpx0tmggOTDIe
gaGZI8DNYs8088wS6tbINfyKaxWmLTbKZ/Ic0b/eccKwgn9y/818tJ7L+1qzBdr1
Cr0uGLe2ntFC/IeQUKUQleAA8axZKYmdXSjgI6BUFLnb0DMdwOlxRev7ttUehJhq
LnrvJWsobQ06tu0apyt89Ty+jyhDczRkGBMR0Jv/yuxwu/M/Z44h3OBp1KAlDi5k
Zw/3fgOptiU2voBxNMvop+J15/L0uag5KK8XgrNP5fWLCwU+0vMpkqhl4DI3JiKU
1ArCxODHFrR+fAw3w0lLQRzBmXbLikR7GaWBj+/KXl++3hH0A7IcY//62JAohmvC
GsxNjTTI6Aacyvi8TNGaNESBJ9ztDxH7s7Q9DZ7/A2k3Piv+ZQCGUpX/kX7scaf8
CWJyp3cYCaxgY9x2cwQCQpLu+6IFKmL46FwYfBbdW3z3CD6SR0YLaOCL6EEOK++Y
4kMuHhggQlJlu9E3Xp6jyrwC65VMU64i1uuyyCrIGYaIIEYGia1FM+gAZOiaCiAc
vUNoAfL0+9ABtW7YLB8CQgBhDTl4hc38P9ykfJWifklzTPq4a8Vnf0OMJQcu+YId
T8bA4pN54lPcXTB+Cct/wI0LQVrQ/cQ5z3/jUihBHl4guQAf8hM9+TYG6t19fBLn
e+uCzJp9d+4mliaSOE9OWgdtAPLMppfcbcvu3CvC365wH+3CRyJesJyufayGWQVY
uymPtsPO9Vaiwb8b8jquqgFUMUby5VQblSHzL9yygk6oqWidRBQsvoGlGfL8SP1c
Xg0qbW1M7HL2BNn6sKwRrALsPNhq1NfAXxYxbDtJB7Be6H6yTSJSGK/S2DO87293
Akf4Kx1v7LLdTTkhKZlAbQwD2GwXmKpCMVH5qApKO5h/5Uxdaw1UoejD3j8UJMi9
E0b9+TO+z3MmsLQLS5ujza/Gb3jmk7Wa3UvS5/VruPayEOA0rBzYQ7mG3CYzMHsl
zN43IWtkV7HfTM6YTKHw6qo/TrNRQrSAh0Ggy57wuqp+W5SoDBac6O1X3n0P9sAs
Pu6mytrFcZEalAv8n7fhGKL2F7ZvQFql2bsp9ULFDVhGubJIwK8NUZpwG5R4u+1j
8wzXEx7UaJlfX6z6F81jtBYa/DgT1IK4JHaVx46Zrzy/176fbqxa5TEif11hzYZf
BCXO0BdDDXexmaIkKkW2OGUuP+PQgT7dutDvp+PcQJHft3E3j/4dpMkDOE6tuM4P
IVgaXfBI/rLM9cvX3k9QTPHnH9SHlM37AlP665Q/l+0vwyksGgvs9+gdMPw7/MuZ
dg0D0p6D63TEpKCFTXhKw3xFX7rzI4ZM1onPiK6YLTH6RrJzP6QpoCp4DqR5jQEB
yfFpdrK4ZScYz0nwErJCZXGMtTPIXkC9VlsQiSOl3meMA8B15goVX+XOT2+ZKJot
uxpC2qAJbJoC3lmBpAD8qYQ4PiBJWYpkjtte4vTfk8LelKWRkg6XFfA4NG3BWl9e
Jd0EDNHgfB0/xZtojp+732M+t6kzf3aW+kp5MO6M0LcpXg50iR9M5IJILitaCyMq
rFRE1aOKL3teO76WlK6C/SSvxeaGT2jdgpXZnaogzqd49qx75GFB0OYJyOAYw6g6
hmhI/y6/pM+z/23xOab7nm9ZfN/2aPDqOiWo9uMX/pQxeEBRQu8WbXU1Q64ss60h
FywRUpYG8VGixgLlLBw5kzcdQuIxOtFR8ptZ2TI3uEDOW+9b1Zhr2M3nZTVZihlw
HWvo9zDGocr1R4euNARJ8hvmEFfJUzLv3QlfOxFoOaaGRX89XMuIZxSzAOCgEFak
OlOiFVhTVnTYq02CcjO3rrURkoYhc8y/XsNlx60IEg4cCgapHoWQoriAYEkANmxo
jMASgUbAdSNpfYIIOE8O7uLFjkEbso9LFy0DMwj5OC41jq/AfylQOxcaeJgDZN77
RUaul7rK9TBIrQYk7f3FBP2u7akhgHZHsZa4NNvjpxWdNNHySMMINr/asALIsnRX
xKqRwaW/5fA+J6uRrTDsZZxIgWFhM8wFGJwte4IqCrG7mtquMP9I+cn+ZEyPep6z
S8jz7cDkirHbasHx/2Fx76C7VQcrkIHWTGGYOxIMQvPbZUrCWMxw4RxvtxmT8BbQ
5UC1a39KBtTt1auJdnWqnnMlYG9bt5ZtlWKxjZxxOm/pTA2xkAoJc6TXXlZzQjPU
jKlnXMeoHjDoRIpnt6zGGP4KPWCkSSI8OkK66XP+uXaExhZ44CX93HSu266J2Zvf
tOVX+I91k5Pn0ojFvBkgXI7PZsK7tX2x2R03fpHCnJNjWp6D+9Koo1DJeThAd3oH
MQSnKFpK29bbP7rapKolbXfYAHQ1ubqqE/GSREakj5TsU1R49jsfsnGXmLIQrxH2
ucnKOZwboL0RAceh34m6F6iBULw/XaniDvbtC333lb2gnC3wt/cNGiZ16m2rSRQe
cFPvxPDJNtwLZ5Y/cKzoMaFL+GNgc7SGCxV9hsjhNw4g0H/niC/4HR/C5wx2X7Ps
+Bczi2bnmrSxVK8APWYmgchvnVOjd+sOdwDD/A6v/pfOEhQbF9v10MtAcnIOQwkZ
K4L8hbdNyV5284Bj9GlrhidLuFmwpyG9MH19yUjsW1WFzKEkyaH57pLIHT5J0dKy
HycAe7kol+dK/OmXXeV8An7W7DU8C5RH7DbFAJ84C1mkoIauxJrSKf+k9BeFKeFx
0Qshw+jGt9NqTd1Kztome85x6DV+LQ0LdMjiAmH8q9GX6YgT0fM+rZPbAbU37+0T
I72fxCpfY6MSrv8VnZebj4EpLEcaHz0A42pNWEFoae/4HJxpVDiYX01rnIFKdnXb
2OVJgCFiAvnibfEtcFV2O7Yi4rfmMU1VLYzN88wNF4WV6oH1xeE6+WKlNRqUfUFa
TkDNQV5yzosD4dJDXNAee7WkfZGZmZtxbrZTtsRSsE8Wo8bBC3NtIsWfJ2L+9jEt
O7lhKLmU4d4rwz5AeFUkINkovbGatQKFaKzSBFDeYd3QngdaK8bnPrjUUAJ4MzKV
8S5yvX4CufmHNsxN4fvdSnxLq+P5WPBvtcdLjuJkI667c/bKiaCmjK29AfKZJnZ0
Dp04udpdgBsm5oVB08dm5krwAvU5rxa0kKDwpYTmWc7fsEaJUylb2tQL/lQ/UH+G
RqPvs1COk4vpOb7BkljtNia9qhssOwSgDXP5XCFtDChSmkLsigANA9qOpL8lDy9S
LCrGxhgaIlFFXLNpWwcSmw8cdhm1kdfBrDfVra+4izCEdp0YZTpSo3rOSOtAP3VP
oCjFRcAJuZ1sMLmN5s/9GDDappOPYpJNrijjoTCNge3U1h3erF0LQFHc1r40s3fG
Rj/hLD6qvM8/UgxDsiEbnxLw5e5SCw/Tg4LxGwaKQ1/AMMrxp6UTAJVy5xSS/Ttd
MOR4eSOhe/dFNJWWxTZ8fWnOfBQ0t19y+2pjzx1UxsuQ4USQs2uLUBgUID2CG+Om
SDwo070tYbFKzPn+z6UKVUtS5KbJlGVuHzNJF6txRXiNNMySniMUdgd2PHnJflUo
xdG86riQOWgDuzta+RIKwqjBW7ua/lMxoC0C7NYVFCOQnbl6ZJa1RvOLATNnAeu/
mjY74T83MDUt0bns0gg2NnyUqYIbDQVlU2LLx0jzT055M5qT7vFLylYZR0aFJAx+
0m56VQbDncqqmwG3EokOLvnDfjrv3YgDAg71G43qH1OLfCW79AGF34qR33DBLpkm
cJ+rxSB89zZAYNbvVICxEciSXssiO5PrClxPydrXDuu5hUyIhP0PK+6IE9tf88wF
AkZYxy9/81foohgMhJfZ1/kiyyIJskYFcHQflsIxk2Zk3bVjnHTjxbMqKIpIsIsJ
SKUoBYvBsCo6ibRAfwABCG6EKwgJIpgSj4M0KCZ+sfEycBJAVDDt9bszoPcyrxlf
jSUZTjDtEM2FJx9lidFCISKyqmsVuzDqKDPD73gZKdH66FHvExSpmqSaT7iDScuz
QRG/cFidkK/6N0u04Bb0E+PPQgsG9UbPFYIe0o7EO3Q5/Z0+uwXoApFwXwNy03rc
vpCKMHEeSR5jCUJXZoRpHu77ynJTVVWzA2MUwyuAFfoyl8px5Z3QcNftOtphReJ/
O6gZbth5OhQvcWjj2KQ7v8aDnPM7DkPcFHTP12f8vG8slNfMKXYvPbXtMQKoJnzn
mVKyfYibin06Xoc2KVh3yyZIJhbsw/8CgJD07o2iRvg480rP+xBsLhOELtJX6/qv
NnP5wOh/t36W4tLs5Bm7qVO0XmWLEgzWdVZRgzb5HyPRSFo6TFUa+IIJPvEQKE0g
2yqDtCCs5yna7wm1drUsGlS1zisorKmfEJLjM7Ug61VSHEjnH3Q/Mair66v3NrHo
S4ynybHSrXRHS2UdRZRE16YIgI1/dsA7kqr166J8KgwcyMVUdTL/HIp7n68vRgcr
60Uy9zxvevYF76oxJRB+D1Jarr7dKpa9YEDwtXBeXgKMn+7/WsjHRxEYcEcUbuT+
fnuK1SQh3TkzOgPAw37s/SXKfWdminfZitExmARA64j9P4nYahGdQvJ/3E10Pg4b
GhWTF9rZgW9kU4VEMt3NZ0VQvIOmgzO58MTsIGApDvaPUcdLhRoooiE98YamhLhX
bt//k+m9maICvDbsLTEKQvOwWhIN7r/+G0Vnwwx6b3uvFHoj3m36uH/GGITXFf5J
GPt0txhT4xepEhii4ewjNshR04/k8SUM+odUW/Hr7FlrJ3qM7w+u5ii4GLS7gsj7
dwImpkCyQsCxDfoh4a/zBh5KDz28vG+BvaovvJ+K0wDDD6qyMFpQxYVD/H3odTxG
KCMOIh3BNah+EL2p0Ca4FG0Fh2fzyky9EHgEsC3EsG9wqLd0M+BHqyyhBCI6CU3T
EHug4QAnYWXscbDutiltd60G9DDZHOmVJPC+ZFvxmZvwQgzOcGikaCe6ShGQygJ1
HboL/Lzk5gTsMfZdpAxTvIJchdFB/eluLG30qh8TOxXpJ1viYvmOuyWPh/vtPBH6
3GJVi6z6n+Ha9UVtkk/mwLjcEV8lua9ctIKAU5Qh0H3wBopyhKbBc5+LYdB8aqDi
1ENdWtR4QaFKZSWFFnPjxd6mSW9/KgX/hfrv2GEWFzy90dOsMJqXty5GyqoaScIR
h5IfD4b/TKlAzuBV7tlX4Dp3A2Ct91lDOElq5k/jnE7Ys0Gha//Y4knjBE/zT1YY
6PW4bGyNlye5xWR9cnJ1CVKC+47ndscmEfcWyyFKMmGqQjkf18RWKmtNrbpb2UTt
bjYk5zMfp0MWkxOnGA5xd3hnjJliHhVGDeSB0ABWZL6cpst3BmHMXY9B5ruVumgm
ov6eSMWqDOChWbsR70nSGTJ3ExFL24IRUCv1q8wwOl7uzV/W1gL378Fw7Db0Q530
4bFOEZ83HWC7143bY9+PC3gXRIuUCWI6xELBXy9jpRXuvscT+GceO+EMJqupmEV6
5ALlQYKYkEt3IK/XypW1q632P+yO1kCdzALINHbyb/UJeXQYLl/d6IgWIFMDCHyp
JJXB2v886GFJCHlgxBoUhoWX5JfgqnbulXnCRBLz2pOhvrOaRlJCPgvXwDPVP9R7
it0iEYCfekN6Oydn+eVglemm4ryVF9xNybVswecHFbUCssupvtWR7SB44Iz8n1CQ
bfV8h1jaw5u2dWeiUMVZ6jWYbx/rvHkBhhlXQqZ4nZLYdy5piNPAC79eFYay0QH3
ToSYxwINBjhrXHmN8L61MZhoJ+19ZitSIxhnJWiIK/AAcYsuE/dTbFwe/xaSzvlt
dxVjjtbTVeTgclRJRjpZ7Www1R/QcSivWXowsTdnIh+yKqGXsD/9zKJUFzPUzX+a
3Hmog5I7Cju84PkdEO9qro4bk7lG2hjIMEfg/CRW/zDcfvIt+3BgnAAvx+ID7cwi
odHGLJDMQdQ/iNqb9RT+WNefNPtR4CicdP638OZ0dOfYxvig1RVQYEmG4M4rIzHj
E8exBy4F3xvH9KSeT1v86m+aqmEjQu7jbiNsGESW1qCW9g7xwvtp3PxvqHs8rycP
zKJrsqe8awtJFTMoCZXaa4bqR0XJCSraivqMBN96Tk4MrDwmwsIB34Q4R26n7kPK
shwZbZGSPnkcprHROvfFGYJJUMnWXGczQIIWZHdpbNEcIr5YdgwacE/FYhSiZPp4
bZrIBvfm9fEkdtZxhf58VTM4cGkI7pp+QvcMScFQxedA/ZUZzrMROB0fHxLjKL52
kzcBITL/I8hbfO9JisU8P3j/WX2dfpFOMZ3p4eQEZhFHkQTMA19D4Nj/YseCb5tV
zfWUdOHhcRivIq3FqzyDJ0oGaFndW5Y0m63kMKknaoGMcatYICugeOOZxEaKXAwY
hR/bYFriUtc55tqhaA8DxiXeyZXZLxXGE973QcVvX3/wFg3kDdLt/O2PnP00bMBE
ANq9EpKSz2R4/n7iNAYRgs/aEUqWObTw+NXtBg/lSpnZn12q3b9B9jlD9WwAg4Hv
q9evg2Em8Sja1SHk/Xjx/KyYO+VVfpO//sI/9seJF4kl97VoRWf0OE6yDkUADQ7R
zy/Ls2sJv6FGdiyl8WY0sCvDzHqxgeWe2oElXUmw3tQ1Is+Hie1ZgOYwlzmLZ+rl
OZtiaJzaO37TW5GyIQhsEkbHFj4d0iWGD5bB4CDrFaLT5EF9Z02uPhybr/P2tJwk
GsKoyf1lt/ZO8lj5TPD3NuLeku1oTGgaOdKHkH6j8ON9F0r48qR/h9HVbH+NLCYA
h+6VjhS9jAgOCiSspVVFPes/QWNgG6hdNEDGASGStONE1rmEaxSkBGV4S4zqNEOp
LclaCM3n34pPSJyZYk1RG17SUmcvA4/ABHzXDy2VKqCSGZhXjkBjRyPO3unoo1AO
SCV0XYu0IhI9DAlMDvyVa4qxpJfOPpu6hv9ghGykxAFC5DnTy1lPO4E/yZ+7RzRG
B/QrSYvCWrBSutI0sQFywyHTiZtGNr36VR8/az6VDFz7sNKn/dPjStMi00Xvpi6V
vI2K6FfcD6eG2KCX6FGg2CR7tj9/AV048kogXphuHPjlIf1S7U7qZQE7KOJyhQfN
5V+RFS+EbEk92bM+tje6CjdNb4226Zh/b4ofnw9CcyqLH6eIYQrJjq9c0w1buB4C
TQPJUmSM6Ir2MNGdiuopKqpZn9FSIBO49NXdCKpBERPKBcbgazMUBDHtxwg0JzuT
iwCHF/5l+JAosxRRznGjALoGCeoHe2t9YsmzGIuCfReW88FlHUaaAhM3+0IionjI
gLgbP5DNWc5i+HFrXDRhLflrgvUnfT7Pe+/nRm0fq8Dxtrh4R5o8YjHYbTYh3kdi
OLDaZn1XBcqIdF9B4utVZSqVCE8DGMoVOjR3tT89mq+mx/4fUKj52dIojGJWQTML
f0wObjTZ1jDiLi6lNAtpHkWAdfUr7xLW/HFN6fwIfNgw7pcOJigyTmNivT/17UjQ
rQtJVtqJ1aufkTW0QqXB3KjtYLQb/BHgeosYhsfmt8gUq89xFNuWaoNLzSPwQdUH
Z5kJ+0UvF7ckERkQXY4DvQRvtWZvlsprWl6Ho4BREcr9AQ+gIQrPT+cIfwa2+4O1
tTYoxGCFEfrkXte+0tl6R5+eBKYnGjGqu6SegbS/llAun/wbEjNhUV4w9ms2G6ki
5n4ypxS2WcNhndTxQn6tmxA4+POF7A/CWtyqw5Qs7HnnhDboB73YGmNa1sW9kGN6
9JjcR3xljcJd27/GT+6Z2r5lg50ZjmKAxVETRLpCFZtH+/OnNntBwBuk7Rr8znY4
uQ4lViYI0RsxYLwb4ybnmq2yUPkw+u3JBaY+3pNlOJanx0mu/SUnmw1KFAMMIVl0
QQLTgnQLF70jQ/lmqLa++EixD+lB3gvloqQaLik42T+tB0Ffj+xp43hqeRYkXi2S
vXfs6MwN7N7TN44JCNmZhyYxWSRvhwdLANHyx3dZ019VyXD4yESm1ENrHUTUa4RM
WFPnIHWzPwIWcbAgxmSDCuXajyyAk5pbikmmSnAbqhlAJBjL0c71MlyhmyBWzsv7
IhA3XH0q1syVm9DBtbW00P+yprEgLat2ibf0h2Qgyl7O5zQdW26ARcQuFiEA6Vgs
hTS5khwS+u8/kuOK4x+Lks5EbbD4Sx8YmW406hZF26kQFrbjpIk9xsPIDWNbeFkQ
MsaRiQVw8LfzVaQWlDXYUXvvLug6ZCFiySiTbTDzZJqAOj5/AIUTRniQ+EGXuHDl
8HGDBgd2jkPhbL+AcJEUkr72/hBfYwbVNaPemOiSYywz8uvWbPWLKGzPkpHRCa1/
38uiaGQnotnGTcoYv7ZRWHYDdFrGCEL1HZmitTAZRkztFKDI3tkksX7w7bGsmzzC
pc52UWVVBMNvpbD9v1/5BvueOcG+/JgDPQzHqp3lQ0lnKFO7U2BFCEmLWNu1ekLL
JESPZpYg2alEKs2vvlQlLpZVdP6g1zTQEL4l2jFh/9QftYDF4cPX1QPLOQZA9RDf
nKQJPfaB3ioUevnJWX8ZQnHXLb1crbygSixM1GOjiWKvqVjTcIQ2+Wjy4r5d3lGM
jjO9BKb5x+DTbtkg157gMqtJTTwRGyrPkO1GeVLwFGEKnatbycHo2RhDiRlCSAcY
HttDGuBMkEJSVaxkw794pdjvzGxSlphZX/aPcRNaM64vZUOJTslXvZJIwTgPRelN
8Umt4MAcqI1gdW+8BfMEwkGtalcgDVrCpgcqD9UnS5jyiNCmQVOD8guUBlCSdSLC
ymBUqNQsqq2xeE88If8zTL0zLYPCjxbKVZeJnDODS92Gzi8WtLRTKc9d3fgwdVCX
JZiKKfU7WJjnjNUPcWLUiWuDwgSe4Ne7+864qiG0cDbjlY4GB5bchbegHOUwbE8H
JD14SFZEZ/zMHZjBj14NpSB84/wdt8H7rM53KP6EwbCwhamXs8QW56JTw0liDmKH
1nKssJIRG7fHB1W4I85NnJthmire5g5Gs9c2VRhZYLe7Ds6LYWpFrHzTVJM7fmsj
WyK5XOLwPPlUfnr/Lh+GiqmhzilAdKfEhTQkU3doc9rxxt1+Bm+ssBL44tYCUfin
8YeQw7+ymA+0Rze4pNeVm2VQzst+iCoq7EKiG5f6Srp3g66jR8V9hrMPRhQQ9PEV
jI+xACqsAZi7MjTfJ0EMztJWdIInaigI2MF8hSwj5pbhEwmRq5qY6igjEMuVRnu8
tY0L0Yw0O3hQkSPx+Lh8zfD3Z6uQBmEOqolu8uemp3FZoYH6a8uw4BVi32S6kGtY
K0URGR/EGEOIorru/J5dwseRbqMH32lAu5wIAxJzy8124MN+bHMKnFSAJ5HVdd/c
tqoymvkD/3wU0DUtlQQyfzE35/AHzI2CKGpq/Dse37KU1TvLwuMl6mWvGRah6MmU
7PSQylO9Max/wNY3hyIDWAaBis+09i0U69FJEAyBkfZrGPrmI4Les13+nxuKAred
LzwVKKZH/fneevs+A+LM4Xedyt5QNfU4y+ZRAbXtxd8tYF5byrJR9X9BpDSfdJSX
wqHZuyx+Fk/5Jkorfnunj4OEJfHese3/UT/v/f3RmLvkhbZcBQkS5Z6LvDZVD30I
y5sIosV7iGe2OT1mAf3nm0204BmDbe/pHspbGSFvOJDq85RJufnlnb7iDKnSMX9f
bytPDRNrN3yBqyIwrzRQw320N++I7zGPqQ7u0ItKJUFCA4mMaXpcQo3veWapSQvl
PWdIR5v0pq6L8DxKELYzrRAGOMIpOdTIONbljRUhRPpn7lw6RMxEykKlsYxHg++4
aOF0OIeA8wmn4Im8SFfN/3oftCBSWeHPIm9oH+wD7uNFP4BZ1HC+AyGsuvGKC6cB
9Uh1YzrwNUUyUed3+rlVikes9iPWCeMc2VrevvlPdz39D8/eE1KV0syfOoOJblDQ
SrsK5dWybG9t6bworYTRd2m8SqfxIq+xctyRITdi7a1EUjTZ4NjzSt4wuyiN2Ggj
BBbjXsmJKkAnMsmDDym78H/jRbH0it6o5rXkAwbPokdWMpaRQSVqSWzZSSRQ0KXB
o6lx3iy59Dr/sKIlhfwbJIyzSGtBmcjzIZbVUTUhZt9r5dmoHr4yNTcBn4oMf9xg
u+gWpxLcUSvJu89iCOzcEqkgPnxP0kOkqepMAkxNgUQnpsbCKXcMz8WAVKhffpTx
VV8ujvhikdVkrxqpVQEmMsq30wHru7GbGFP3XyXGPVebcpZ9eTO4KzoV3CyljOVf
rYQsPyFre95VGB/YIjWcrIQAIM8+9/IeSPspdecdw5iv0md6XJ9FfY94ODh4NSsN
iouP0GWa10i7rHHfOBih4OcBc/XifatyTCRJwJlGTwPKIWpwyU6RVtF+JWH575D0
mYXwtPbnRdbnrrrEBd3Wv48bFoVdQFXonJPuZjYd9D97qP4w9+6s68PkAxda2kTK
5g9PreDUEY6cpvrVySL7w9kbyDsBUjKOxmoOncX+rTh7oh33axoDvJmrLDlFRo/A
yomi47+OmpsAdIfDoCWPrSl1202BL9pi+D6gejAES6KyGVqlsafNjoEZpqRodyNk
AdwBcHJj8j5VALOYNd83EHSlymMuXaz8u85tlo/3RUIIA4rnJujVPPTOZcRuDkKY
ZIYg16+N5Vp0EP5/SstbWEd5/qKPCSLWGG+FywJlCT4HcjzBbzFiRC9dzDA38ZVc
Njpv+1doSmfea26IToz70I6ftXJKk/eMzIpXcXNKlzk7Hm1vnCC2+iEyHAx2R3xg
2clE/HJbaY/C/FU8sebcJ5tyXUaEkBwBb3roUetpI9qVo4NOutsG4po7aSrss2hw
rj4NDMoJsXU54cluj5CcecumJbo5r9kVX53ylics+8ehh5GJzlsx9/NhfNQz96Up
03q+Blpt9qOkw4EbmrRYfIurl0eeX3EbKlikRky4HRyUeW7cCGNJtqeS7SJcVt1m
lhAtMJADsOVeLQOb8S3ku+SAfsxVbZiv53ebJ0OjFtPYoC5jz8yw3HZ+1PA1h0WM
zPbwLhHmtWmldUwxHJZA2DQDEerJNlBkUAhbmhXsXWzbreq6ySdVTUBsxiW3Tb60
n7EtZ6Il3OEvGjVbwicgSuWc8Tu2KvJQm2XBz/678cliJV/t24LOEXRBxsBcJEoP
l5CSPjMXslXOx8dF0ZQ8VK81A5yQ+HFki5lmFeJ3xv4VDJkROQ9AVUIcHBXGtb+i
egRCrYsTF0sQ35VJk+BtrXm8ChU4ksPERrHZovTQOnFILfrln4MN2XZtL+lxFK6o
AawPqqiSQNBP9+4YZw/aASe2k/EwHMwruRjHNqCo/yfDS1NGKvKc28JhMGLiJpfV
i9fNIlty2KH6+5yaXmLYN6TLjJtRYuf+8Fl7CIqRPxthihs8kTHccXDatnZCbAtE
oBEAp05i+3WDbjisU0KJU1uDQ2ByUyRGUxcHNhyDUfTTpspjZDqVC69KAuA3OoMS
v2ItxMWiVndpCjp5OlYdK6kvWswBZ0Yc9vJi/W3pGSUp57qoFNOnq6r1B/Zf6AxK
qUzXtzoawfeuRTyz4WqGl3LyOO9nqSE3kSvRSU0JYoufYab66SzzZSZtNf5ggtv6
cz27BexFA4SwZgPZLUlFL1lrOM2MovCtyOkKrq65sFxhL8/FhmMh9cZpBQR4YSf0
x34oLvkJD145TgrIBsGGXP032dVg7KcRL1UpyuIfeJDjeKgHQUiwxcVF35/Wjz+z
Nv+gx9Q8yMA1XEoSRReQCk5ejfw4sN3Prn5PEFOEm//mBUmLHFO3fTKSn1x9Nl/V
u+3FPptZeYB0zWAvPOsPWEUD24COQl8idHbluroUdjB89Eq7m/Mzs4Rd/YHIG0S6
OlDt+R2i3KzweIWQF/sNOmXVedQjRr3r0pjIND57M6MwSqDy3zg8ZJXBmZOo9Fj+
eua103Swy3FnXrD7yl3Xz9X803SdrEmxuvOzUpWKug2VLt0ULiG4jqedillX0G2+
BeGuTZ/zObDJ8yTeIHa2yzXPZG1A/EFSMeWwmqMoi47Si2aZDXARJO2/8ynE4SYM
exVDcWgA10oZC0PZ+LC3lAJqJAVNaOpWMdClmh2J5KTjojkV2IcEchRX4OUYuI2U
Q00LVG7M2SO/5aEHMHhbwMKRUJu+wbKNMtsle3CnXGbjei8DDWaNSeOMqvZ/uy/b
pswfTwL9V0IIBAEpCH+/vID69QsIW3w/avA5s3sh/UFzKMyrnrgTpMAV08U1ikFe
49E8YyufH5h6UNExFVUVReSuqOA6V2tmDFautAaWAIGRl6UCbSN0hl9eFXrvCdHV
taOJgATD7qwAuK34EXjK5Njd4vk7+aHUnU7OU7SZMxG5pjURxzFpBCvA/312M0YT
LZqlrXliRWYKmeiaRqd12PfkMeQY4whkqY/rOfJymkKknmfUfEk4+ZtI3kPMtcH9
HGrZSF3aIR/H8g2MHFs/KM6odJBQxgk3wyf4nrFOnEkV/fv2F/UvDR8I9o6hsqKm
u4Q5F3agRRFOB4jWbz9LZExO+VN1dDMCVpNXujuoh5PDXYhygBcGSx/h0dANLUi1
fuhP0LtiHWVbkkEfJwvgdqXWux6z0stIeDMPB9scFt8/xZqRR5ahdYZDoFYlJ1wM
kEXrq5zWGojF+P/WRd4t3ZY4oJQABXYe/OlAI/lzw/xSv42QZ4M+SDNCbsQ5Lb03
OkkbXo45WRx7FKvAF+P1nbl6I/87vWo6Vm39GEzSzzC7ewF3hsgIfyNnsUZ2pi/b
UOGyRepggnUeJvVrfuB4YT8MfKI+ybHAIyfVgp883t6o1eN8/DmWtpSHSwKDJGcN
fhN0UhkoXqr+eYlxyc6BnwwyObsBZs3HGjLEIvbWAzgrrqIZeiWcMH+eqZY5w2nw
HUCwNpu9VPewfGjPgE2RGox5sfYMIh/7A3EHSz7DMCJApHJFg30b141uUIAquueU
JtvEJ2FzRfgWOx/C4U7e/PYuMMuzGRXreC9FOsfF8IFGc0IWtOR/tqUoHQNlMldZ
gp187vGBSuY6pxfyG0Rm2/FqrF3kk1Wa/h3S6G6PcVP0smYPmxU/AfzMsS46DZvc
T8RvrDqoCYRsUYa0VrBGkXYNvOY1sLtcW/1pfPRlwEJ5+yauJkjkvInGhlZcxZm9
fC9pHzuVopDlqQJ8v/IDks5OG8qUD873iqYZjDfknTpT5e431MR5XQIqflKnxHQV
7Ce3MaH5uxgQjFiXQozsGigzpHJ9GonuyQxAplfWbQLRgyLamfgQYg2FrBt+wv42
rjDySesM05VS7QyDmH8vSsfUdtNDwC+E4TFtUUOXFMRgNPZB2HHPDcdeWz+1f1lC
pkKdL5V6aYNRVE5fzjp9k/We8uxaK4H4RpWHLV8fXBDZzsEwpZs0s+0t+KTsGGZ9
vXc8xxsd4W0bErD/0vS9L5gFx1W3X/s6llVywh96j0i1x5nl9xKJpYWitTJGl40P
QMZDdi+UJoAMoyuvIwGMyPZ3PgZUqlwbnjq6rcEz1oFQMkyQRLCPGq6mxxd3mBZI
Mq0VvHZg/WXdjckoO7TQzdGiL9SIocP46nvrabQP3+IN4+BEKRsGlTyzfb8Yrcn2
jmD5z0k0YW7XA3Fw7TpOhpsWTK47ATr0kfmKNxH8J4xJXIDIaNqawFY1UO011xWq
7gPB2WFeZhTaw5IPW2pTqpJJbohK6/jp0MbyjVfSkMdBNvG0e4+9cTjxJDh8SZFN
/JIJ+j/Z3B0Fo7gFic2HUd+1a6JpKg0QBjuJyviyRRjox6djEE8a9TfovJROdwvd
L13YFVZ6CcecXuxzpmykAStiQmc3pc0+AmoQ7gF5cKhcePOAdRFRkfaUlNFVnmeY
YmpU9SLywYK+IMW+tg2HlI5xQ4OJ7tLKU5K+U5txQmEdzClSulcr8wJRGkIy1I2A
daEVFQnn0kjw62BkfnmycJCi5nCbOdSZwDN75j2tq1XBQ+5ZPrCIqhekFXmMobWp
d0j9VQ8kaqcFvJ6uA5psBQZNchRzIVbLytCvOmux0yJ80/UmtCbH1/s5tofmENxJ
aNvptxRWQCb/nKovAD4U7/CxdgBvHV6GPfqP8qy27OQuof6hwlO88R1KtUv4sy16
nsuWz2LJFZXhHdHojVhgUYFHntDxNYily41m2YQZjZtpDuUIGejc0Jz25NifNWer
Z52n+3gA3KbXPhwSm/lNMjhRmvErI75OLkEtwSawZgijSiBy9B/R8Z89qFLGO7or
IRPZqIbXFPUjaeg1XKaXUK2SnasjtBJam9j/F3Ajm7pc+qMfr24OkBynB8aYQrkM
Wxi3iPPm/gT1EfD+w9ReSZLzde1ZNtHTBzEJJfkcCPP/1ROzTj2oy7eEHr3l3tTz
3Pb4dnyHqr5eQAlsJPZtfaAsg/IBFDVv7v4pFZm5yug/sMOCMb8yXfgoK7cdOWMM
hb1PzsF6Jrj1XLd12cLEnwJiAa0f94KCEXi+Xpx/wYIq18XMVnSYT2mGSoftxlY5
Jx/NWWLhxP18BbVlSDPyyj0f+vFwgPOZ/mDLkyGAYfbP4e8ktymgdL+u/bink3mF
7MGbD2L4tQEoABB4zrOVq/cMk/fi38KFOLOY9qHF0YVA4sME8Q5VbC3SRZjkDS2p
fFEj8ePNc+RiBKKwiBCiTNbPt5tNaIr1ZDjklUwZAMSCmSrAEvIav2MPBXSZdbiV
QqaDNiQIfMsy0XoTopoyold8r4IkgZkwaRMDOOuiu39yR4p+HMKWZSNfLPAtLgn6
eBGno7ayhF0TI/QxARh3/EXNVbpGSNcTyiMZXlfkz/dw+VfYuacER7PNXD+1r6h8
uygsQtym6qGA//8dzzo+b38dfMRr39ywbTwzs7oTh1OFiWA8MKuaaLL7+5z2FEIE
yAnThUtDtDwF/SNV1NPTihiDBI7p8eK88hKieys/NMkcKnLB8DxWxDg0pZL3kCjb
Ege2zpqVFRliG9ymyRZrr1r8kncA5KA2GjmbECS/087R4PsPbhKoZkZdEpN7hHbK
jWXl2uJF5Jk/yKMf05TDAsmfAU4i8nMhCQh+YY8vYTjTWQTWor9vj/taI+m3e1S0
5Z+2fQ/BkQ2LYl27/qyg8S1o7owuquWrOzcXsNg49ARX7nxHx5HlbfFRNDq9ePLl
NbW2LuWIrfFBHR91rCqW6dRaUeeQdGHTqOrdr1dx9fwXUCjRyc8hxvGTDHE4brE2
L8dE6J0CthU5U5KR4Tpjgg5hCmj2v0gzhXlgHklwEQluFV0Os2wSASdJk+NDizMd
quG2aeWCDjIAF3tLBK7pd7YD8/DH58CQbjlBesRRdHZJn7O/cc2X1qWEeYHW/DEM
P39QgZNt8810icrbk4hhIH1EYTNA5Yp87AdB9zVWLvXDHWRvB4ciSYIRkxmdiYh0
bGNmGcIk2Sus+XCWMoY9Iz4jm2Xmex7Vh8RRgoeEV/wAVxWYYQgwN8wYSX+QhHsy
niFOYsW0dOX+6EloDIffFGzpFPsBYUWJfXKcPH4QYVQ7duUvRb4VC9jpdc7YR1KK
Kx9Y46KP9Zig5E5vRwEk+BZNKFq3rSGIZEKB04eEu6gNI1gvM4B5TtG6Gw9VA7TL
wrc3StYEoca443+sZOWVxY0dIYXJXh3eLZ8Ne20Ra/TMLLEKKaSCcSgMpNxjp4Jd
JqqfyJha54pjjHzCtbw/i3pB87pCa7V7oRqeJZhiqrL7cXIThPrqboTB6NtsSTmt
8xcxlEHmt8kZ2FF9RwREyxjVRlpZIn9pdxd94uNftGMiUpqHfDPstk2TUD7aT5qm
x03x9x9FItUhL/54/60Xj8h1WcIDlHXzEWBxKTsEVGwdje8xdwqkgr12KShr+Io9
dvFyE8YJHPOtOzwg+lcwuT6vBmPeUqmOVSDQckx74vcxbHDNTWV4yplxGfVljK8h
rH/xfcIehL4tK9KiX97WlMvevPbnuuyx4TBkhsvFz3FRy9T9lrOMGFP6ksqkAamG
amwQFPgZYGzfGojhMEpAl9DLhXEH8ED01XftgEINF86Oc91gde/P7CCUiSZC06al
rZPY4VlfWOqhTnjwL2h58IC5UPXg17TmSpJvP7RJ2ELqA8yufBZ3JM5WmejCLLXX
koeUiXKU9iXgWhI+qjyWsLfhGI7cRe8txTLm4PAnZ8kvBWixAQ4ckOpBQ5uo6Hch
/VXoTuvKI6076vZMO77hbuxZYUc2BvC1EXMT0F1BjlD7PrOdWyr1x0J7SJ5bK5bx
cl9Aq3Ibd/ifYkC7Lf/zy2msmmjp+xfMK8cJJXXYu4tHyqiy3v6wEpJ7ZB6rVfNc
T7fSVokWwPlgRE7c/ldLnHdNNi0QmnnLlnsprsIwQiR3EaNYbTN7cSIjohTgDjT5
JxpTRYWuxS1riKJKU7ciHFpBay92Box1Xc2SUh2NlH2ejdoPR/nVqS6p1Dki9xxd
wGCl+MS4bR7//i6PYhl3tKnZFY+LNHdaR2wdCUqICUA63jeW+tGGKYD03kPXNWUP
cqzhAt6eUJzcNR1z2CC0g1cCSgjxSO221Yimc4YrbXKvQTZchM3WjncvhYDTAEnv
10qAA1Ioezph5Y8xpMjXeOTkt9RmWqw1CTGkE6UzMZWNX4aNTQy1aBRvcj0sL+2S
gI2qNkM+eiDoBgdFpMutwZD2Rwd9IOpQCOPu54tAbzFt3W2QCjko+IElrdiLF9N5
RB4WzFAqxIRCEsrgbn54GsOz/p6fCNZm+4ayOHPLlndCH7+9L2Xsokmq3XVnKAR0
lXSP6WyEVhXK1YuXGkwtp8ikIMdOLkMy9Hpqh5EDTRmmCcHEicpuBphqgMi4qOoz
u5C9mNW/XuHXQCTpg24OfjvbY0e05LJJTrm186qIYB1Zg/12xLhyUr4SEC9NeFAZ
oTfNz/52clHF0o4oQnUUEz5yghvlnErcT5yDW7UydA2vmwSXW53/iiFWbL1evZJN
yS1yZ5zym90+GHuACXoiTnGOCyY5BujYD7Ch1WvfiUCRjCnOPO3LtvTKW0QNRoX0
ZJjroOW36qAVYxAgSQfQMQaIPhUxWz6faShJtUibavd7LCaPLXZG7dw5fXjSajJM
La/7j9x9gQ0MjHrS23N9o00FjFuW54Rz/i4qjlzRr0FGr6F1Dmh0zexCArhyGo7M
HqtCiZLf2BQiD0JhPou24iuMEXGMGZ4R97uJrV6c8cp8flZ5S9W0Jy7PusedYi6/
fMen8HbYnK3pC2R/ZU4bguQZ2U9DK9x8dk91fIwLi7EPcZoq81FOBOYIPICzYf4f
XjIaUcQB7Ps8dVdMetLyuRqdvG9XM46a/xzDMNaJpYA6KuHamGKsq6pbXR0NQgIQ
lURxyspFH/SKjlAs9KFHPJwpWKS2TJ0V0v9Nq6CcreavdoerrWnyRL92vqa/Ngnw
Rfhez99SXecM8/MMi+kJpcBUe7veoltLP3czvBPW3pmhNHccE7ZYHzdayTgHz6z6
SgfRyQkZiJRMxexwItigM/nB9XgGCNp/oXLX/iNnDC6Tyy8bn7ur73x+ayqwcuyk
79/04G17cdTfkWC1JdVLeh6cZ04qpKNYy8hcebgfLDBtWdycU5zFAQi65VMMsb9j
NX0nvZplQ0O9TJ2jSvNamoMG1aD/achC/CtyotiBo1R4IwtuyEhzp913UBreevO5
GuyOgyJ2H64u1xXzpltvUfNZltPCciByhrMQfWxlU0HgXb2daNP6thWLbgVfWqnR
pIlCX0w6j/MKU9FdwpgRUPZR7valBDZNlwY6JYFvVRTq+rIJHCRVpVa+HZIvVUxJ
I1DNPFaena7umlZVBSLEFXFmMg8QyQDtOSs6wYuV5Cj3oOjpo9JCNOJSeypUxW4b
X9JXIq5XEmBOixF2gpfKyFKf3ynwGZsA5JRVbpJs3IpPS0wpqKObWyX++6wUU27V
BcuJ9XdLQpbgZ4KN2ksrBEbjvrvrAvSvLy+zmhFwQB48IXHKDb9wVV5RQxHIpJvx
GFj1CRs2Re6OAkJo48COpfgDl+S5OMi7EhXA0lpSEitWovwQAvZupxKMRwQJeXkW
pbn+wCvP0b+AXR2re7ft4N8CmRHKmXiiOKcnCwwXX9wtLjVVrKtIZnNDgN4PNIr3
Ora8VD1wE1I9/KzEu1OzpNxNsZ97qSyDGEQVIIG4weQCG2Q/Fgc9DD3VWvp9QLA6
M66xFU4qiODCR7B80rs0Gz89pErugmM2HiJUmB+hK1tGLy8ZWyqyXMtUL3AF2tRc
ixSjZfyHL7UJ2S/Apq8oN4LxdmpmbidEcL3QD67FzB0M8CBuERwSXyvEMDvypmRx
jqwlT3GZ5296jc1kyTh2MNEscp7YIg2/KjPfk6rnFwxuduedPeuPsoDTvecfdhhQ
R+aBe2sGaEY8jG5b15jb5XEwaJUaJRVHdPUBE06QUXiwm5SHXBYyqCZ3kroeRADm
rizDGQwxX3kdKLMC4T92Ti0ApjETPCXMwgTz3aQeUNttw17rK5UeYcP7eFERxwJB
BrZz6eA/rl1deZkRCgVJEMwS/MBEyGf2QnfqFx4p2kFVOXv0X6QBJPr/PbKZ+zXw
LCq/UaYqZFMTbYWLmF98sST0f2o7oyDesjmQ4VdfFZw9xBpP0MGuVUSAyWU1IKhu
ZzWg0pOKCGNVYtuao4DwfhD0wis3oEO/w0md8jubzvbxD7HTyXm11f1X899LsWlV
B0KgJL3uB3Iv1CgGCZgsKNMG0z2lrQe3VOW8rhulaVgR9RPGReDZbdolqnkA4byI
6FdOg2JF0le1owPdKEs6Ka69j/76rm5qWS+0AJwQzxjhvZ04yDb5+m0GgIf5WiCN
AiqRr4Iwtoij8V73jxoZ1G9V+B5yB9e8NHjPRm/7NQsN40MoAOoZRWAy9q/hB+om
FQV2us1DhlfChRW+sWHcHKghfi0TYXfBzFq0+D8OWkNkEYTP9rGi/4hAxAJLL0oj
s2/ZCvr1iGZx4JF2UymnE++gBY+lT2C+P9ZQSh/fZ5EPeYVtG/5Lq6GtDd3O2XwH
VEoyDKlke67FsoWq0xkRLi+0E+TF94bdh1SH9HYlRAZeTfY7eWRej5nGFvk8iLRC
svv1XJH3r/Y6yMal3rprdL1iD1iPIZ3jgC7mcfSO5MHyE7N9PBHcW54aL3xryKzC
ax10yrHENWlQHD6c5m/Y+r4VP0QTNvPiV2tThU+0qydw7GnwAx6xHtOZXR4sI10J
IrvJqMnKRRRUS6S6tPoD/YSE0XF9RKWhGpyWwW1lkkPSqEvv0j3hLQtXD93ZYiep
2tHBHBYdUW1rJxXSklSS770ZTFO8YusN1PSCLRbp1CxYL4w8teDiQKNK4fhukhGK
/jzcqGVYx3BucEdJfNgPQ39qXyO/PE2wmaW7ppN3tm4diUoyH7HrRt5kEs4TIKf6
tsC3RN0cTct2hQk2o6jhxTTJI2E9Mso9D78cF0ahzF7n/a9AB4orLOyn2jA6bEJg
hjagYV+8JBGlBnHloUm/DZFA5yiN4YDNPrJfrmDIMPF/L9bYDz12OYfBEwSrAlV9
8ZFXiOhNRPAzONGV7sC3u9NAmMeCmOkJ5Bj+79mD5n3L/+YDAT5Q/Hn3ghrXbtX+
kVAaAe3SmITLASdKJdJJzhFD6i1nMFP1X4D6Udoma/+bUZC6RssGmZCm+IRIhJPb
mEiq5sOITRvIJjkczqkW3WeIuwd0skLFVjix4X6TvOu+SKG/X0DhaI/kolT3xEV3
cr8RLTWkmsaLrvAD4ZgcKKCU5DBZ80hQGfYtVbBe2gsen9eV0HoJyrzCnQESS+Qx
37C1Rnt8vCEHRApYERj+N7mlMP/7CWT57anbgnZW40N92xsS2sT5ELoxmB6NyHVR
CUhC7ZIrYFaAuEuOtWB59hKFIZo5vHIjJk0P5cj/B73z2a6um9pte0uHvZacJ5jo
o1yUOIbw7GWIt8P45Upx/rPHsATIZDTfcGjxeWA6w0o/1lQKNM2UTUE36cwx1gNh
UGzHKVvHQ4NdkyAWdjuGUhMXa2nhG5d/yc0t+u+nV/q9fayWZGCFA+tAgYCLue4u
rVS5+PkKC8j303QMA6jRyB1mFDn0F/Bw/WzeDK/nOsgcrWxu0glwhAwuOSxfJzSa
YjrEyab67SxmDU1GBjoyPBKbSqh/54UtkwsSXUsL266/O/W0lFpiiKW34Z73aPK5
Au5ZwI0yJO0u3JGPsA3IHLk1305xJxDK5GaG/F4t9u0hQiPQ3dfDN2rdHClCwyxK
0MXVl7mp8J4s5lrVjdZU9LYfnFtOGYfMaLVZzeGh7JFO87P/AgWH+ymU7ODoQKvj
rwMPNc4A3E9Dio2WyF2wd0/BouFcUtxPwjshbIOSjCvGd2kIEj/wiPHIRBEEyMO4
nL8YsZv118aItTsRlwRBOSUYaNci+8s75VLynsNqlpLjE2ViHvoGuC+gW/3VCFRE
f1P7pSCrHm/jZRM+2hnoqUZk22XUdw8WB3hN0z8WuEiiyJ1aU1Kcrr1M5B6+jjVN
xM8oRIqCoGXM2A0915DIQDkXNtdZze4YGb4Yl37Z/DKFlFap168hGaDQVyoe2QPd
v2bjFAvLD+Flj0qlKMndUe9irP/j9H+rR/Wdw+P8FwZVLgVZqDOdBBNLU0kHIe1j
uUY5s0WLxjY0npu8b9TlP7AYPa+InEivSo/ZIlL8bUJoppqEvcJWgYxIlamympfK
T8ahS28D7u8G76suCaJ4UvRwvyc/LLurgdtzesHfX/YBkU2L5VFtlhdAAvqEnO8I
zRt8EHYWOokzCJsLWFGbYFE33ruHl35RZP5z/yWCZmEcsHwntG8LZyP+X5PGtUYk
3TZea8h0eykpejfKTS3BQKcYw10MV0pG55uEYplNm+SbFVQ3w10FtQpezFsjCQfE
/ZmkftFervGs7egVdJsYSTIJXOxKIEaNVgEAHMyx2l71ZBv++CnGDNOE4HT7Do1L
PG44hzcXoDXLXdR2FKbaR1cNRwEVAjcqo9w3LXjf1f1PBM3R05RGmHUZxO7FXl63
YXF+SPeeibuTGx7Es3PA+X2wcNOdlOPRjiSPUM20l6SGiUyTqDPw8zSubWWioEai
U5BM1LigRT/eiN4xTIl079CRn7sLZN0ZDemJHyxe8OiWID/8muLZpqQUsMGlRaRY
Kkt2p++VJPfrC94Ngh5ah4TlCie3ytZXQmlIxorVdz/ckyGiOIfNGRs/9dubqtK8
/UxGsq1v8FoYW/8VHLtVvcejPzwfnuyYGbtGE04U3OD5VR7riM4DRQpFZUhw1YS2
LpqpJCC8JoBIyKT/gZP8k5X19jBLZjWB4sQm0Ym6xisvPSD+elkuj2OJDMiinoZV
6t35QptCOclVFEpyDp1FMGFvOTpSAb2OJrFm1a4jr5Tp8uDWOhTwLOHjZsbFI8/H
Acmm6dW7dD+xm2zsVNsKdg2t630dx76/3y7lHlZ8zmqOkW3PFErMFP19mJierhSQ
pq/XLQR+2NkIRx+8CPE5j/6cDx/dvwJtCpwO5psTZbz3AOlsVnc5ewmW30l3iI1y
8NxRCosNjCNAC8jiUEsHr1TgIb3MNTGvx1/g9N9FTVyZ4/eIVYdhptEUStip0x92
45gnv3AXH5nJDxOP0PzR1Ao62bsZJu1e0f31kZ0xCWnT6sowDZSL5CJJCzktfHC3
/ORP0KoE5KRcihrp/6VLSYSwxdVA7wG25XX4MlIvZvuwKfxab7hv4PCH425kRvX2
EAm6Z7qqVpUiaBDHkXlAnX/39QDN6buCwUt0yNwwovdjGWNDI6rPRiiLka2wIMQn
L+l8Uw/rQHpp4XIZfGsOM9Uvxn6ajT2aOYtRLWtVKIyCICL79KW4cjNkS7uPwK+F
hho1Ui4PtyKpK0gdaLjtEHL7GS1G9LcotEpCt1aWCumn1nx6LOIai4jDKUSE2WWd
/pEFqShDshvjjvrXlBaac4IClOb7ZTx7b+0+lkbPt2+4ZJQfOTSZZ0kWY4LGY5ip
polsaT2+k6pjZQArsjm7v6quGELKRKjK7CKzE25qDNI9M1VBO0TLFX0RDtdVW/BO
jBnWENw4WkxSV46IqFImcES7cURc77TlA+XVBOb74VqFv+5YD/id3WWbZ/TeoBQY
HIzy5epUSZ4CJUMBH4qaXWS+TYw1FvzMvnBDDUQIs9JvGmn1SecWLC6rYU42aa7n
SGTTCLLVjkquPhydbGlJ2dVKy7JY4m4NloAJUPUdG4IaoukpfjPOfddwIdXcnVkH
bA43vKiI6ip9bVc92FyyEg0euZPXLzzFqDfTPa3ar86Td45usIDWQT+oXj6kyS5T
3AWfG0UPxV/rviFTY0WWpnFIU5VWiTePZWHEQPWslxdukfT7Rzlugw/GesPmlgfT
wRDdQbrL3H8EjY77ETAszAAb9eqoMCHmyhQlt1BRVFC9MdbrFxpD7vx81ionAiVs
LhNmqvFD9uMdAtK8yGvRXScg0jpLwR5xlc07IZ23nu0oSvbdJJ3ZyLN1NFzJ5Y3E
xHaUas08QRBNOimr3RhX/pn8QJ1iGneb7eb9Cvl7kG6RqciCtOTZSLsmkgpYYgiM
ABorOEAmjpKD6RDe0OXZQzvDG+SDvJtoJtVWqyZlv/3clRpogh/oraPRA8aMCxwI
g+BDnuVXDwsWvOFZZqPjcwzl/FfOzX+KjwRkg7BoEZje8f0Bd310KY4BIFEsRwYs
8tp374k5BZi2RnG+UPG+BJwAO9dPUETO2i8fB0aOPJNUF+k5ob9Sy3cahbejzeQr
SE5KG0F1CME5zSTGvBtnbCkFsRJ9KWx1YFj+GDyY7jnBul3vXHyoJ8QovPtfwF7R
OUeo3+Imqtqh6vD0hHd4Yx82hYiaseN+cO9sTEtZC+TbTAVUspYtkhV2+0HNTHqO
iGOdfuRdzzP/cWJMu6T+OGFA0FW6vcMONSbt9tgOOVgEWzAlORvdZ/IxKLj2rPXs
Qlinumr852XmU6oC0DN9xg3wPko3IQx4c7O2Tq+tscBQKoxukPYWpFdz83wpoB9o
uaK0eKTS0TNcigoq5Azp0OEg8PTWCNAKoctqTqRwXGwlIVqPAiSegp13UF1LcrmQ
Y/pcFbNChlBpW/ExhCC8bES31TcP7PCrbrK9KXMaEGFAUHPPsmYXslqL3ZwtGJB2
nwgs/4+TVCntpwxfbLWFr49WGW67ng1uwpBS+03FqwlBWXNlwcp/+34jaKnvCY/1
0/uAJMoPosk3e+OG3E2PrUEle5WYCFVMsMPAGuY0mN9Xm5Zodu4vi37H+FcKxAvz
NyTfe9djgYgu693W/0jCSEDYhwIykdMYNr5GSuaq/D7wBoD18nh1Ku3OAuPrl92A
xAeO2QveCOH2PCHacY+bu+y8BMawvvXnwbgV09639KGTxPM4+XKjepRK0mKbEghG
ReU+hQ0ADxMmvpTGJF8skgTQBDcbx+UKsTF5NN9mcekZ4eNCf3qZci6LCvTeoCm9
Ve2TW+2T+7wcCZE3RyIzN19gW0JTjInk2lrEy6srpEiPalgRTv8rNC3p7oUPsCtP
0BPfwl19S4W0dw0cT4cRiUgKz5adGLhoMrzbhwOOwxXA7IVfQWF8xwJ96zl1wEO1
fipp0QMDrLaUW10RvBlsb/YQjo3rEq3qMdFGo82trKY4+OkNu5z9KRwuzPuKuMmN
8t02yAmza81wrUHutzk1ucr3fHTCpj0n3E1wLc5HcjwWy9R3EumHw1YXy/4Y2aJW
nBWRhaJQoTfyLguNHTBqVROfjMHF7tTojK5q6HUvJ8WtZ1iEyK35fa6jqYmTDw+u
x7bdSAItgu8VLMLWuRlfvUG2SMMBfpTsj46UoFYH+4Zp7B7pMH2z5C3dRM1Dltm/
e0k3O2V8Vyk6ajgAv0ttlculqH2Rv7cjIfzHKMq4q6MoTUQOax3+jLcC2JDqx3eX
AZjvwHu00V7jR0bx4xpXzZcghne/j2nqQJdAWwhaDIEiDXbYjCkPCbL5wN4toDUn
maWJwc7FniQAblY+kz5KZDcHW2NFyr6sBZggws0TSxSV1nmph/soGv5SRQmoiLFv
y9vG1/TDn+ARxNgVxwtjrYmVK2IjTNT1P13fdovXLj0AwWAspBzFOff3tp3CAYrV
PvYln9sqJcAooiAp8pb3fOSDbrUHAflT4RZ6k/7zkZt94bcjfpN3rarLBxZLhIjW
DvCctg3zB6N5Ky5twdVc7NUpZ5hvZsogpzwd9uXGbhicClhjfPV1YjAy1eUleA1u
VcpKmcRyifTwWWv293ZTjOgyyYyviuKKW/0mJAOdhbXabLuSFSSdDsmTu/fAYqLO
1yFp6ymD/zgRBnl8N6of16UoeealtUWx4UpTFAI1o5xRLK4N7bLN29Ywu7dS/XGf
M6WVHbVkjynXbWhCJUmWGDsvsAnuqkfQvgtM4+Iw3Vt79Ltt1tUyIl6FnerQ5REt
DiErZP+ln3qwqALQL6Qm5dRGBJsCAjaTmZ/9LhuMHMIAapXyPiGTF9L9ZreI/R5H
dan9RASpTXPcc2LMuX0oQe3RydLVduzoP7bk3MTHotw4FnPdyTrDDfJDXpN4wOeU
RQDXKIUj5w/yAID0DfOS4Owtw6qWDJg4IEn1S/gALdYl3iNTF00EqEEEVdZvO+lx
vIVOTgIoxUYa5BR+/+39XUo0O0jCXvXOzGxI/g6bS5RbpQv278tKJUmMUGHK7jX9
6lyKbds6tS/+dEAOy1rmCmJUAhSUXVDGy3aQ+Z09INRveatL9WYfYPp8vR6c5o5F
8Rq/Y34unmnXFfAutGppvtFvUvz80TQt64ntVPa+bEsltEipqoao5TZprGU6w67Q
Aj0i5HkZX5yhFhHzST3xySHgnlhZ1dvhEMvkvCIV0qS/yUn9Yiw1rZU+6yubSLhI
BUfWs3YgoGGS8aq2ytKV5ORKPruzkU8BjgLepJ8v0VgW8M/HjIvR7v6R2CdmcmTB
bSdVsxYqlyvzoxqa2ob2ANnsSagu1xBuUzlpgUNKLxzcnCewDqccfC8kJDdTZws5
rb6Rlx3pAnY+Ezr7whwzBiuThBDZzGgDdaCAZOEUPLsnXzoNYdN3Ou/HjDglY7lH
pDgkgWHFWCUDYYw5hRE/BH0lAtFk5ojypl+yZGbeSPL6hhpzm1T7kDw3E2zEXAnn
yCjpJFOE7MydvBsyw+eReY8bfup3YM53Kr/vWT1IzBlTfyupvMZLU0gxMMth5+Bl
sxzslaqzGYPO4I0VHsjcGXDjXxwiUYaDfR/C07411i4kpbnOuwKmuKm4hTNA7W7y
TvyG8PWQ9V5hqzdMeXKrz3Jk+l1c1NozlCrZDkxoITLIHVNMgYzGifMl5la03QeC
muVYYiTxX+Lu1baN5UfJkyYl8wblAeh/XCikBTXy3ww6cQLd6HWrw37nz9e95Tmk
FmHab8vSt9Mhsq9f1ox3w8e7nG4tLtOgRbbfMsngC3VdCz9OoPdN6PNOVWLX1wLN
Zr9FcOGVLLqcGGEcYKE21JWlxT1aX7L9/MuqgcBIlRjLNCv8nZniESJMgYOgCM6l
xWX55LEUUcX1/IbkBodcVFqM7mXOGJjTMO6KBCA5LE2Rkk+QpsfCioJPA+e8J/o2
Ab1sJOQ2B/EAe8t7m0e0wsK/L3Vu6lUu2SzXgU/STH9SI9v6I5i1u3uxDYqKzmp6
4UI77wgceqWrTvc3rQuF2+qr62+FQzH7skhpHZaRcskF4Gjgk+mjcd3sZwNTIWNw
q4PebJxgV0OB4MR7u8bBDxmZKnYlquZndv3Th7d82AWt34SjvC/764XIYGsw++SS
/KYLOcqZCNfIvDLI8yP3csDwQIzJ34YS1iidQpPkPbw9lAIFZFbPFSH+EBItu4qu
4BpLqylfCSGaJjZN63581hu3wUPCSTHxpcsug1yCm8qKXRfK/383Ss67MrXjLRyS
CURQ45Fg/8rLpBpb8VOe7jejYfBO4va6Ovf+RUBmzMQ8VJWMTlE3YFDwONmXLh/6
WDgb9oHRGHH1fs7VSDg/9PqkZcKgX8f9i8TFDGDSfiADnTfixBBJxzTERrFzHcAi
93XaGZyaoRBNv5x+xJwC2ckGkTJc4tWey20YgcGgZpgQAwRsUjdSHOb6EnrQ7MA7
m1qVqqqH8bwBJqpMpKrpjghi0EPtnX9stgUFtvQoaynfFzNfk5tzynaVboslZC3E
sDFszf1XEljcys5X0iwakaZQxBxnyF4a8Myw+QEZogI0mD4v3USHxFsDCL50n7a9
1jRn/ITZznr6lE9yidYINswXeshViibEH2Yryn8ssQvcg3P2Zd/UPVK52Cjy7x/q
Cb14DvUllNzaC9kv26oiCYTxv2uMx55DAlkxoMQfLdxHQjdAGYpo/l8T5Yl061Qp
v505ffwdzb+YSN22iT2VcJSgosVFd6qXdgL/R3EXImjraXSggK1Dc+wjd3BhSama
79cT0PEVM7+v3gi7XpGgl/oaQvO1ZUPLod9gLU8alEtjQT7hu9b5kOwbDk0IROjx
H0cTauQQA0FQLI5gXGpZIxzvNU3208e29EbjEGZlCC1bp2N/q7mjVr90qRHx4tqT
L47/BLn7hVyhCVCR23w45wh6/zoAKUDX/FFL4GOTXoXnnHNpBx3cTQ/ON0O/1eDz
jadiuQer2wODcvaWobtAaPNDgZivzcPUJzrSNjXjjBLMYzU1vTgGM+zCDVng/1eK
pQmvGESkRivwUFNV2y+2tHVoGPwoRkfQiO2mo73RKeBY4j0ge/1RzvHEozEXeInp
37S1+AexMUIUgV5gXF4d6F2Odmw86ZlTF75Y7j+An0pYVIoX4+bBpQBnS4+RAv0l
+laPebifciO6jpFoTkFyUqxmQNk6+fwNKgsd32+fBpgetecmmKqiTmexiNw+IE6u
ZhxGWhmJ9OPebSuqV1rpRqg5ktT+428DUcSwqPvg1b7ZbylEUiqeTfcN3tRikfU0
6kOxOyud458F22Gwym5/eVU+UcCuZUd+2KWDykCgzgKbQYSiSYpO4EKVBxm42fQz
GkL/34+vHl3E8H145xJ+MlEOChtxbSeFDwJR3bm2eZJlR5HYSPPJsCBSRo7U8GpK
vj2lFZTmyo11B7DbsmzVlFbkXrx3nODnLPyxhlZublz42qbZIPBKsKWmoD4j1XLF
pZ/R2nYR8aoFBnL4imCokepGEZEbAtJCQPNoVYcRZecpX0BriVrTXVId37EdNiXn
sz7wEZmBziCJn5jbPR34kJXI4g3np554Y2wuKcrIAKyWN0vPCvaoJ3V6fe0HdLWD
d8uCWzkRKKbbw6ALG4+GXAVSDmCNIm3W+mBBFTUJsf/zqBfHTvXiFL3tITHiTFrU
XuUBNaI1K91KT+5Ntn6TShGBNRbNPpRqUQEWpW3HjTSfmdqsGsg+MzKE1DZk7m7e
NnSCRV68hr1DH4w22P2rUgYXKI7BaZ6zKft03GB6mudjRSLII2r/KSx9lyCmJal/
WclBMmTSvDoSpJ3QEi/ILjFMHmOGs1tfESvSUHMEBOJzD12r3rN8lPUMNM5Sm1r0
/aTHa41R4Vgdk564vxyo5cRn38gAA2yNUsR8Uryh0SCt7uKDDlKg3k/Q9HfiADES
m0IwYX3btwFL0PRNH4SWqG7pG8VRj5j0KVRlr/VY3Di1gcbZz8amW2hVH9kFrr5E
5Ki+zLOjRCyaU2nBiVkaQOOwPoD/vl9UO0zn4zWeOz//iVsKdqoS/9Ep/jRw9VpU
MHGlI6xm5RBqV3w1Sui4K3kUW+u8gh02JRW5gRO6o/5+aHsACaKBLkDjlXhhs7Ox
N5wekvpLEjKsvP6qCMWPH4kWVD6YhAEYyENEzz5ZeBLzOu/FSeDFHB0Ndm/Wqw1e
BcuIK+LyKYpXCx6cl3ntVnz/NrxO9kLWjl4E+NGitwp8OfKm6+idLAQWqPqCg0FA
x5za9p3hSZxzndxQG6JR1GPrg2oi2RXrbWq+HkLFJHg/VbpgoiY2uf/hVusPQuV+
2BM2nJ4iVkUlkujK2MUoL7n4OlR6ygSVsXPBKUnQJZbem96UMil519lO3BxZHo+I
yr3JhWrz94a9tWwcueHTULGlJKkUVp0ngpjc/xzCfkUW+vvyHTYYq3s37Ppcm18y
WHHxiFhGBvty0CLPOayC7Z5HEbIE/VVW/rSny6F0pjwti9fsYNiL8zQ++cBxKus4
fy4dZlRbD678K7IOoq4H+brRI8Xy5WF2nuBqrBUTOaDYnD+bneappFzF8su/GVoE
NXT08/LF2QZhGR2qJNYBbFMBUdzgUx5FC3HyVJAaVQL2yc0dbESJxMOKNd2LG1/m
9H8eH8K3pM2P8Hb0PGo0E0X61SkUGFBaWFmnG+PVMklUaNQx7C/fXnqTdumRfexN
hSkW9PG5T7qjxwy/3RC7rhSsCZp8g4KapkcC3mOAxsza2g0FPBOMNinS2oWQ5dMY
ZAYTapupyejxzIYHkD55E8Ifkzls2FHcCVDxodhiEtes9gBLJgUqjMxDmZAMd+8M
E4o7bhuJaPgiFJCpPEOalo+mtZS0ai9ywTKV3wjtjqZSYPJ6UZnwZrCkS8HHPndm
K2fmBQdMnxJho7Yiju7qnWwjxEag9YaLngND9PqA1Ue22LIVv6w5Vcxl1+VmvIGC
9gPsodl/ArXOAix6g83JjBHtSAhIm3AKC+Rk7Nsd0MSFLrEAJWffhdgSACOeRbX6
V2HHB2fNGTKUNdQTA5tbidmL25x2HK12BsnJkTaLOSpIZ1XqctVnAXAcnFw3Ay66
uOLR+WOIgK0IgcNJ9GRqc978Ddb+RI5lZ47NbmYTa1Wjw6DtKAQQ01rFYSSs/GQr
N9jW+fqt2hMogITOrYKoOVTnITi6XvDaUOkqAK+jZtdL4iCN7wFrtVaTWATWDWNX
+5jT7h4BnKHCa13wq60gl3+MU0iKoGDYLR6pTviGjCZLMszmboDASqusCiq4nnja
jRAuJZXYirfqH1F3fGQlhHroW+5NVb0XpBcqqaB46iWhyjGcrXUG8HrJXPmycB1W
Ipl9yUHNAVOKIrTcvlqvvQJtf+j67WLPCATAO1kv/peCzb5MsxKDvYxpN4AujcEw
moJCgNioTk77G+mn8Bpqs/Z78XRCN297D9BPsFb4+5bezJv4eqdr7ImQPoH5nOo+
3zjngUjxtMxlppePdx3xoUs8RDXZoWXnCg6kPm8SnPs2c8X3TmKvWl93Ry4CPsUb
g3oxDW67v9JxU8n/Uf2xr20JA/MYkovRSxCy8VVqQk2ciGNx7KkfHxW2p8RLfpT1
UzagF/QWK/dGuArN2Umm1txTtPPLgUB/SnQQH63chsUiFrFQqqunNLKYiKwmKcBf
+fF10xkXskE5JuhJhJPmZ1lMUFSbtEK1kcJ6HkwYryOgZKvWcgcl3ebIH2n9jLKU
XmT4deZKHg/dL+L8qx9tLoCxiaQHWf+dncPaaGSluwPkPXd3tz9dzXUYlb7WPuFB
F8EPjYLwrxNFLwyTf2xMXxFl831ByR6m1SXo32cVcH2DtcTySlgV7ZEMuseTFFAn
SwTHjPae6TiiGvb9hsrx4XEr2hEuDyf9MfwtQcBJ/CzYiuidZcG0Sj3zifFufFYR
DhW7CClJHRnfXc6UdNBKoaWmJqDvTnrPzY/kEboqcEXKc12udz/9wgTWGEO4mK3g
VwhpqZ/1azdiyGXP10+Sf+XRpkMNFcyqEeKRRn60jDChI3k3dSk/o/egtsJlE1kb
IZLDs1R2S6/8btPPKQagk1bN9AJuDcBGsUYLZhPSskAEj6Dtws53/SrNKPlIsTSp
F2PlnfvNpPdHe47PswNYuWZTrxN+xsZYGqAnK1nzuD7Eif19vKhDNiUyToQbnGjK
Yol4NNyBuEtmiEXMU6vLZp1YjitZMRdD/uNcZsX1EwgG11XiZTIUuGgpa3WiYMPS
qsrHLekjzg0djPYNnfUKzHRnu1eoX7lJsV54Y4yLQGhRbLFJE5dZnhO5v+uaqf2A
m0B/Mft9lm9fz+TSGNW3tDZFALafOROE/+y4HyFzgP7LLiewaN+EdsLa4dLzJmqA
cIu1TAsahtFmp8UK35uc3d6C8QHHj7fR1ZXvcF7HnuRcI9QWKe/3rBwrbDBUABuo
kwp2ARwg6eCqGRtowo/IR5k/yS/ZyHF6DyT1xezpngDIOQ2jiu1N+vE03WW4nBGA
Vd5fVw4rDBXJqqXadWCn+CGc6Qo51LR2Fcf6zunxfXzoNZEGaep5l79XwMBDOS78
mcHvfUBj4rkJxCWSXNIoi+Rb9KD1OFCK54dCAlL8ZsMgrYuwjywqmX5PTenQNfjB
9LUnL3hG3mTZO7IHkxVSyhbv2lK3quU4hgtsZdVxoNMoQRPI2IU/RmXMeXFzh7bO
WriBRYDbAYuLR6i+Vde/iyup9kqNVT5vwFuKqmfvcikvVl52wPzWFAiuTVk/hnZZ
jUqsSArBxkYs4Vd0lxP1KyEGfTxTYLomVqbSG3Lwms7yJpNkLBXBhZyklO276H7t
E1UT75BPafkHJ7dN5B/ZFoaElXl5YcGfUYgB9U8RU6PDpiHsCZeeobHHZjW4OdM0
9/AI3StTuTjlii/tYeC8PtrWEt1Pz1Et8/5LX/L4yKVxdhGV1DL8T1whGAQUY/cu
ZNA3prYnF9MqMHsXcz/lAbI9ZbHfERz6FBwp1fXew5AYdB3061VEF/sv4HdY51Zv
gTXQ1UmnQy2U2/X/Df7dubrPH0i38JVEdud5LN4ZRcsXN62WhOkv5MofUqFTF3l+
X2gd0D2Qz11MsSKkyF/aomYPhJq/jkYALLs8IMFHetlz7RujzbUWl0PmH7VeX16X
8MQQwYQflRy5Nb9wqEkIAWlZms07LCoUL85v/o+wdaYT3Qqz4viP/8X5il9SfVGW
AXEDRSfYKOWvIRVvP1IeVQLw0J8Ln8AzIhLeSW8UVCf+ztsbWWgTeWjaePbjZZrR
mwjy/b5/YSW69BGhPcDXzDlIZJ0P7fWs7GIeq5EkfbNmJzn3ki4IKdQtQkQvQEX/
owUHqRNs0SOYi0bV0L6jB0H2xvi7nF84BpiQXkA9zdJxqm3nkrvz8Acaxkq/r7hk
nnyQN4DfYpxuDBdgbBNLmMPZre36eJbskyYcnsVsASwsd72PMtiYoQxB9lD2aKxd
hayIZm56bwgl2UXWEIFLxEUh2JgaLx8DZfJY7mPnhulnqDjQL6skJqjEGy+WcXhe
h66jCVQh7jlgrDznQ/UQuWpN7rA3U7LCiUxdBi16VNu3zG1wXt1/iypFv7Hevsjx
Swh3nHi2t9M7SpqQ+mStIaDEuoIHuUh0Yau7122U8xOzknaQAq08hc/VQa9E/MTU
0gsS5Smlw5ABgLbtjFQKogfDItZlwBOewBPkixVF4e8SiY3s0H41oKcrGbwuwYLa
4F4gJhJ9VNkFQx+Lz0MQAoOQ58Mq9HUlehnh9cot3S2HPtXCsX9fu9EgPJsSIO5N
4P2H9Z+CVil0mIKTPlH4LDdRbaX6g60eBmzM0qtNhPmRGP/x3Ps/3ZNpwREblHI3
MiCM/TsIwcTRPE/hn+sFbIF+QREjrxPo8j1iW3goE3MrGLeiZbi8OcgU6Iig10pa
dNx0sBrW1Z0gT1SLWDCBXwtTGpaFONEvQzFLtWsGaKDrqUieBG58V0dco8zbFpRA
S4AXjiSEVI/sXTPwboR0AhYdrIKmRAEuwuyeCSWrpmy6/4d6lD6sGDLxG1HQZ+Ms
j6DjFYRKvG6/7C6YWzzFYPOTxyZo7rrYUIIwFaY9NUahR6w5M5UQy6oiNFYOPydW
fj89z8fF4SmWVPX1ZdXJ8ZxNpQhB+5VZ0nOJLb8nmglpS+LqG7iFTbzO0IXZibpT
cYuBmzyyyRgckSI/+QE3LqwszX3oeT1x1wNHwsyXFamRb4shkhO/hdXx5Cv7vhoa
vlBmZCV/jLYVwyt1jFVqUL3VSJ0Kmq9gPYv/0AwU9qYAKgpGvpVEgA9rjwfwFG+d
xgDeFvjG7D1z+YGPsUV8oDDDmS+WmPdn1/EZU/trE0rgbC4+yUV5HsaChyiDLw5q
8IAL6WVf6czWvs1k964PIIODeUePOPyBNvEq2wo+ebQLhwnewEa98G1irFzA5JXb
PXc0IMY58I5nzLR1f7X6uKj0zerwVfpIpQGjvga+3kRgdg5SqEIrBoUoCAZsctSe
KS0Yfwrslu6JpsI6UxBhH2Vcm0qiS2fCCSQiPBcFgNocGi2iT9ZR3uLVaDp4tRSb
q6iLmEgrdJf9VYtnToCxrFZP9dLXPqHPmORfIyPhRPiEPG7MaOUaOARzo3um3HYh
m3dCpOdOwGlwocir5avl5q1/aD2F8gNCNRpR9n5c5ZuEvj57Ms2kctsLVdsJX0+2
FjhW6PGslt5TWFOqIACpdWD+eQMmvjqy/X7DmCGUyQJQ2mNTbDj8tlna7usAUqMy
sRodSIW+6BO+bHMGld4jc4rGN8wUm7UnvAIriBSTuVbphOsoMLQ5wDlO6D5m+jAL
yPh9uL5se5S8XVBLhX4mLaaomT8pq+yEmnFvh+ky64qHkEkEnxHum6lhJoFeOPtc
8iebMav8VMkyqJ2UftUa3vHyQb8WQiIMqtI9YYnz2Gnf5/Q0X1r3Qz3gXRKWZ7HK
BsPF2Vvq88aM3CBMPOxTSi37VazNjKPNx7jLSTU542m2r895feKlEymFhkrdM9om
Qm7KfOCVVoOxwjU5bIFRiulEA3DCsrbSdrgqsSnQExm/o5lj9a4F409VISOi6CRi
SeANORhGEAXVc/gk2iycjLOIHyijm+xdIpbmx2T5ln9uFOHBMYlYslQ2d8gCRVYb
KPT5TcM4fwhCf46F8CBCQDSin0QakcWDbNh92GqC6IJVTbqicHFcH8wiiZEi6o8C
G/MwG7PxeMNWtLSfPY6GF1axLFfGxKeSJxSmJuXm0y4HzVpZDjriKe3CCud0MGlz
5bgeWOXxLb5qlAFhLeL1f93dQgV35RDkcXhbkaeN335f8swEOrMOOqzPx1imfn9M
0Est8/fc+p3EbKTVkpzCo+F9oNLGB1m7ihYKQkfN+WcDjtY4V8C4/fZA0GNMqchd
yw1GAp16VVxthN4UwGalNVFWN2rPRAE4JblAy+YVkHsxuQR4+Qu8wfyc7V7K2fFU
Usx2NaVNEsPg7/ye1JucaONChEoqEmL3hvSqpEjwxk1Fuf8ZC3CUWcMt1rb3xrtd
zBgtF5q0C98vGc6J0+EFiwkEzOiOzgt+kUuSvBBklFiNzGyViIwy+IqJCWHI9lEy
s4NguTZMFf28TVlCKg0XsVJ4D4N3bbsbz3HDAtgMt/pCgZ18wSVo6Esx8Nkk3oF6
NUEZtJt5OsF+1EcK88DjQ56KfOHCTY1HrvQ4TP2vAd3lfqdOyer6c9Z5Yz368xVb
qo76nO66eN96sFy49dLQQCRKmOHF10NF7G3lbLQdrNvVcrDeXlnl73RIh/Ez3JLV
lvnOLQBpTpSI4wfqOOXw5g1zFWZcyyorCcBdk/JnNN8axDrHOz3fRtJ/cswUkV0D
q8TJu0sw6abopFisrkp7CjUMNjD0Leq0mVHHVz5TeGr6wdMRfa0nZqS7YL9UKrxL
UfWauu3FOTe544ugM2RxK7x8lE9Ks044PV/X1hLT1reARU0tmB9ESDf+UJvE6LtF
J3qfTkKWCTRiMhQ4wUCXYTKVk6BFyZ3mXTCad1kee2MQai69W29mAqW3DZSZjE/M
/GoBw2+oh0HlRR83dIBXf8AsqkGGdWLZDgHpe9B3dVUsVBOvsdz0GNcPvJHbfe+z
psG/SipWxOWdcj+7rPoGa2tyZ7slRffgd9fBp2YehTil4OsapTFV2KCZ6gLayIox
dufBfV9hsyUql/+AR3XRFoG51J/zQdK3ejYI67G9IHR0JEle4UT+FIJUHFmFVoUM
ckryjQbb9vDSemW5EdpK5V4bLdMyiHytLHJxi83HmzyhyRmP7nOZFj997hmytfQs
/Dlx/2mOvKDyebijUqlIRBMIjV2Wqeco5LezAuVT4v6LgA2kH8epabp1dUGEFuRw
bOA7dI29ud9JzM54Isx/6CgL3D95ZRNUR4YSjoE4cCfasu0WJ8vKmn7kXAvfLeWe
s4teCUmkeJI49hmPEq0Pulltw9rk5gFEzzlqF/kB6AzhjD1lICOwccUvYuc34rzY
jagD7edm5ecHsi9Tz+V7d91gnVhJWWkFhUk6ptc/l+/tcLUpcqyhKVQcTNzQFvW6
Za+yWbqyZ8NfOAk5Ja9xfDYT1Uzw7RTJaUEplUZEs+IWT+GzUO7wi6mySxl7GKkg
sTy456YGJbxxHpWx3hHITYsNass66zcJAQNbmY7Dcw7fgdO5XgdRQ4XwzEGBwcVc
uwetuTsYyy3EXEoTtbE0SCyQ2xcTe1m0U43QENqKJ2kuR0y+gCZ0qqoFWCm3FHZU
L8k/tZOLsd1hC9gHgQ5cE3+KBdpDzRvF51JFDImEoen/qDhcjIG5391k6S0NNluf
gIlOFmHiSTklB1NTC8GczFDS1s0li6dDzfyyPCw6WYAOqDjS/YpRRaKmji0EKkmi
PnvXLykH2VdhdCJKJKDAWSotX8PZAD8k3DZ/fJQ/2/uflzRCGZX+EvRhyZlLsznA
GG4KBuzSNWNw2RDGUFUpAc00HXxKnuh90DqaDpOfWlBdG/KxRZfyGQSZEBY07Q0Z
GsYoWsUUoiL3NON95kwLw8uRlzLMu4ackGr5eaK+QKg6vX7Km97Ndu5f4q7JcGAr
ty++7pkt/BDgTVIqpXy1GdDiqidPAglpLdFd6Szy+EBotlSPPRidKLNofhilBBQN
LFyFfT6pWKYM8L2JJwT128Q4U+GbIcyEnZLDl9ATZVSweBYOm+zhvUwfvbzPWItg
kPbT3esNMfX92JAuPZQZMMf4qE/vdZ0EE9HxRbPwQ/iS7OSV4ay3tckrUqO9Pzyp
xU1ptl8jlJGgqNJnW/iyiIWWeO7/lI5tVFOftpBfOHYWGpZ4ulgqiIswqCyVQCrY
8jnQnrpa3J9SgG73W55ipyqORjK0AA5xu/idXNdNGtbnuag3OezDvqwjTQW2O7Ty
SSWUCgVDR25m0hrbFGqg/rq6iZrMkS8CqDNGeCn9zgifa1zE/rr5qdWKCgbk/1q0
hcq0JAqMQHeXEqmxJTplLb1NOVmCikbFHHJb+VFj4QKd5j6zo0rE35ltq+w3vfoh
kwfxsmi3T+GITEmLXZRTiW7ex+eqElbLeyXWE83QaF5fhZDjOpi0xgu5J9lFBMR1
+ljRijbcl4/yCS9n3Tya8cjoW2byhpucXPi7TTgD+FAW5U5+Y7bAlEI9jCmgYUMV
7ib8y+hN6+utDhxMEI84vRCiBRuJAO2lvUYw/0bN348Yhlu4cxSaFKloWzWL6AnP
HilDV1wVpk37vAuqzby9g201ovqteof/h+523auf+os6jQhAjy7HsRXugwzM4Ovd
xCNCNYawrInNXCkto64UwG8U6Llsbzmd/H3LkjXqdaCCoP5kfk+YfmrgVwG5CskN
R9dE9UNiuBev25cxG2HOmmY4dDNB7Y0dbUqYP75kiH9DTmEQaj7KaW7+E9lpsTok
iizo2qnEcNwcHZ4DeJcHTo3fV07LQF+TJWotJ3DnGgB591PUvxlclQky68+eA7fq
oQp7UyVLzPjuZSH7FKpPekAW7QgFCOM904krR0ZOJ6Vk2ouMh1oaa/h8rroEWSD4
4b1uUF9MtfH44oiiqs4q4Jb0sA+89i6ffy3X2DQA/rbOQtdGrkrJ8A8+7nlpDQMg
McD+OA0tU3qq38tvSeI4m0J92uAoQgFZcNyZOJUz9SHMKpkxO53nCFaTGjW+nJe/
uJsGW5TgJ/WvKLb9WK5AITgfYRPRA3+C1sASwzCJbK17JabwkY4RBfuD0camsShu
ilqb9N9+Db41ir3MHmxrua+0u+4HOKHi7mV7Yq4O90XhpYb0Fuc5HIjs5bmYrIhb
dAT/l15hk6Lurj2KRIC84ma8FOLovFGMrB47e+CvPWY8QzJ7lXNeSWLGWVKJz7qj
pwvNEK3MnFgO75QeIXY0PX9fFi4rhdNVFYRDdMXPOjIQhgbnJri7P3Oa9otK88dc
NgBz+pg7e74McAwqIPjP3oswXmTCVirm/twzjo4U4qhuYC7YwEbb7J/PwSitnp8C
Xvjd/gWRVeZmGljOFj5nZBfVrlUx3GeXuB043M76GlpKj1ZOsPR3STu9wSWu/ByM
IiKnPxxieWY4llDxh6BXjng92d/iq76x94QmBxHUUUS3u7xxR/HTKOVFOl8oZO9O
g+qQRFQy43OSR2WX/mztZAdqOSQwDmpSjfKy64osf3T9XiNvxdRtei4czpjnSCdg
qfgiqeSX/AA7dRtX1k7f6HYuF1C1jdQVwUx0d94uDnlBKGkySP761np6n2gVeo+e
B+AiOtK9Gsl0TeRYbom4wxr8P62deQ0Ghhk4yJgWjCsQLqfjJTKVK770MhKb6Ngy
FmW1n8qLijvSHSLI7L9ENH5TMOIMILei8I15cZFyU7nZFqz0sqv+K4afOnAXrc/4
d49uUgH1CVLLFu5u/LhRdtw/pYxnPHr1ZeQN3CM0NaBCGPG9rwZ5gLckA1fsdzzH
3ZZcKRcLe/kTpXeQO0HCpaZjP0NX/8/MTc0PQDll1Zi7h2vjIQ69v5Pe6YvONn4X
i78Z6pOWpVk34CA/f2F0XvOiMKJtl8I0VkEvJkp5DNCeVWtcsWph0Uh4lmT/yzvD
a76KBxJAX80J0S6iLh2SDr2EihDJwH93TWlmInU6j3A+fcAnGft2UU8Jyn8s8ZFv
2wNitUjQAi+Ctl69SsQ1ZKk7HlzyqPpc19W2RKOMkVTPAXeVzFi30unIKqFtH2NJ
0ZHxGifK7lyqkR9fi4onNHmbBOfUrrcDyxv2IkYrZzP8sU6TxeNRvFXC4K9qxwJU
62ajnC+9Eq04wDAj5IjkHDHVd0aR+1tnm9V0/nnq/SJWTQNdG2azqcAbcaZfqtmd
Y708NgDmNcsODBEIYy7bVZRgF0sVpmk47cW2xph01P1ShSURLbrcmNSPyhvGwvgT
qetBWV9nXHkQf8akDs18t5XLqOYuKzEgNj3mTKuRC4S6EUExOTx6SLqqYETT22/I
S69aj0bFYGisemIZYElaiZ9Dcr5v7Hle4mxM2a8JdATrNaKBJaSL1kI0Ev5Z6W7X
tKDZV0ZyyYpzEZzlhn1rLVaiHBmSGjJIMfGMK0kC4IpQwNBMG1F7qKVLRekuSG81
WIAlKkvZe2dVJA2uS2Ui2pg89thZjjb+N/cxr+tiLlU0eO9CsLp39vai2YYP4ng6
4IhgENg3sjGppjX6/CChHhWsCXWLDEQyciafVKBYaR+l8mAtAUS4Pw6fgTKW9rPD
TK5B7xE3e6HhQx2r6FceigAeyAZ/s/vvvZHue9J7+402l+zFIcRhbTYeGf3FYdoY
8y+9t8aYtxDHs+2kcknOsHmH+ahLEFeDqHHee4zSWQzCAX0jH4nTJ6DRBF3DE7xy
9mtyHtzaVaTjB/LmD7+pcY5OzWQ/ShaYObiMcyNez+aI8jS5z2eKJlvYUPGxG67v
Bd/rb0NhbFBAhkiUF/BUo5f2A/r36ATDOiq4M4ULjAiJiiIoVO8dDxPrfgfYZJR0
TdMd8iE8tO9ZXcjWifdI2VxjjOpx8aKeFUYEBkU3rPgOvnyqYLqnckSwQvkV3EvI
dCOvmFAcOuG8ae4L8F/P+pqaL6XTN6mIUo1sJvTwytMqN602RU/MjzEpjAXa2G2r
PMa2oPI7zHgHVjNAvoxCftPInYc2/hq8e6HU9hwZyzAIcPtv2L5xwi1SFL3MONRn
+AiCVWAsqE9SN9QR7rluMvMh8ZM7ZaEapjg1yeCenG0V/j3+ETVWh49cm8T9BIoz
AMPS4sYaB7vjVzsEN5ZlNQZXyJgG+fS+imNqnXkI8ZxfLOUY4Lxu+17Za4gT/4lQ
aGnwSfLithCM3jM/Y8L8jcX4K2rDetdkOHVPjB/KzH/4uW4fbCpzJm9WTwsXvY/v
DkyR65xbj54I/a30aeMSLsGmyn/h+WCBCi983Hy/Ov6x5t54A3pPP/UzYSz1MUqY
LE8dg9qM4iW8MQv4LugdK4VStEcVrxcwRYrv0ITnM8NbP9rOh1ups1cScaRDulWm
SkeS4NHrJMjeQn5WWhma94rru33BpReeuipdFvgL5rA+QN9eDDBIKm+xQUKxNmIZ
NNVTAEnIClWWh3K/D6EXO0USCFObx4pDC9Sr5GU+8suyEMHTYWNNpB3ICSMqN47v
+0kw83zpHm5ebEnJo6miqUblpGDFBvuiTunv1SLBD+LnmJHw7o3Zq9zcfz1OBrqu
yUYmo/OXpETORZHsvFEn/nHgjQIeQR9peCJBQo8sgbTTsotipmlO/GYz6uaM7r0D
jVksjDEtwQkNTfmMT8rhphvzXOyY6zf1Qa701oit+j8xYBu2eKmTNgTn1abGgTFb
iBR/Z2bV9J/kj/djnPnpBvZDWeLRSMjQhJIjg3Ik6f+o9iDqKxFiPBgPVY0q28vg
0ddz1Q4YxlNozgsxaf6kTn2xGoXEB5lWUQDzNJJ81wKk04Yx+56TH64EP16sLMkU
un8H/jIc8cQK4QwrZWxbyoVWakoEZrCSqlEGEfRVkNGvIXlkWNRFRHbS7mxa0Wrt
OQTjKSk6UCh2xxryv22eBvtVHI7TsiUFMl73ZqtiPJvvc2OjNGXRqbNv1mNSjgrU
JrQb5/mImDXsqZwtDG9197chIoAMnLIfITqARK2vu7BcIp0ROpGNWbKFu4v90M/S
T4+EAIsOLm3H7b+NbF7DY+3dh/6/DGbW8DyhIzeqFs5aU/MFCFkG6mNoYIOSnT2B
eO3pMenYCv5guvb08taTNS9z3Jl8Q4b/Vc2ZRoaWApNi/6GWgqzUT/b9siTmHcdh
pJTcbyN7KSmOmyt2WyDSVGkaMhEa2OembeHecaDwnAxZTzJPt4icZZ4EOIMFZW/f
JmK4b9ALZ3nNITs8oUjatI20y1HVLBvRkF9ZLZ/bUHkFbsF71+maHVgqHP2U1Ba/
xMnItLo+DqQQrf3hyPuGBHiWOfEUphcCVdTeG9CJDHDiESN0mShRFNIuEhTYD1X4
B4+SlbZ97rFFKmoiVUfnKnURLZRlhHZgd/bSebBsJXe9o3KpJPcLt7SBAoy8bs7i
l3ute2/9K8EdxIiNxFYv7hQMJWwR/gm9QyDbgzUiCWGZGcR+yHfQx3UyzNZTECLu
h/SAX/888LG9l4V/f1bVF2+lSYbOiQzk7xFwEH2uSkupCAtknnv7vVDgC+HPKhOr
zfoDkBwAGaHVELBOUuRM65f8hbwUUjCWRGIBC5M91BvwGJNF/XwRbB6Hqs97GMWk
esQqbtC8V2fzcQqRpedeK+lH6UEXYtpYuVtoAzBabmg00Zq0d3qqnfup13iRcwfk
VljFZ/sOBJ6Fmstz0b6s+eZ09nSvl1eCB3+ehDor+ySp8XEvD338comyOl2FZUsX
3kN1VzwRsE3jCpZBQTpe98icft9q1PXrAGLog6Z6wCotmDt9daq5DAG2wpIlL1fb
R6dFOp4KLzKRe4wqAr+qUTA6oJCAg4mLMjM0qIYK7eTd3G5B1xyGdxfpyQIKLikl
cikOccJsMaKJ/ZBiNsL04iaE6mEtnP7C7mi0MMIE4KwcbRBEOXLMXRN5AkNR6I6s
kVgOJxxoyNLAcEW3/w+6a/leQERkX04HGjLQrdQD0+T6JmHfwIdt7+s1+FA3B+s7
VlhuXyO7egb6iSKzzQoiFnvVppm4zxYMk54dtCfyObyZ5gPelS0/6uSoDgP2yjkL
8lAtgCNKV+CZls7WHO3v0noQtxYJfcQ7Vz9GtdwIx/ZlOGGKQz+15IFrlz4FpjQn
4/xcSpq/LtHGgqtNXjYPPRBd9IW0qb/IiPW6nW7prnpOqmRNVG1ZvIMpP8rklguE
DjjX32V5GCZj/U25SIBo2NoeL08X+4MuWSbS3AA8jU8larj56PnEoUT1Wa9QXA/r
OZZkS51r8TAQEMtUn8QnONLGI8S8xRn9WEFTnd/AWEOYVR9467lLbWZka5qK6/Zv
wL0it4wvUsEW3oQ9Q7o1NosVlgUOOIiDQ3P3KswG3I6qYyZMhzYXtta7GmEg+LsQ
n/oMHcrb1nOHNiNNYH54tUqpINJJwdF3R8tzR1DcqBPT4Tzg8HbPvdrujI8jOqiw
elb9MP6yGfp5jUK1b/tBDyqFesfFcMeOVWuig41i9OcicdGDDpskFbeLtqAAmDuj
kfZIHxlq6VLNYkOB70JpgmhFeyCmN02ocuCM70WmSi0i32uAuB+yKMXnLU2tbZiX
K5JVy2n1IGpPYiRNNhuOJ7ZBhlRL2Vz+/euOkz1O0V5krqddpplqqLOjy7bkgbgc
a9eCK4TJeT7tDCIm+SLkuSliGuVTr/I+nSM0ufFa86126BSK537fLXLNb/Ok/FZf
F/bumRp25u7N6BYLYAa46NWuUo6AF94tMHifqUH5N2LzcDcLiE9JG/mSQA1kMq0R
T3cY4l+Qp640u8AIWmyJGy3pGwuIW/ko4JshiUG/Inl/9xZhVVxSc5eZtM0URqH9
dZ/yDV2/OvUnJaWzmeEbqfP7VQJejP1x5sN654951vl0JgoHnlIAeZZ0zvhTbCZ7
tMmpHDttjeJLSnsGGsCs2oWiTJjSATvWYKqvqaSt/7io00VIhditiqgLHQdv1lob
gscB+xCpr9YdkiSJyRCmzxMO0HkUP7A2ZnMae3K9cp43Loc0SnhvNQWHcoGwavCl
3pwKovA0rlFWlAuOzACWNOX5C3IuFoPEuXQ9vpEmF3lLS+AC3nrOw1f6wU5YArc4
gSlYmId0zetP2oHhjHzNlYjpQieSHbfzETlHWU1X9giSbFN8fL1KJ1rlQe7Yd1EI
uwzNV57zsH2L93aBCA8Jt/2YPXXJBo4OBfrbppYWReCUQwewRO0EWv6NSO+0nCte
eV5JiVzJogEx0dKtBGwBGhFGcoTDU5YyXs+U2aXkIzgsWwERIDwj5mBdwzSX/dRW
k11xvUTTsX8frwFykzJL5/VD0UnR2z+eCN0v1sm8nMRVvtKu1OHRrJIGcXyxI8cJ
m8IHP2XOXs7bpuJul13oXz/Dj89V3cFQxV32b8z7WcPZKzPlCBzVGHbde4OH55RZ
NCOgNQJROvhlfNygmq/j0EnQ6D54eB3qLjnu4ambm2Q/puV37CsWqG7kXQH1XBph
rdJHDrfiFgqpwRJg9Mm2np+T1U8seiTLScnDywTHPGa1s4zPnSyecUe3wMVwM7Uj
NNl8uK7j5+jzMCxEVpBtqNZhZS0h8rtzPQ7zqSBOH5SE5PheD97y5bDc6hzGNj1T
q8FiIqe9FMxtqtNkjXI+LluFrsznFavMaSg31+rJb85Eq0xmu2Kk0dqXylRo5eAN
rofoiAw+BcF7yL6HpqoiYgjwOspCiCDA/oO2MBveDnGa+m66jlUZKYTS4noIhPoG
L/XxQQSd7NFIbo993g2Jnul21MYoVzJlhfMdxqrCES5uH1gjFwZ1WTriid86lKLQ
Ro/5WvzmE1t5FsCH4kzI023eqghuJuIFdYDdIz+Ejb07Q15WOBvZ7Dt6t0LUnwOR
oCTSPE8ja2Fns2icG79Pc0m4qqsWB62B8M+tMCL+QTFMpKyFfFtlJtxHf2Ilcaz3
iKv5bIx4U/dPKkFRjC2tAos2iDy6buvgJVwJB0NXnR3s+ez3wP3+VOV7/AXdon0f
2SJFuR2L9K/3pX9O1Pfib7qmq2tNssJunhveMR19q9DjpXMlhvWBFLMyTb6r6qWd
RSTwWANyi2hdQwKBFxLzxhGznU/aBNLmtc/qY7aLmnWXBWBP9yWyVpqDNqY2TWSW
Wi4y1rCvcxyY1coOo+qYmT03TL8SP5TmT5DxyTc4cEofScffeFVOgRMgONYI+oZb
B5Y1+iM6nHZd/Jl9w4+Z0Hj/90Wl4EK1LBTBUgtLVfeR7fo8NE5KSfBtEQF8hvaN
1JVyMI/d3Hpxvu9gBmaStJ1fHEJlWIHbRU0uR3SytmH4gnFd2AZsxDquYP5BrzKy
8hS+pn2tEX30/H7RB4sQipz2pjv4D4Cmya4RX84lvJ09U5iCPa2kiu2rYjkCahA+
f/gU/0ekYdKhwUuVBikD0gT0Ef5qsXLj23AIATcw88kSZG29S0cmxborc7/WbtUt
5LX/26grxB5lHqjPVvKb+2rLn/Rc4nx0yCjBF7hY+YVYBROwdcZQRFKzENPvmmxK
1fE+g+jke2KAsYEeGpslcGK2Ba4Mr1JEfwhfQF+EfFYpdJjOLHtSCT3Ipyplc3sr
A2SyaReUV1MQtKpTiq+BBQ7VxcNvS8cCpBbkbplicI6ZWImdzrKHqrjo1oH5RCiB
+4na/cf8K/yNEuKfK1ThURg6JyMUMCOJi0w18onLhzsa1nSSerKegS3rdnOs4xIc
17vxck0dv52Rb1UREm72kM8O3UYg+awjGQXelj3BAev3rFrguJcXiX+kVBjOVyel
isqJIYDwVSOikMKHcOFcdFJfUcSnwEowQ1gAHrAIHDbCRx0mzEahbOlXGaWlmw2V
PVZz2fUfF2gPk4wPlxBJ49NsUQbNh+y4n0NnKem/N8O8beqUxowm8DIgeexXCrZu
2lxJZwywypGs5l1OLrNBjZ52/9CgvLPp54Gjz1l6SKqULxVlor5DJ4wd2RTq68KU
1P4ONbvWhZ+vSZYgORryLcDsyZ6cv6aND6ev0xjH6TP65ynzLJk8BsA31KjFNlSI
FRu6Ck3eVBAtl00Zd8ZG5a2lxs+Ftnkp8dxhYn+eUo3M1TkUhoyBVVNZokl2uZv/
wAlx8Q/DdJdkmUSC2F7pU1vZhzEcaz9+YBCg5/c2027T03CRL7zXiDzmnI6mYNNw
ncf13kkYyDxq/eGI6RkBWzJcLRxZnroafKPyJ1EvJ1vh+RBqPpY3YhgMWBrWk9jc
9tEyGJyQA4lkkLmRAkgalfBwwMOsnvEXxNjvTRI92R23ahHzEIZE2FzlConscwgt
/fx5797qGDulQ7psXGsRd9/KiX69UMrFKCuXJzkqSJSKMMAlgklRTdkMfW49H4dd
AF51FQzYonirFfyGswZkFY5osx7HfdKVsYJr9tyNZ4Xlhdog1z5fQI2dSNKrzCVd
KY4eoMX8mi9UvSlZpEqld1A8brIOGyfLwwxRY1LHTcSRP2kt5n+y6f10TYBxRGEy
ADXYX9cUdpTcjpntXgRqD2bSxJf9k5lSOPCxfjxZjiwq/biv9iwES+ObxKgFhSc7
IIX7codLAnvDOEsA2wgYaVoDu/7kPWv7p5B604ogf0+gDRUfV9fSTZ/TDUqhvBha
LiRJ5hZSn6qrlNp4GkG3Herb+ngG13Or7ifpexOS9iuJbWm0QdSszihyAFv/ca+o
5zUqgzgpdHJK7wPkWy6aWXW1YnFCy7ggeJHPX4tSpomjW0CDhyOj03kCsruz7d9g
eZ1x8+PJdYliPJA+Bo8e4AW8FBUgdypTdUhWrruWak6FajG6qIlbAf7u5MTwGiCb
hNODVzLF0gUeOXaw1UziwZaDddXvodEJUCMF63dEHp1Xyrf95ZjhVCOFnHMpjRom
oANRuGAST7eJoDd43q2Aci51Nv1LP3GkfjIZTNOMmN/buuPE9qkOzGOVXHpoJwLO
epEukz7xpkO6T50GNML4K5Yomj1lyEum111bJUyPxisSCjtgsos7xuGPHU+q03lc
Giyeat4squ8eOPfeQVsmlDpMq6JgWhHWjwKsJ2rCsSqGtRLRVvRTO1m68ajtZngZ
DXg2t6PDyPTCvzcrBjsZSCxMLZN6Klq39lqX7tahDBQxcOUsoQtSnjiyaHsDlczD
278O6fhbk70FfQWSqYpmbYnSjfuAIerAo7KqPt5sRJfuO+MZMtdtWWubtcP5Milk
G84xUwIFUWXONqlPkhHKJkW6w0uk3pW3DT0bz6oSsGgb/n6Gn28PVFyKQ2+eGS2P
CrV/z1y1YS9Fg0Qd4seulRWlRomyodGuZJ4n3ngeoCpwPjF5WTqBMAjBEl5aUKHM
aDOhrwML6It4WFVKaxoqQyBgVEprkMqZdrMuQLREQ+QPQFUSMAF4CpPfuy+cJWxS
oo8ZXYqTLTDWl9aHnan6UUJm0xpsfHQDSzXWowDLQQICRczcmACC3ds6i7As/Kjs
qrLXqNAoPb0RDRSpDWD1kSGNxBP+ADPaZtrfdhKawfessmtgl+iBbn88js7kpgaw
tCPbb2PTBENP+7+NLOGQakCuUs6HUn1DSVqD5q0uxInVU0ZSfR3IoaoVgIgZFNBh
7KY7xaEpuHEKAGr4/sD3H8cpw2WvJvPwjE45bq0CBfVllEA0U7jR2iTHx8vrbw1X
9F1Mt6pUeHSQJH1PoWiV9ILY2OBJU9TV7Q+Bmszl8h5XxBPGqGfW6fbjTrX40t2k
4qiuJ1nQfdrS4knwF3BpNDkJ6LHi7mxHJCXurMixy2zDfhdN5lSyxkQvcUMqJEXa
y1+DQVuSvYuYi8VWXDL2qPZzOaztzhSuFHR5/xolt7HwncoosahVZql558b315Xc
YZUI3TFAFY/9Khm11p14kdUbxu2xYu2F6zOZLVNWrpRjdaT0BJwDVP4kSBc0ktmT
bzse7c2itTFPDpLmEo3FI0G0jgnNrQFwzP3HDONQgNI/hUDJqY1FbkUQocCzwn4U
YrpQzZy3WuW06tTfdjq0ONChw18XZGB5zqN5BrYBeA6NafduJmwlP7nUGLIRGZm0
1S9a/c1PoWR6hvySBpOodlkGkIIOJfk6iZ0U+HR31V3nEbp1qQ3k6FvdCjXAC7h4
/IttFl4ucz50zo7aq2gKpFMCriuhS+DxRphR5Ge+xEZ+jB+qVrbsHf4YvMJDQDCS
YPVQgi7RsWugtKfmUuqa4xju3jXywCD9jHe+zxNJY7WI7j+iN0L3oF3brb6etH9e
YVDVwCyvdLF+L0y85BJ1YsuY4iBpgdcgp61hHU/uuQPGFaDkNE83e4sLy1Aiay6r
mcANBVePeXAeTNJFu2+/Swpw1QLtGsfoAto7iPd8+1KypY5xd36D85k8AsEc6ff3
MRAzzTWMSlzvoYtOXoNImMgmrScdY51CU0PrjyWtRxFE0/7qr3LveMHD8xw9wA8x
TbKgZ3wM2RqreIsnLUnhzZ1ZZvb+qfLMKC2D6153Aheu5Nu1qiyKXR606sPLvbEv
HsZ0v/CsjkI6OPtSp2PwV3HZS98VK+utKV+lLrEadfXCrRCnCrqzZ/eEn6zYCRbS
QJ8NeWhFc+0eOdCP9hHbH5iK1wl+xNeOEkMCRcddhF4kH7U/52UqaYH2hp1oJM6v
bZCkrbgDQbpqBm7xV3aB3QS5hRVXwJpvgZDUlfryEIS/lJvv/k45wYaXknIkMMDZ
NraXsKGlSTAf/C3Z6akMazXzc7OKB3jlvvCv1gdNzcnUV05J6iFU3kQUjpiMkZ2/
tXbgJXbqau3QOskZvCGChQ881XxoTgBKsVZ1jLzjZ23/ROn7sTUrseDGBT7KO7mm
fv9WdMxisFguQ1i1JCn52npxPWaql1LFfjinLfQGhlW7Hh89V6zFnv4Cvj6q70Qe
aZubQTV4CxjsGxkapVM9TwEEnMB7wVurNyFnu4DMZ4BQkeSiDI0a0lmiwmZeUVh8
MItOuKyHNsz40d1htcc/hRgpbqjwJxi+V0V5TPLn9Gq4R/oNdnJBuqjQEz14Qdv2
YfHTu1GnuUqzXkVQmFlQOHFB8BjmS0uL4oKlVaxEpBLQwufoPNuOPmEMvrbhJvOF
yhgEvYrnrNG17It8tsITqQhJ1A0ofrCgDuFMRKF8/PTaeNPedLPw7pUGVinwhJER
kbgf3XIc9Dj7ul6toY2DKogJ784QXJGsGHpU2AISPcLN2V79Ka5duNoUxIYd/QWs
9sEyWOzQTr8IUu/Ufzl6Ew7PjUi68TGI6PRF8HcUR3l0qnNbqbfkRHjK54e5codS
xpMt8ge3iLZ0QQq9NB/UBsM5dBTeqKYwg2zi0M68Aix1yg15zL+u3Y9Em/olySjQ
teGisX4qnRi0qCqMFT0aA5oGRjOD3bNBtiSVS1BrsCAhsN3N792OelX+rdDgpW1C
Qy6Jxln/r5vPXR0SwNcAYO1JnePl83+lj3qOcceg21IFHDeu8tZttfmxjDwwFJz4
sDE35XQHjmKEaV+2Hy3YknxnqzsFSPYZ29/B8tbGjvlJJQF50hTkUBLRq0iNHNHe
03qFfZS81vljwm35h9ghen8GfGCoZS0J92Fekd3a/WYULzxeDTTo8nsjKXgUhPY5
ZcFZgPnrfi7CJgHwRQbWFNgWY0YQ6rU3UFe7X2zOjV4jmpWYiVgHoHq4RXj0ZRfj
J9Y0Lyor638BtthckmhE+afwrmK4Eltg3deMrh8MzLsJKUnrJ7n3VRwF9upTh4UK
c8umWC8N6dmk3FCgeWa9pxyUsvxPp1ZNzDAZ71jIZ9oOXuAuCOcrSIaXN4eOAmPE
Ee+bqQXvlIDxJLmHvh5LcywRODFZQ355BmfFKMUoY66pEonV4+FX+tcgnbxijAxx
zAzGVQxdh5oK5S0KFomvmTP+mkPp8OpxchvcD7N9cUQY+wd9pQXJHTUB3uh8c7X+
vKGa00nmYx0FplG4/a1NKeDeNC1PQmUO8pxAKzboEEyx2c1FWDievBFYruW1BSQT
gbp6PzSZmJ83XR8knnzmWD12S8G+5EoKM1vLQvs+B/rLQ6uJNyr/OfLoyvu6OfTM
bmvcnax0jzv0gDt3ZVvsaZyRotFPj6ziIrx/Swmmj3eWyvsgpLmz8dxp24LrLs9o
iC6c/q5ioR0EqFTQq7B5nfyTlTcreNnEd4rnNWnKVyv8zoiRSJLX/Qbd+LrAbuYq
FJfNGXOSBPGpTqzCRCUKfHJn+i13+GA+5iEyrCCEpQHm0ZGgEydwPWAURdYyyW2p
xr/AAnp0GoMPL/ZBos9zQLnY6Imsula2l3wBuMLsP4iWmNy/LzNa0YoKzEF6lEZN
N85A+aIGQePmPa6miKBtr2GDaXT+3oMyFKDc6wHYjzLBC4eivx6dgcefVjs1tbIj
cf/pXWk3CHLEjZR8le+VPCJ9nwA3N/GhFYsRyRPFM1Pi3eopxbLPfNRrLu29mfys
XxsNB/B9YSRhS85IaZoOAohWsADUU2ueCPNJlzpQVivqy+YtcHy8/SyhQmidpzxe
+ovglm1uacBt60NCAeKvIEyRLG/WZgUAUzJcdFHY29wiXKhLAAYCZTNB4MEv77Ze
BrsR8vc26qNmI3k+n0LEFrbrNtX3EyFloJHF0OzCY5Vx2RXinO+8vBkUOxVqofqf
o6yLsL+tb/1hrjVf4q5ANQ1cvJ8yiKNsyRWKMKz0I4FqV7gsrndwTzlbVLffAkEw
Tr9mU7EGteK8TjEHpPw1Av5eflAgrvRb8pfU7Etc2twWmAhwczMAwEGgsLlNEOxd
taiqd64kJeB1g7/A+8vTNtTtHKHNwYa/TEaLgSghLYhoFPpZMZa9Pnbq0jA3Iolp
fiPexvVWX+E15K5AzLKHQYiOl0jlTQ3Z3PvdqkVGHMf+drUDWKvj5SIobfHb9juI
p6sbVCiULGCUP6Gcfkitl0QkTJJh6pbh+Pw+L3fxxT202oeCTRXuOzk1LgB29Gom
bpS3S9ED24cOOcxISm/7uJL3+xT7fEIw26v2O5++FZiFSwq6hZ6R9Q095eWZ6xb8
uZNmIomU9fUGWIDTRPjr0PSICDJ4gxLD2eyWvrgJP5cpUllNu32mpX0vimW2h+0b
1pygJQxuz+1g/kanJVUu6if+hLFXXkVudvryXEK0GdrZqOoQ5kJEHolEsVbeY01i
BkkCWMM76aLCNBQXLGFF84NNECMqo49AcNa5rA/muxktNll82PE0vzsqNMTBwEJn
MGAcYHerD1T32j1vZS7ZFYw2ar8FkLqOw4VNj1ojQs1Rimxt7t4ubBjWVDO5ChZt
SNertQxhY6VSovNEfltSLqgJdMc8w9QA0TH82q1cVkh8s9jyBNO966DpL5+9BgQR
DkGFT9MCd+5usWW9r56HDw110hTpVCexwuR3mZL1nxXC36lverBHKKlO5g5po2Jv
qU2cmHAFVRd9ekWL8LuQNFyommlH88cqRpzkr7SVb/vTuOSSM9Z1ANhwq0/7sB4c
mZ5RvjDRBhk3yZdHEN1EEOor75dAYiUQLSWmo4eHvA/YyaQTg9vaaDkTcVvR6q+r
MdQV+SHWdzRqU4BVfcHr9bXLLME7yGKcXBMtFgEA8wzwLN9PcO4PCnmxzuor2rbL
lXO56BXHJPPXTKaJMlEzCiQuKYyHT4iaCWA+BE6AvOshpaAZ6vyELITH2AvYDD9Y
4cfcGo1RVa1IuBLeJOEMAzDygcBMusI1KzM8ehfT1/sChOpV/xfKgmrogeUGakdF
ufB7G94WdGhyX7I1UzhHNVEF2GdJZ/QQRl5de8PMaYOhx6H14RCPE/AXeU3wf2Go
cg6Ay6SWY9WAUmp3LZBMgWwaw1JJel5YlGEkJHucHigKNrxmPaYBt96ap4ib2bnE
+wpF1AKkPaWBOO0ygFlq6AJWGUXNbcKtcrhp5aNJMm9oBGOAwvhuCB1VQa1kikQy
7nC2M3jWyEk92OrXoKd2ksfaRAs6ZGkoHSX3T/TjVNwXEMZLZ24DrAiu6Jmqw3B+
KUNk90zCXg/DQw7MGPx8etthlVV/t7O4jOvUaGbDz2cS1tsRic0e8dZpjLJ+jYvA
QzyGNHWOUOm53M6x4aymlp7yhZ3T/mBNcMtc563NerD/q8iWoR4VDFBRJS6+P7yF
v7pEBZVgmuRXB0WPcqZN9Paga2Xq96KYWfNX61t+5Oc7riZ8t2VrJRdB5TvlwRgx
OdS0aVyMqJ5uOtvLuN66iBldrfuWkLwdc9YEny5gj5lXFs4A2clRN2/+iy48z2if
Y1I6WOH+q6eTw3R7wYaikajSUpLtNk+UyJBAJrP1oiuDRsQbP+Q7g6sEMcBcNBCo
Wy0Ui0wpfuRWcpowawAI0EclWZ/PEmhnwsH/gZ+LoDKSgzXWFwToobHXZlJ6cWyO
CdEsas5qCY41YbmvSRkS4rclwRRKXtpae78dNu6bW7289Z1giP3PBo1EYq0D6IEd
+8w2Hbus0XjBvm+rx3CEcjk39DAuD+fhfgpvHEbtaJEbIRk4667ZckoH3Z9Tl7fu
EVljP5CRGvGaj3kCWEfFN2rTPKs9P5LO7YlwvGg1tKqVcumhz0VKP+z6AZ1Spbqy
bPNyxrSbo1PfIrWCo7ylE1c9GNEdYCgCmXKV1I7qNr9j30gMyv/TA48irTi/FYOX
pNcy50qfnil5LXUxjN/lVhqvwG8LvYA97/Z7ClK6Hdc0R+pzp47+A5nNBgvMCq7D
Z42EakM3RhA9lVgtGoMKzWgdlY2GLsZWco4NhfNjMJff3K1qybDtEw4GeTMwp30r
oWgENlZlcj9GJdDh1QO1EJctzLY+Oj8Md7jjT4JjToFdsq7vO+jxGxxfwlsjAtWz
/0JYhLkUSrbr1o7zzuB3ohectVmtfbExIKyKAvvyKgDcp6+0n2rfvHVa01kIvRzs
/rtPX4qQW+WuuAf2579G3VzWtl6iZC+i6QTHUFajplxkcom8W3metH5rHxxDgiUH
tkGiunX8GOMHXTAooN7HvBXSsPdYUuBKDpbvzdwq5VwjRX6u8JiOgCC7goLufRU6
1c7sYJlV6gAir29Xsd0t1C+BSQ/ZzvblP72w4TdU0Ud7byKMP0YrFJ0MuIUVooJa
tnd7GpaU8fpXsm3Imm+XzrYFGkmskpTthlwfp6mT3bPaTbeVMEmQuHZ7eiTXeOZ+
uOzMO1AZj4Mu1nktYhQmB8YRL/SP33XjU85dBiqCbfAy0efAUbtrmXRrGR6v+X03
8sLFqBM0H97VpH18md19q5T+E0nOzNbWJQ4KFCJJlYuZjvxxGLnAcuHbmKtFA776
RZ15Xgkv40D01izo6dRcOPwWOmtBD10CCPt24fkAd/WV0CYEDjokXhVkYlEqrxaA
RPXLXsXw9TYxRG1lEy4L6LrcY5fZmfSSoDUUljIThh7c7yF3/W+TLRlZA+/ju88l
Z149qVmxJV/aQ9ugfTn9m5rMwSi80ddN0n3QrqOcIpYzp7nEahbeO1qt/Xkm1YMJ
FsS2CWEh4dlwroO5GgWStnBzJpWzW6OtaeBJ3hZN7s6AJ40yVVmi0pTPvcZVSPPO
TfLD8wTXPUZpT6txBnlGADFfJSXja4ghPVBBw/QKl1KSN6ZYnYmOthTNdHIGZISG
KMzU1IFn5Zp0uOzoEGPvj2N9Ebl8swq/b9UwJ5CiUaqtvy5mbId0VcpGiIxzOsE1
DTnMC+NAa3oG7pgOWA22K1xeU6e6W9tbyJ67IEywa4cqKlWExNKO2uS7hUWZhMi2
w4qVLlcLuhSJahndrB1r5dM9qQ23drfnw37nxixD3jwB9NwQSE97yaWjQgqRfdPa
QrTjld3tHC+IXi8Zx9jCN8DSA8NLMuwV0UMAIX0UPPRDta9cqrUau9E9GV9YWHj9
+cKWj1BYmdAbY0Qzziat7KuJg8rgzLszSZNPB0KBVR92R9BNlZgheV8SRWJuuwqO
2xyfSHn56N1M6q7DIMzDn8Wh84rjfuayKJgI0OtgbEYtj17+uflRjmi6Nn7vPv1i
0NS0YZmX2z+2BZJ98O0hIr5RokHD3JrmgxfqbkAb50f4+PgGukeu8xV5jrtA9Gsz
PrG8NkI7/iEuJrFnCL7vQRyvoCGTOAatB1B4nm98wCJmKwy0aTS3/h/lbcxW8w9d
13hT2n3J8fk3R0tpVT6TC4FrSUfv0Ajy52EM7cduB0H7lhqaxf8CGwL2Zj7N5TRY
k2pKFoG4d+MWoHAqYmvEZPiXYPmQ+XsV6w3HDtMvFpvE38Xn8Yrb6/Xtu2oCjpKa
HBTcfdWOLOah5I/AfEt38zn68aqSLYod8hwuwaSR58bIWCwG7wYD56rIxnSfNrZx
ubs3GTUyYqFgodiXbcFtIOc2BxgpcLTe0eHDpmVhlTYXK3CQ2vxX3E0/QYjFiJ9F
RdBsJZ52dU6k2zo3A6pwBvXUe+mTRGjbfizpANMK7U6bHWhTrbnWuKMyXjC0ObXM
Dzoko4TD4g9cLxCnr5eEp2iwQGl0UpdOimjeXhGU0Uso3NrSpHE66a+5kAwAsOHN
dMc0sfMSBjMaHSFAVszwWfX3/lgqFx1ptbCc/cupDVTTOADR6+0NZkwiIGPP10FE
WvVatC6H79SO140jKakwVbpEsKkKVoPzAIp9tTGzs8Cnk+qTzPpDeF+E4jBgtsTN
uQ4YJFrganuBEI0mvp4qeK6AWC0yj64FviemDfwiFuruhZuB0xbUlWOVJbS48m44
FLmUrdgrFSsKlbrAyo8t8H6eW8/JRBQoCy3f7uJqFeIcrwd9+AQTyYtXnyl+PNgo
h+dktBK3ARwjV/X64oQgKn8NGLOWyk+ARcaL78QeXCyQOMpnXBkPcMZCNYE83xtn
MNbIUyJUy8JimOyJ43X6KIsigmY4j1v8kID8H4tuIXq0x84qLhLIjrnr1tXfyP+q
yk8uHNSkuJ412UbXlAEYwusbwf93SupnhE+T6qRcPSjPuYPOVSmOTPfJjCh8G6PZ
TbmV+myVb+e7sRUuUaMgDCpE01y9xZBH3K1ZdMDBKzsAZDSJqYYSGghwPaDhYc2a
vJBCpGxvPSSElRiC54fgIrW/nJaOYeD3RrWsnfbyMWEha9MHppKOzAMvZGY2wuwP
kSK8rdYiFnPgw1q45aTxDmKkKjz9Tzl2uQbquz6fnvlaVV6axtuFPcHq+/cmAiO2
zl1A9nZEKw0UsD2J7hhkgGlzUXZbgkfY8dD31zH+YxkK3duHWr23B1Vu70UnNGi9
dHwIfDHWBHREyRGLPVsqFpvn04K2EqtCjvD0FlnTYDmuurR+Ki4JgPoe+5H5NQXS
/4NcHhAOG2OGoOGPy6s8ru4Ztj0PtU5MTsqnjkJMJ64W/qsH/1qGRFYfybtH2t3U
9aFmV5VQ1BlOV7T4IwhJypit0XYswBu6w16YiYYJtoC8QNitSv/l1fmIBPhF7Yfq
XqUntjQW+/3gunWPSeGofSNfqkfcV3ghCV1eGniNwvCba3saKOBbWKKorNdqK1oG
sT/x/Dk6XsGzegwSe5HvgFp2cilVb7kW8rG7dW2dy+M0zb7bkR/h3DI0Wls0eNL8
MjoaLYYhUqgEg9LmZ/FlP2zWSAIOzOPCeZ/DLgrBMTZVnHjcp6jnPzCWIdUhKDY+
eYiwYNItCPmcn/opjSgoRCsqhsGjkBIELHmkew8JUWQYTfhGROj5GToNJ6z6JfBo
poyUUo3bMr0t+82i2nb8vPJfFWWOgnNqBIdlR/70ob1pkB1qByGwaf/qsUR2lZvy
xLgPlmul51V4VgPrX2fEzzmIUkR4GeyK+BzsannJQhR38l4H6I4gjRqjT7tGJXyx
0Y5gNln/Y0VPZAqB5y4YOm0hpUnFcMYJ0Eb0YYjZWhHC4FOcerLZZh3afucRvWaS
om/5b609HrVOC+NA1jdFz1NXJSBRDdkz2r1+6WKkT6bR2b9OlmF68eCJ9n34Hake
m5jxOt6pC/TBGrXsz46ZDnM3+w1JcwPju2YSCfJgl63yYAsKCg+LIuamM7FE96tS
5evQRpFPgTGaXLx/wOhg4fwbr0JRa5APSYgHXCmQayZFvWSfuFUYvj7+1s2Wfzoa
57jYmdqPoM0LHxWxNmNHPTsgxZKsbZv2gjxvIV/SAcUSx3kTY7ofb3bBXiIibsxL
FV3xWqMYKfkwSgRAfLXHvVtT13mj6c+946CxLhR+BjYBFH/Q8FXmJ1sjg7z3Wxa4
l38rmbNn9zVFihaYUuztiBRdcsx4fW0SI7HkvvTiD0nY/M/mnKygIwmaFEeRPRbv
bTLoPdSOgNfI3l22FkWCRSgsywFUjLIN5Zfg5Oci7Zd7fUP7dz2C62l4ZvMkanCV
agnEJPFiE+gzojmGVO54RDTJKy9XhkL1uNr8fcFpZYGgX4ocaLC/lYDDKkWVEnS9
S3rDU2DQrKakxJTnR5yRvAM0oYjgD8FxvVJiB/hsaTJYB5N/nn7biUlnmReSkkWZ
i/GywriZ0pCAUBoEm5BQkFpiwmaweJoIpJ3QErYwH8Hh0UEdMhg0oa3v0vSvP4F5
fOt/kzWjorzVujcD5zqDD7THP/9aCp1oSTTCBQGNfGeAj6UIh0EiwJLsvYK0yoXW
+uPM1/WjQC8TltIHPtX/TA2WN6fZ32RK5sMEfSM5GYPsPy034vg7eIL2QFrd9a8g
RIUn6h03gjwOiNPQzZzEEFKXZeWkckEOr1iUdlC4wkzWJNsuIVn7NWyQ/WB7maBE
4SDijMATbqJYCON0kZmfJO/SdV6n0BfkvEIfQSI85aKhTlTk/Y4wudVU+6PWIE+J
3KjtKybdjA4bsHDeqvuVwMgbwXyjwiE5+Trn6c3CiI/3ikiX3HsickPjyHn4QxlO
eP2+K3kBoFfiB+72KJGXRM/IFGuZOYjwvAsxkEUq4aI603zZtrZIP7tuzQfvD84c
Hwfd5j98jG6dhrXidtCyyjwHOJ6gHQYRaKxTtGt26lQrsLmtBQajFwJ0dAf23qXl
q+YZ1sm0E0yo3Cadzxv8j5ytZeviK8O18CH069Jx8aY6awxLE28A10q4/qRAJth4
2zspmTSSIECwX2mfE17A7f8X1Kac783cOc3GbHNJpD/GgJMAsBl/la1udRvNSW0D
/188QnZPJpETS9jiMleK6beWBK8mmINQtZ4XVMtNTfqIfJCZnS0yEVRq9bMUTIVO
lo6DQESJWYSUy5tQYOAAqE3p02IQc2hVh20HqwWjZ/mr8ITGyw0UN51ze6cPrF8w
P3r5f9J4pnhj08Hj7gE3XXUHtWVzb+Dxvd/V8iXsh3Mo8w4se8urW58adrMS625h
sTam3aqq7XHDsQRfrrPJC0wyeRzCVRwuj2s9+Lf0q23L9VO+PgWPu7pgj6x+4GAJ
9on+OtUup7C+YJQY1XiyOjlFlekk36QOH5AHMbYIP+bZLbppRZFw03rOzXEJkTz6
Ke+uSCCMQOLIkOZygoAhAZZqP7JFh3uBJK/Q8yBypkij05rrt5/mwqQRDSdAi8eA
swsCbC2R2TTjLdg+lTroILt55UEZ9KYubTOJoQ2IQCmfJq0NpgJCc9X8jYDp+t8T
z7zc/rVAsIsYdKasvHX7M/+PnEfs06UTCbN3zpWcLPR6ICBzF87Qfb/KFzuUFp25
JyY5tQLyB9IsBCuIuY+Wgu25w4ENwJamQKS/qpGno9cxMIQ10hJA+6oF6zt9fuRj
3vR3BvxoMApzcQwNLWQ6zcIWcopti8x+rlMWqZutlYs21UlSyQs4smCpBwgsqUxk
25i893bLS+wxSF7DU+HAV9DZ1GrnLslxiJGly2CWjI8jmgboJhBI5G6VWthOvzI6
qPQ6y+SuAby+OBQIHwLhWXgXW8ac2qweYSzngTotAg9Au+blYv4OHj40+vFQbuEr
mWdx9MGKB8PnZea+yImjd+/lREgrS3gIcXhDZKwLzt0q5BZuoOTTfEyMBLiILuzE
xfxL0McBiYEcrX2REqPHtf6FrHGBjrqT8UG9QCSnRy5iwrNqdqwBOclVoE3Tnxcv
RfnGqmfEA0Hn07Hw3HyWWavka1D7JkgnR/B9Eji4APCoi8G+/DxDg5F0ly1KsWsZ
qzDR/5zWlcuRcyib1IJ9cbmr/EPmrR+3yOxQZmz4ujvSxfiQv+82o2axpOXhEnz1
ZxuOZFcdblj42GhZk7RafmVVMZCr3fH2itHhXh1OdsaJDQwvjfcwDWV/0yePPFFR
OKoeNGtfv7QDwYFVqlU4x20nntgLevL0WigJ4ojOo7O0tI90hyShAnfIfmhvQPS1
ze5lhPxtYtC5CvP4NWxPXWfwvi4ktaNXLN7LvUIzyTQoDKt7Hb/yuS2Js3md7Nel
rgOpZ/qG0urn+znI24jACKEaChz5oWs4kO0jajtij47KzgTXHoFV5yGickFIo0t4
g5dlkRqUIKrW//4De2crHMQkw1V1LkwSXw+kMIcazgWIGNyzRt0IqHKSVEW6q0O9
+ecgfdJsJGvFMJIGFbJkV5rx+wr8fKY5WyPCs57NRV9ol9CtG1G/BxXXfQM3vFo2
nCnkb+FdI0wVTINUPpZTNvV0p9VudgzqDdNvJ7+q3K4U8I2VhO/aoDdD3SST5bSI
0NiR0QcLaaIdqhOnW8yGMd50XgtrrWT8my+a3JMaku9K99DW9zwJtCKn/Esf5bi9
xhVNWz3jLiYYxbNYAEHgFlcT3zcPDbKgnS7IabIc4x9SnQDeNBx3tS3rMFBiAzUy
XqupJNqOv31ojpjss+Jpxp61uVZTtaeEyuwyiwFYIeEbePBuXCqP5+5gzSi5PKdP
x+YnF+70x+9thQj9EFI3CyAsbebVd5aGxWLrCncDetQKMWthbc79WcQ2R5NPx3b+
00JLpjs6cgnSl4nrEk8I0t1lwum7ZnQmZUKPoZQeIYYXnoAm9h1yNg5+3m2Fqre6
N9UTI4bTv5hh7CTxpq21CuAxZENuOt01Ik1yOrtqnnWeNac+oC5C0I5GUyKruDJR
4Hft7cVagdfLSrTYAex48lvswwR8xiauWR4Fndz399M4NKCz1wf+Lqo9n+tDvdyk
Xjk8xh64U81mZNHcB45YFpQrZAh8EmEnJ9l8tRxb7nhXeGGvv3OLkioZUExKy1LW
QA3jNVgRTQUCIMeDzFgAWN9jQPcv06j8fIDDgmdK5uoGZghih3mIXJZZf3nzuNiQ
hp8gJk+BsTzCOKJzOT5F4pVBVEUkK0YNeT6YNNrJ8AKuQAB38BeL59Bc8C3wS1i5
KIUCiMPxORHJeMjjwHAOS2jRN4auHv5MYLP5dDWQ+6Yuhs9LK/LZpvaMDhJ1ZKD5
bu4uwvw+45UXtmddsy9XbPkI7QR5aqAR1WwBY1gW63gyfEhloUxh/t+Frfxh5yYB
3MCtEzjGCP1LGGTiqT/qyum60S9Ryypa9fVZvgHqYTzQVsCCkVuGiToE3vGJ7EhJ
LZ0CQ0O0+5pOxlV7z9PMxCcUMZm0dHY8gb5sMnaaUOZ7ED5BBpbYPgFG0TcP37jm
ApjEOSmq1gxmwazymXUpbUMQlUnTI8CMnkNhktXBPzw5swm45DR/nekhrhPHdPX2
7Hn62Nb9q2fQ+3CGbV1QfAFU1SJztAZDxpSlcRhyMlK0lnzGs/EUynxs8BAm6sJB
0L4XodBM8tu161vVgH34ugP47yE/HMgNQvPdnAI9u12steO8Fl5GOPhTwOk73URS
pG0CxoBA/BarFCzLdM40vqK9Yr6ZThdMVn5jeN1kWN6XPs2AWGOXmI3D3ZVdlKjN
J16Q+1DY9dFQPY9/JYWEfPWwjrCiREyQA8p4jSsg8CcTXpBeAiAhf+lE6SvFPv5p
dh4267y/asgDg8m4x2wfX3w21EHtzveC5FEnk7nso+HSh872pJD0W5DLg758JxKS
DISuImtKuXRphZDGNbJfeTfWJKaAvHTPL9rU7pfJxTOiuNsvVsMmSDxFFzr3BOPY
t+A27UBGmdgPepA1Rmc1TIt4blnUsrjq4fRabJBFigEQNMfx+ty9cM4GEJ04ylNE
8vWxZX6HjMciwsx0A5GrXVI4U+e8srrGya/gVJotX2k9ZxMaZUOpjgUya+OdUFPt
3g/7JAPfsEfjzq8Fxr1xOJXCopCPScxgqUhZpWn6jsgauN5os57AG6KUf/qKg3sB
/fhRz7rHRQU78eZ8bc+ChWqjN1ruoZihgdAkVwztZ7Vb6hvM7T/mx+2ynz9D2j04
Xx88e0YzTAdGD82utOeVRJv05w2GddQCeekIcJljytyayCbpgz1dqsRwYsnezboa
qFj5QTjnejWvS0wfq9qwKzg3LEu+fxj6SVo0YPm+zsAaRWhfD4sUfoKngaSe9Y9q
g8loKnbR7aHVNm9efTfY3dHnW/msgqY/V27Ok80E7SO84WeY/4vKaEGNT2ZscHz5
5NAGBPmMAu79F7B6hpbf6/dhFTt6FiIBDnx+IATjBwdetahD2zAZteHB4E/Q9XSx
8Hwwqb7PmLY8ZWYkIYjCinDF7WkMnxk5XhJk91LfdxunBYpAp5q2nekMQyjRET/V
bIcaoq8K3i2b2mVU32cyX3l7o4e6SPWC9Kq6xRdhj9pbLOtDVSrwSySaer8QE6f4
/Jb2y0XGOHSonp91AoymS+pWoqc7lg1qCLy+vCjPq1jkNqJRbB1tkwobRduxHWXy
PGVyw9Csa4BgXTiDLkUnk45fDJVeQvcJxwKtVc2hPSiQ69zvvxP9CxM7y02z9tuP
yYYXdyrRQZVMDZJJEr1zptZX4o/jBpHWwhrgiuTBVQoNOJLsG0l6BCaHjI3D32gX
J0r4rpBBfP0scM+QG3YCRQ/y87JWegg3pm/oMXUK4rqEYYZJ4pLmz3wZXYX2yeCu
Vrnp7uyslpp5k6vD87aS0+bc6Hw7+bkWnmS7rj54VXt5wtrSFrMNAl5vYhtf0E8N
H6kDWPKw4BZGmzE2gK47NIdR89N5NIsQhbAdFc8aCR8gz7E5Ndg1cPl9p42T9xrC
iwTo2++INLWTAYxu0zCyfQtNe660ir2Flwa+4cdHAQ/DorDV2zQoUGaqeefO54vh
YoFFPXi3h1mzUik8pXnOEUovqk4kztA1aZ2EUlcvbXHnCnBuayREux+0XpwhWRVT
JhXGOYWGBACtrU9XXAo+C5UbWINRMM53at3tcJ8wNDp7BCp+WMszkYSdxlCqrqSp
0mmE4cDDyGykE/EvYqEGUYPJSqImQJsdAiGql227w6Zh4ljT4TaLVvKXgJ8KvgOt
357m9akwyMFeZ2F9VOrBNyBvIk/Q20w69AfKgQexzYNPifkq2/Jml6LI4+b1BvV1
A6rdfkPwiShWA0pJ3XPjVkdrb6tXorAgZxaubSljBwMpq88PHjTO9hX72TrBAnl/
QfD1qpLYvvN4chXNHD/PPd8nsA2NTxOPkj/qD46X3X27p57B9FyeXAJ+Uf7vvsaz
c/46LLRHGcA7HhhYhg9rixi7gfPd5rJh/WI/XdoMbc2CbJ31h4WTlwMMymCFPZrQ
UVYCWykyTw8/l6QStjm5DLE+Giw/Jj1EoiWEzv+Lo7oYxeD6IaenEEOhR88R/H4C
iOpjHZhUKV6Fq/k3JUw90kwSPhGK1lEi2q2QhbfZxFrCInWYxq04cTES8VlA5lA3
gMeexhARhlqh/RZqESkTHXFmN/fbFe2KwHYA1NFZ+WqYwFXjr+Iba6Z7TLyiPkyX
yeydwhUuFD2TV0gPt+uaIfYM6JzZ7BYDox30dldGrFYoRQ5me3KX+N8JSc0wMbwl
R3Vv1yj3ZUcAmQFIeyyo89SjoUPAiFlGrRRn8Gyc5zcz65dDAx0D9HheJB1oeIS0
ZV4/TPBn7dRIViqZYpKlRJqalKvbYX5kH7MaITgdsn3udtntY553ALiOjGQc4ton
S4btrciA1X0NpSfinJBI3H9NmkfC4whUjExYPsHKeh5lstxrCkoN5D0gE6/psIBs
S513Tirjg6l4iiRrqOrHG2Ri1LAiw3g4vqoZO+z/ktOBHsTLd6ZlGuf8TlYocrO6
5+LYvFC0QP4yhep0xRo8aETfFNuCWoKGRuJe1t0ghjhjSgee2QewjbVOIA1B9jRc
sh9/g6Z8xo8Q7flrCbnY8IC8RFM3U6XeIQNsvVS4++J8a+W0ZXt7puA2ImCEMpIe
ZgufUZD4vY9TKc/EqJuq+FI6nL77y5Dl/e+Uy/4hF5VN0EST9/dczcvSg7eMZWVk
efLfeqxZAMtbuXGdYBh93injAEXXXJsbs975X/8GaHHh0JSPWzd83JQ9UXzSj03M
BO46FzjityfvFKiGT9G9ut9MXGe1+fZL61u8SKkhk1sT4GYTGOKIZf4nRw6E4p9S
0ZFe5edBbKJeX5XMXvTpzXXNPk/P4H5mEPIcmvCPlnnOLzJUZGs5PcR6ccdAsWnR
SnM4Ar9TU5Q+BfK2M2a3QZX/cLhS0yRXdRK+AStKVAINcZhfD1MqsNxGdAOgYzlw
w1SUFXoSQn8n/WlQ5mQnbhS2ywTpWfcUnrzgXQ7pF1GM024QzH78QE9myEPC/GWK
1euACPleglxnJm6YXdqe+Bn/TJqeaclqdmDsy7eZ1j8i8ERk++1hJ9RifmSXHpqg
gXHjLLw6ic5+UvbATKBIBUKLoAOOOYKvVAU+9U/ocxS1oDVlA8cWjKCODqNUKJgG
v+HgRyI0SkSpL56yjLoGRrwbWSzg+8Kn43OZ9JEYmKfo33prh9nr5NGL3OtZIO5S
Uu+ecVd95RRWIP2eKNNYW9hF8grkuAvj8uQMpNV/CC8i7tzYOe2IpLcoenOxbpAe
H4zQFTXoVQ9h4e+tQhUGaoremBacDwmAAe7Vh8epae7IkxeDDL9Us8czejJbFfvo
0inLvzxpugV3m3jpQ5GEGjNhRYJibATJintuIvLWEgKYPLUJNdf+OTJb6LwfYZxS
jf0EczH23TxV6PrTotao2wUOFitgRiH2ih5+8L3EALglcOiLCS56FyIwoauoWluk
SFF5T2q7AmMAWptN5u8sEuvU45yFkYbFjqp8rU51KCEVIDA4Yw3O/cE5E4sI/P+/
LwwY8n/IkDweQyi+GTHbJCCWOWi5ac+xD0S2DdwzIv3UYhaeQDp32JbGs5xE4LsX
IZwhTKUYkKMDoo7VfEmC4A8oMnw7kd1RitbPVBYw0Al1uTaPzY3N14T03DW0FVad
iYiZv5MA8yf68FovG9Kr8yGusDNFNHnQC3LjAOKwlsxFmPzSNUccWZtbsjPJPnLn
pwgDzuFeq2HMp931mzwBYPaTDt+jDsKQTUK+WV2HVFTvuFlnmbZmIeVRykqNtZ3y
tHt7KzNWgToqWqBgwkVq/DTZxNyU/S7JdKupjGHAO76NRGVr9XEkCWK9t5oLNtCg
SzRowkCjrgO9WJ1GNNcASqHaqr4AbIZpfrYYCp4OPzJNhG3NhaXWO2+XuWeJDYB7
cHbub7yRBaO1QAOYnP7BgCHPO3MzkXViKVjIyYS+KjEBH+kFuNpdhPfGwfOG+E9m
Zg/EDgD6OcWMAwh3NTOcwutHqEUg3U03wIO3nz/wnlECVeMboIFmiSnMseFSOoX1
zpSf3+gz1+fpn5cASsh1Ek7b+TWkF1IC2Sy4dNL9sS+Lnrvdum8it/NI379o2IUU
XRzrNrvNUL9vPT53Q+VmoeyoPf3hlDzUHKdVfklhXV2mYtQ8N6LU7ZttOvqt6iss
f8oeY/Ab+bOsO4B3eW2quyw9bZvf7S1s5qFx6RsOKwXUOPkHkhkKm9TQJIcwWOW7
ZLIXH4p5PIjG3qghlCQIvmSQh/IaJU3q45K9TLpEHlOhVX8UzPmMGoYanfFVEKSp
GclCUpbVFZ6qDC+oYBk3ppdT/Be2EpZXpbLinyhy+6Dr2INjaJrhlo7uCL7ucCcL
2Rty0uTkxUQ/Hcr2EqHA54JNfS4717ZhVGyD91cLxE7+6KrtTeSsa7oEgaYlYmgu
071ip3WKgRoZ5P+VmUrytLbXCU3N9YrXNZl6u+0KdpD5reLEd4/j95ktW4ZmySbS
lGiWu2ZIkk2S0bl054CzRyCmojSN+fyHm2MnQk43Nvi0FjU8Pc+RhNsRJBG5VQZk
UZxh8WeRW00jAB6KBJvxXdkj5DPNV5IIVQHDijx+FlQdmWW28SrHoFB1PzJgqbeu
C/92oovN3M30xzlsFUZJmzK3NGM6hL5QQ6eq9kgqIlafQif0aDftWHSz/dF/+fL6
BwhrrS9lrWevi1gt9smqdkiktoj8rxWntPle77v3qn1Js7AoOF8shpIeoKzikEHq
srPJAxJBx9BJP5E0MmjoPiB+8UslJoc/mU65UdlSXabyaBAKykBNwF5H8rhtv//s
lq/qCYnKrAiEGZ8+uLHZZLwxKlqZLxULVhwTMK1nH/wC5pecX7FxdXa/jdSY+3IA
sPF6Z+mMrZsNg1fO9ZVWrG9juNwq6wiyXjEXQpML1WCK1OhWxOV7DPOP4EKdHMIg
+JYKGbVWWZH66SSVq7V5wYMKKdesh1r/medEXxnYXSmQ54REPh1p9VU7ZS4OMgpz
Z232OW6FMd90eBqHGjJFm65kdCsbh3HGeiYzqB0oOv6fyPxv/3Rb/tRCwZhjbba+
L6OXALvhdraeMB5Kii7guJGCS5jddDEUu1opx6k2OozY+yhgzKBh6IXIxdN6oEPx
5iZKUw+FF5N08EsqzmFDKyY5FHDApWlIJV29YHpHGg+adwaj8Mv5FZv49EreEruW
e85Qt5OCtM6VpjhaYwO+UqIo9vx/50MitwDqSuGCD6GiX4wwxQmVJod2eLFm/XVz
JYqRD5+PuT7jQTsFqSBR7JUG1itb0FYMEBmDUhye5zN596SR3MhX0vyNQti1G07+
8CSXtwjD55CBWVC+RYzoN/MhYEEcjpl+vwMGmFQDa6XZB+mfB3FO3KlvyVs3MuI0
CgghHbWYnjiX7HlA6S/qZzZh3ETwapfd3koCwPl7cnlELalG0vbVJgv+QUFyENeA
2/eQvRDuaaOw+V9A1P4AFFklXwFFRy7/muSEx5tQqHHW+O2v2T9zldWNTLA7gr8i
tYggy9auqRFt84s0htOrIIu3bkJg2E2/OhmRKRSsbCcOFJE34nqfPj5z/STlDuo9
CisEhcJzkQozruYs/5d44F5foTCXTgHI0c4XcPEojRbhqIQejCc3D7lRHuMeZ/Vf
ME8cr7J/2U17NB9EGSzkSoxFdwFxcDNWM2kM4UtoT/cwJfmXwVj3lUv0OAZJB/0H
iOfpM8zQoAbM3zHBMX/vRsQlqYYrjehyiKGfABbfFdGMwyRw+8FS2Yranm9VBUxp
P1u00aJhefH9s+qqCHmB1yBcMxyBP7cKYa3c+/bUdgOLDDEOi4fCrMHah3zlzUU1
Z4AIHrWbvpP4+D+NNgzWPRvJQ7mp0ZLIEItJwfchtnKMd7vrLcOfZrkIGGOp67H0
v8bpl18vxnetRmbs04rMhB2bhdvdMxvgp7dX2QGCwqZDdgicOyaOlN7fQmeFtvDH
VlwOarqWs50xagOoM+vC0h7aZ9A68xTysClzm4WCmOJAPdL0U7JuBj8CRalS8isH
cWOeMOdfGlOL+er6JaD6BCRPnGgrz5Q2ZHzmxDNa79R9G1ChH6Rzw1HA50Xf/srN
lBUx2BwaapYvTetvG7G0Cxx8r+3BSm4Dz+KsRQAfF6oJv7m7FR1p0xJb4vsbYjVf
Es8DtS/ujb9HOTekeyYH2Bc+7Fu9ujL6lLEf6fn0vKTJhtt8ONMU+8dQnvS6Gbde
vlIIfQNp+zr/8UcUt5yaInPYlZoSNdIxUVhivhEhq9vOITReVbDUZmHoTz3a1b5H
HMW4O95FeF/1x5QL1MnZzb3vgyEgFym3jO6pLBLFXUkWLPsZGKqKbGWDLSXlA1Lx
xbwqq1vouZdxDERhAbHfcoCzmk3qTogIJ+SxzyUATBOCpcjI2S7p3tknOnv4a9lW
ZRzR/wHMndFEJbAH0q1TiDOVxpX8VLx8r4+5Ksd4OiNGhp1wpmOA0FYVSL7JywI3
ZIW/mRVPVWZ8IJIdp9rce96GMtdNGrTGTVrXdNxGtqq07R4xWijLO26q0D1KtL7O
6Sl0OWfMnit4P0h6a8ETtJJZg67YC+4bL+NmAIOah9DjSuNc09wNMFJEsEZuh2xo
EV6+Fp5CtTx7sJkECw/v+jprRsw+tWEYVwCxz3jf3ct7p4AlhirZQDQtCCv5CCVv
EG46orL6gc+Yvu3z70GXKUt5bWCGQiGasRt5RVoUbb1iW/5If1hm+Sj2MT8MdnZ8
SoZaqeepG+rQ+79GzyzlQMH24aLTpEqn2ASOoAg+4562xj5FpUEMedjKSCYecf6j
elcRZXWI/1gh7qX00srZVBYhrHAsdYx31edRIEbyhqoA6ru6mUP3hT3PCZiNNYDu
3kWvr0SKfufHnw00ycFlq7/l2xlt22dNUNAcEGeri6OmtzT5v/hpsZrYSdaYrdxB
BT7EBS6tzvag29nLQWoy/j9yfOEVxNiPOSUDPHEzH7ph9yC1zfu5kAdwH9e4Flxd
fkI+myEZ+DeJA5EmGQ9wb+2g3OfMPo+mYt29t5PwNHHUmO4aX8//9/igCRiXDCPU
2lqoSnGLUhCU+wiSHJW/DYXEYK6BPZNgWfbe12Q9/yIfD9NED0PIMIVO6SAR22rV
W6KEvUG/3zYCTLYeZAmr933+5ELGQBcxKVLyFHyYLlO6lSYB7MY1FY8zWf4fy0aO
f9sA3mYz/amfFr+uwbYkmRTqZSQ0HRYzMbgIg2gkcn5Fi8OcbxlYWxMHwQMDXpHq
MUgjznWkZOOtO7Ot0HfAnItjm5+BLlWyMaS6iCrbpxhptgBLGHrorcfmtnhIMHLr
DpzWKDjFgzhuHQKWkzRGXzwmYDF7FI0oDWgoutceTP28eOqJmbxv2PSwDVWMkoAv
Uq9HRyvr26jRGhkM+IVgdmFgDt/rrtzVJmvcoOm5WI+uF+AE8vqjAdX09V/HioWu
N3UsR6W1y/FeNtz5A1zCUF1nsrsn1GCeTRSX/k2ocn+vn2VbeoxP+CKUDKyPtjcd
v73nlIT/YNQIfo4SLDxBDquUh7PinuhvoOH0JXK33rjuKDzxsZcuM5x68bKfYS2w
DVRGlg+Cb+e7Rz2z+ca7wqxd5UENtL7A+B17bul7BWa5C69CWshttg9q3BLd+wjt
/eTTVUNawMrRDsrHPk6GpCq/CCPoTYoHL8LSp2QheqHE5kBvnHYh/Vp75/+K54jY
jRgcSbdmRc9tEl8Wx064+FESlrS+YE8JnfdVbLsx2jHFrlDHMHMxlFVbo52Ke2dP
aR+IN8RR81u3zffGx45jyhWfXTR0EJnr8KNS3DVqwW8VHY8G2TWrMymwsxCNomm9
XHAW4zjsjhoZymmNpb1qH8NHTiwX+cdcXp6wTSuqZkjmjo6m6T08GG4i/l58fiEJ
ekLWQr+8Fou9kJ8MSRe5dzk8ngSjNmJAHgrixhaM17pEkLmzGWgIPvUyePOYzMpG
3Fn5OkM15H2ZV1ZRSqI3ATU0CPZwIB5sKolnLzn8F+BoPmbNvDYpvEmzzmyBhdbF
ZutOmEJd4r/XZk2owoQ58TxnaaW41h4fLPo/rSZgDkJA2AiQWNYegj+XaddD9JOE
5LifACqYv5y2cArxTojjQDcfXJ+lq0RX9LRyAw8tQdGbysAjZ8uSVh6zvBtgcuAD
yeUDObGTljC1CP+3XUrjRiCJgzHZwEV20cL+m2W7Z7bnCXYOk8HHezbITDtARuGY
7ILkdHkkwbjKaJrIgUtOm6/nMgYc9HNyhnX6deZvXZ4rNN0z3ZxjvpuQXYbjkUkU
trt6DtiS2NE4Rd7zV6dE9a89MBl3s7rHhhJSIA6tdWR7B4LVyLjFGTKNhWHjeUEI
giIu+mp4yE/94zHk+zUFixbzXaVvrzItdxhwPY64JAXQnHx+skIZXDmh/sTVErJ3
jI8ae9Sog0wIodAZK9PHL+sjDs1Yet46SKtnsb9tsWF8AixwSKxzVt7vNapSw1HJ
FxdEXVn+aEvIuJZpW1gNBZBLdgFEqcAV8xfl1JR8rYtSCvBicm4cur5J99X1wlHh
93yvFNIccZ8Xtwo3UyemeaWRw5nMZrI7RTjXX3YiKRC7noAkYkGoOHRFybDluxEU
iZ4jhLQEG3+Kqs5NfovQ8LvpJ31/FKJRn9wrdnXlf++EQJRIP5QbJwaOMTtl3GsA
pPB0giDBo1RCOwljSKWDmfEPmw5pddnlwWM+UG3SqZPrNgGfty9Icix2i1DVM8Fk
eTAcNcLWEfaKToVtXRbP0ckgKujxZBbmU1IzwWhrD2gSiyyIt5604EjcNdjycdjT
RD6wJXHYIX5UDp/ALGnkJVK754RQFyaegfn0ykutHKGPq5x88wrEYDv4Sl9QMZiz
JhMPcviFgRP2jZHxWnx0mFwbt5bCdmK66VNZCDqg+asdDACXCn7yLCbxB79L/+/m
xzPzyDlEZP8AC46r4AC8Ty55WDzFPO5h5eH3b5JuyL2sS+5Py9LZJFnbjq34Hb7R
Kjb6aHckH7xNFF4Zc7ELlxS53yNpx6F6ju3WvIckbwJYQgveflERcLJhpHobZU5l
JvmwfUsl0qTcT0TvNV0Q4f03gdMlpm3uS3i6azrKMlsUgSxgpXnCeL2XWB5IEGVz
JVLNePnyi47rvWqXLmeHSzGcZDFBz3rm3CcmG/lj92/YvflANZpdRNT/z6mkndMn
sjX5M+FY84kTe3NXdJRuYorMdT7vgLxrg1SYyF2k5YodNnruZgk2P0+a7cplAOt0
V8QtGJA24dHh16w/poXsQolrsUibq4Y+9FD8qqX35r7cYM2F6JTcC3Zu0wMXMQ5D
8HYWMqisK5BXSDE/RM7nFMrTWPZtQUD9hdXMIuDjJe55kTj/gaS1bVKwR7kH8jPo
BNKw92kEe4Bn37ja6qNI6vLorg5G7/0tUeJj9Ijl/eQpbDKvIGYzqGJsidBocZKu
H8db247XG9T12eOyz7QSSfNrnnQLYza5dHuNk2UpPVwgesCbdxI04FkrHBVZJS4/
hHQd2tWoje5nrKhuYmLttHrv1cel5dgswS9Ul9PntEy+QCICon90jmE0I6Muxc/X
HGUf2to07HuG52mk9lvaWQ6wq+C0X58m+Mgg0DWpyFrV73ZuwSfZZcQ+fc1yC5mG
RgN4P0fMl2zzZAOyMNaUki8nikRSBQZTeU9cu+2h08ewbIm3KdHAiaYtT9iLlNGL
zVOw7+A6+0dFG6xFiWBUfh9sgOjjfrt/efHgR54QSs8ibTUrr422WWAnm92WBTMs
PJ1G+iqr/SFGNK0Z0X+56UFoQiwAb9E5QY2tQexxxgCo/Go8XS/ZRPjwaDBIuj9D
aZZ2ZWuRC3nFwf5vjk3VU/ivoHRJOXU3aueXejMriZVwaT2YKNsngUUywhiLDuJB
n9UofFHodO2b5sV80P172DLU/crpAVspvLSPIo1KsaoGBiLgGF/pDFzlqmoR4zj+
j1xn3pgGOKO94HAoy0Sq4O52q0jy9dRSoMdu+MYsOK+obfeRkcLM1dPNYtSVUY/+
f7/Ed/NhSjwbB5/MtEPDeMzfL5JWX8lr/YgHxIDf9r7BJKsotyjagvyCCTPuR3t3
ZWwUDv6lNsa5dzd4O31j8S3ppwX3/V223zWYkybPvVyNLU5tQUMYbh66jmvkVs2F
qIv4My6sv8veQLwaALUcTpy5OMfdKcUpxr3h576GkYSySMLydkvXqcdSAsOkWQKA
XaBcB9w4pmcq5E3t4zCTz8wip5Ia53G/4NJK31IfhHN/7knl6Q338YKMPZGKwp93
BRpMk0Ayb7AODT10xAWtUx02x7XPKduCmAQ6EUknNpQujc/gKOA7JOGFGbOWamCB
ENyDjmJHnQhpONyVrxNwjc7FrAAlFIfnmeXk9HQGqjRFvmHekydeT28aZT9My9N/
cveKl1/zsoqi5I9foFfZQM4DJHx1Jb9tqe4HgevnaWx46TxHFhfgIWa2Ixdx5kLO
JsAwp4wsw4+3urOakAxb561H9iMXuINHtb8XB//MxcjZiMzWHvLzHaFFZKf0Ph5T
vOkY0LW3DUH2/ySg5c/FUGy67Nv3p11Zj7ZbhNcJbs0u/5QRm788DLcyCrpUON2d
O2qMQ721RGWQAqn5/4qB7XYba/8WcAUZNTaEmB6BEYhNvwzQfwlXH9E5g9EhkRLe
81S26SZFSb2YHOUOoO6pXo0Ojf31+K3UuPMGkxOoUfp8A5d+vCeQOHF76O6iaMIe
AKkdrUnDDur/gdqLDhxPKkxc+/i+CBgoGQkC/e3Hq/jzr6ZUXjoCXnXfoRJk21vn
shSoshsDtJ4+ut+l6KpvxPUxRot06agLyc7X5wSjzTVdzljx/aE9VDpvWt+zUB8B
ZMuPiPhy8pbqLme9akvnmbAj3ksGLlyWHB/9douwQCB3PUx2cK2BsGTIW4lEf4y6
UTLqg6alDqZETwBYaw8V5VudHdroUb9PQAViVf6gCNuZqVH2FhYs+UUP6btD56ZF
7F7qbXGh3yydxfjnIBi53WklQ5faq7ShCbDswfpilHFA7MOMIEBOw3CxXGVBVIwD
Wqd2nUkQOxFNtUcoOlj2H8dYz6MggKxXoXxZ1GMO/yeok3hL3ls+Q1/EZk8z5CgP
Bma0VnaNTrEYIx5/RumkkHzrH4JbbOkhSUQT/rM9DFrccQybiF3ApvYwioY4B07Z
KAlM3x6GUTqzpCVhEnV9QD4dXkW99h0AhMVAz3KVaNqRkuLd7oL28+67bq5gmwhh
sFFroyBxNghdneadXjc9H4lBhbOY5LtvFGnsQGc0rbXuAvdFx1ocGYoh2B+236MZ
rPOOvSP7ODKZnlqUgT/8r2K1DEaPZ5CZksH9EuazfPVG0UPB3EbywT4Bvj038xuO
Dc4tJ5/2iYPsxfOl2sMHxbBh/o1en5bf16gEVAgS7uvFYJz9ypJ+JIUxxEDx/U/V
cbqwNVHAiDSvyeoqYRAQ4oOhqHvpD0jyyIx9jvGhzKHtRo8J79t1037DFDD1uOGf
1pxwrnUYq1rgSje5JaDR9LcUHN3OXacFlNKzu4X6swVju7J06RHwi7yO7i78WOh2
J5K+fhUG/esHkTpA7wnuxEXljKtOIRk2r+vqjSnsWWIj8hs8SkHx88h37n+GbesB
v1pY3M1oR3ucX2ka6ivIXzELsCgsSshqGXh/r4+v609D8R/zaXym0hig2Vd5nMxa
b6uCQjZswnrQTR/KFASME0RxLFyFsopOHL0RrLNY+3cHyWe6jeXgKZNttSApTEnX
gB2Gq1vWZL14CvJOF/PhFcRZZsweE+LtHmA//MeW/VOkQROJd30wLDvP23mBrMFc
7w//1cKivMPyWCNbgQ4DzTn7J22bHvf5LUOqPaZy9YqA7iVjUhiKrSpQGGaSN4oK
IwBOXPEalDBIoi3cweJd+wYNxmFue8wPTgzwq9ZOT8XYm5SQ/JFvA0HgfrUNHwMP
1oOn4pcIZq6gItHZLFCXBOwU1ZrKdfv8MYwluMdkulh7wjNZRtN1FXTJMVitH3MQ
GZepHp8Td7X+KoAVuIQ/4IHGcEQL/9eGlPNtGXr9qfke6Xgpjgga9IXiispuNWl5
iUeKdAIcHmxySz+xUfXOHdaCxWnmb1drao3eQWDr+LaAQXsKbnFuCvBfcluQNTno
bWdc/HSdvVKLGmxGvN63y5myQeQJSb1Mnd0fe74HQe4b67KcLsOe4qhgDAZkWW1h
+PidvigIh1cs55CjP5MiEYld3kS6+TbxjS8CXYaLRVjRci3fVQ2Orp62KLP/Db2V
A2pAJmkWDug0I/ATNzijSXfoOC9UEPmxRGWb+w2uksU8cUTxZ9Baf1QCEpIK6rMg
3F+WwC7zLUS4+TdWphcdNcuQDkAcT0qfyGt6qibutg5QdlviFFYDnfzGNiUKLPqn
TbuDnifaVr//8JZEHDkgtaNmhrjPvnjvhsrC44s6F/kf/yeqQ7wCKyfl3xVDpZbv
HVrvNFV9aSo9rVNk9J+7wBYX1taZrBqPdtp6cfH10CDxzq/ls3jSTc3p+0vOAs39
4y9sxtwj+kTluEMqRdun5CfYGOzMKq2lQ2CV8usalZgsRlkStGHBCd6rbD44U3KK
xIixaNcNG8fTrf2xCxqluaSJZRlZ6sSPSS3NJpXbBcynjgQgv7N6zFwLtj/W+i1f
zAt51jGWRq8vAcyWTHrvrEr4+wz0SpFcD9iO70meYjUf3VYKDF1qqFl37LOqB4Ze
GlCroP0tICejgHf0ikvoPaJOBsCTLV1hQdgOcc6PUZ4GblxdqdEeLjW1SYR2TD/0
G1jgOesarZ/OLQ2yvGVmyJUISRgpC45Hj+P5Kybxnv+FkAaWu994jbZSZ8eQiQnd
brWjbLQRtF4V077Ad/ftlOTWCq9ImhVwaCOxl1HECQeSfWESsMZrCcvKLjMYsgKj
cHicpWqjlxRf+l+AHj3HOm92lI8O29GKNAFakWYUnGaPsIYOEeArMtjDsau0hNSV
sX4t7Nl/YyZD0hZqOaVu0yD2ngHXwTqX8jzxSHG6OuC7slXaY85OLJ2y0/Dvwbpe
5HbS7A8EDTWtYeRDUgs+RheF6ppEnK9B0XfoBbGd9ZT59dadHoPtC/2M3+B2mziF
icM+IkKqHMoggPIWju7CziIkLASluGJ0Vl9kse7CA0NowzDfD6k7Vn8lp2WhiGyq
9JDGg0iHunuZMXJTD+KJM5RfTFddvHc0n7Q4l6n28w7sthq4KGSQoMFvCc9GlQ/1
fd6vKJzUAoemxKXE2215kMJp3oUSvvlLha1dEPfyq6zjz9MWDl39sXVZm853Yi+4
+Pwyr9OTT7wx+JrupzR09wJyuSj4x+TG/bMZQ+TJmvXNXY1iaxe1JyP79aCiqAv4
FgJjHWFHXmptuC1R748MhhllyxC4pBQp34F19k5+bfAJ3BWRsbahUdS0GBwk6jMj
1+fkEONxOvIZ00Iciyo0eoGi4HA9M1wMVGTB4EUU1sIVP244nLPYinfDt+j08ae+
lqoRlmWrFWgvdJNn4SFXG1zqzpEhTJYwPLqTQuT+Ru9IvfQcv5QBFWULl0nmtEzR
1myp5vsUbdM+hZsStH0zZyldjyeZBZxXBsEFlGE6cXK1x3MtNolGQ7Q/pNKhoxju
1KQPo6PohyK0dw/iRn5j5ezHuGKN5f0tM6hjIRQeE7pKVciHmllDRoxzVqyG74aR
JrpaEiJqjXafmO5KeuiYTvYKpHJRGKRRJj2idyM/EVDlr7MVSkJrvta3ZrsoouNP
5HcWXX9hLxvx+qXXj7s9jC1YWbBPqGhjbahjthbU04+U+RbhV9fitBSUmhr7jiyz
D0Lm0jN8edXlyt3yE5RuXoWpMQlKJl8jso1XXMWBS1g53BRl4cVjgH+Z6yFKiplm
NOOTpkaFA9cpCvEeZUrrksrJJBjNAwhLriwQP6bZiPp4mY8tjV1qttIZdICAk9Mr
D3IYQs3QU0oq3cS4qfYyxm0QduQyuxj99zn+If0BOFQcc7PU5rYsEspM3oD+qI+8
yGrZwOMn3U8bBPo5geBTvjbBzy1LHlWLBhGVm2Ief3wO0+wQdcURfSiUydLJjBAk
nJniBFeOMV0c5s8GZZYfnHcH3eokHd1tEIH5/5lsgUKKzhinPGWC93/NEii91KIJ
9r9gHp5pvYEcv7conpNQr59OfOar53anMbmaPerJmf+txgl6+yL8q23+ASBcQqpg
Fz7VTndHmjnbaW2d6uLCpI3rANyo2aOpGidfwHFO59uln0pmhkR9twQmrIrLlrL4
ntKPkhYN4PsirSeQfQBgw/oPd4O3Dh/W7EgKA1J13UpjB+xO2UCYb68asu1hISq5
55rUKi9wFEcq7wIZT0mdI0DOkoqy9Zd5qyGfBnpyCigYrV1cF7kScycGMTwl4ldI
pkPdbWkoZ+n2+TBfvZrHN4Et/Mw6HJPmRFou4wNNsnxCq4qYXHKDE9f3O3HPa42Z
lxotwWuhe5DCNi7htLJCOdkBPoL4nsZoiz/r2vd9hZC9lJrYMheiGu1YHBb93+b5
fmClcFtroYY3BN4yuYkCdtnbSVg9RIFX9J+uWzjWLrkGGjG6yCtyXda1jeJ0IF2L
XRBj8QTpBAS7ShnAQNAv0SxG1nmwWT65eM403Q4gF/r+XUPmBabhtqt4PF9eaj7H
OO9myS78hKZjtUun31Eb/VBwewQp2Gg5G+CEKgkAS7XjrVs01MXwUpUSANLvG7K0
1XaU9b9j1PhViB2Tt7AL03U3L2WhM7b5fxdIOed5brlOnpC5NLKvueg3be+LD/uU
goL3G2/2ia1poqRq6sx7U4qzzYb9P2STw4nErxCQWZnH8hN6rOk1A3mj0ZZ4Usu3
Sb6monY2qfpe7z0u20jkoz6KlCAsruoOXlPAl1ZcvGz6tWaZ7maFQrv3adOvKIfV
ntchjJ/3NcSBZz/XvjzfowuWlQLA89z2dheUIRitaEPX6nj6Tlk/LHHUgAAjKua6
3v8eELO4vZhTaWvOcjbwVjCJth/0QFTq/JMZBLkLLCEUC6XMZv/bmjD/I6r5+JCS
QMOse1eVRCcN102kcn0HNj4V1/BOKUiLG4yEZQ5pP+II5DGTrvUiWRdN2ID4VtXk
+DPxhyx9zE+BGA59d+YOBKLja+uxDE/T3fNNbCEh/WCRewuzkii7ljxdGFK8oCTJ
y7t0Q00ic1iWr4Oq/Z8Da0cvpGXQ/sJoxw1olF1895E1aRqUdYUBVVPCkpjXvTp/
N1XBoiLiKM9Ufm8tH9VIvwZgbEwmDs9wpbnlulvP6Ka7uLZIMBRaJXmP3a0Ne3fI
y2zND4X8MEcWWQehODw1uVunicMwd0iKrEbcACMQ6azQ3XlBzXLvvCX+kbW9iVND
bkDfqveiT3hOu+kh+AZWMDWhSCr8DiIGdw0sqcROK/HinGcCqyuiIzyEf444z8Gs
S81FPnfgbNZSVG2Rsm+KsyY05nMNPi1c1ICTpLHCDyqlGTFxZPUj5ImL0bskBD1d
JViiz55+8/W6ts/2dAQQ/ltYDHuk3EU9HiV8fBxtE2v8yAZ0Uje+LBOB+DtjwwwR
a/0sRH2HvvfUq9sc0JZRZsKscypElXYGSVFnCtIsZq+KFDfEjeLeqYdc2vQuhde6
0tSBrJ8BduMNDBSXF6MyaoMzo0zId0ytozoqjBE6So9YA1YLoc7MfD386LxR7GJt
XtgIQi1z+Y5LaGOABxNswt+OhFuP9qc3EQpH7qvGqzetI/PpAHwYU72DMFuksRLc
hhbGbUUw7fJFsW1J7HSBH6K0W2ceon7K8U5zaWSQREdaUZOISG2OlDmoYUqt+eL9
tVj1xAujM7Xhontvgd4fdBL66mtEQfLZuEwFj8UQZG88ktDt7DNzw5DEHFm/ed4x
LX16HRjVHep6SG7Tirp4mqgJ+jY7HDt9K7Y0iPCGufDb3sEQK9MtXGs+EaVsFZhY
ViPKrtk4HvcanbowEVUZxnnf4JfFrOkz55E5H4nPGH04SnMzPEUqbtMofindmtdp
tRDUfhDYYyBM4EFv5hGjzCzdi72drl8wwx1paSxSBFMLnj8x6BRgqzP2ItLvmc+Q
PyrD43VrpECpaKbcoseNsl/18VAJBK6JRzCngYse4kY8x0nGLY4p9N0/SMyzwuFV
joPwgYM0pXiilN37haoNRaC930uxbhA52+n6WhjPTgjFFbKydmW3C9oJTsz/TRNl
ffuYfy9nDILcRNDNuVVJzMqa3AjXE7jca3HmscoYdIs2pa66AY3s1jDA3jT3xNqr
ysmEv/RwLIX0oxeHbpee51Dobr2dpTHp1S9TGDT1bzRw+RfgsdK6r9cLa3Lgcs0J
jf/BfOUUdMVZJ23cMntJglNYSSILKZdf0wBaL5VRdLlVCfk6fYL7M9CObzO/NZjv
bmyNBdxEMO4qK/Uk28zVqEsEstiDpnmwsERzhkFSGNq/3VeHSxOTiVlAPcHK+y8e
FWtgUiv017c1gEsnxIda2/qb9bZ7Vt+LumFtvULXiozvun/MPFBIce6Ds/4VjCkI
sMpXpIVBWKPdSAqQQ4iILrN6EO9G2wPXpJYq0c2iZr+eDUqJHNH7eNvJwFaHgTRU
mgE31iS1IMPpkuMP+O5OWLQrDoWUYv7uEdIKp3DLvHweQjeYVHOiq4gMSX+f4yRD
lLrpII44Da/cFKbpF0ZCxjyevbZJm1RIZ6TT+c3sUT8voP3tj24zyCjKjEGTGrsX
ZlPWkrEly0cvn4ZwTYKLKh6vaw7RK2V4bVq9GiHD+ayEXVoru2AIifSIt8d32tWZ
Onv54fTjBTHF8D1DH/19bsV90nq1jkeLCpMUXZiEXl1mbYMclb92ggLTu8jGR+2B
Ks9E4GNX6+TgRU6wHPXfpyUWxCTohCzFXt9i9WDPpQCiUJZg1SHZiTuV5ttHEyXC
6TOXONrxnSXK/7rd0el3OdyZ8U7Q6VNx7/ti+vmFLI5kv4RF4pi6d1FCZ4i0WUiF
RTWkFYoyURa3S1Z+NLiqIEKhPe+1K6Fb59cZRkua1NEmxyNnWZqaLovUNoILC8nZ
b8IZaWIkDDu5mebRPrekpzskVa77zYscT14XGxpJI7CNCwaZom6Bk+sEt3gvPH7V
O/6AK+tX8Lx5jXZHUUnrWqs9CkbfUXv35c4Y20EyS6zZWwp/bfWES5OQ/qcUMhBJ
nGNaHBehaybBdyWzr1cyI0HafiienJitQfhxlwcFXtYf2RjEl6h0BbAMDq2gxrPO
Qf3CWHOv+zO1nDZVW/v946u1OiEV6NEVXHFCxeHuZQIH1+46IIvO/dYTzBE91cgb
Z/91Spx84xu5oeEqjBWtJyOsQmfywHe5T2qtlj+WxOh3hoUjpeTeDN8lmBxSHvid
x7eciVQEsuRXlZ1O4aiJi+NvfWh6YQ9tgml8HlBysFSKmkcscm5Q1SmUNARF+pYZ
r+n+xqrOAFcIolp2jgWjmrrlcnwmdHDoHSkh3dz3VmJd+F3pB/gUaQ63e997k/9V
6wxwE9NDb4zWN2/Y64x7+zfM6bBUBK5OK2DonmF5WHDqvEg2YQ4RBu1LlR/OpIfU
tXS3i+5NM9H/NJu4PFVGww85DoFj/GMsIewHNlIbhNueLJqo4Hpg2jfAULDSTRFZ
c/Ggb4jNMLBd1IVLe4bkUK5zfDrJT0yyVgs0jrQ5SOlCTrjN1qTy6BfHUiNldQ9D
Ax/l9+xwu/49yJfCwxDzLxF+JB9yvo01K8PxfNTzg2MokQ6Y67DPvOWMS/JUsuca
tE29KaEWu7KNJCiN6LEMVpzGxBSNT1xsey7iWkEinSXXFT8A2iWKVjjbTEHtQxTI
qHX7HeUHS/WS4L5p4GXWs+EekCrNqFHWqOz/uLUPGBJ1rymU3K8kC0q3Qp90ju9/
My2SJc6nej0g9K2a3FhhERZq6uZJhb2jXYEjV6+uDkT7U4nFQs2pCHIdSX7FdFso
EcIYC65k9zujlARNC+yMz0QZbydRqfEHqmKxmG6GaEXZ0Iai9ZuXNNT1v1aqknx+
sE0uvPtDiVfdRKCjDSO9VYR7NsAqpDRXD5yj42KcxrYsU/NE7XMRtH+wvOxNWNx4
GGRE6TRtUKTd2cv630Ao4QDEV40RgsP8YJMPECy7+9H0QBzFVQQKeESyTBQToUHL
dHH2EUutcF2mIpzhnLnr99tNz6AkXVKXpUL8R3H88uShvSjx3wYkDMfKH5R3tDdh
uminDwfMFL5+k4WiOmIrl40mHbRygztQg7Q4Km+erHiNDVA3hsppPOm2pnHc1Mvh
GTdLgVGzI4zi3ap20SQ1qCUq09QP1kp29JheDfeHnVTKt82NoUxok2oFazqzlrSB
koWzMaR+xjXA/o+LDOV1Ge2xe1TCzUQpZ6JsR/p4Zhi0ekCcLz8LKEZygXRTeMpU
qlj+eRDmn94m7eKuCwkuoipSdgnkOuqReRmNPyTp/+Z8mBnaJWLLxpzdfs06zKPj
zu+TU2lygwddBrKt0nCifmGcGBrmt1zb9edPzlEItJzz1KFalKOunoCtUKEP8PXJ
Wt8XJQcDyWzBZPrwryh4LrKYd129zLdq/kZp8+hEnvCHyHl2H4p3fjKEUvd3G8aD
KUlaKRvrC1h3E36UPMcb+PhMeaoj/x+31XBGG3zZ0jc4eSt/teHQzdx4A6a6krmr
fjSTfS9KdS4nDKo7bkzGPHPkZrV1KQgnMf40EhsEatuGwrNm+GrCt2nY+OvCKG9g
R1OZzpuDX8WMenLx9OUz0t50y0FaqaYGm5iQe9OTcyXemRGGT/GA/MJ6TKaH03In
lq8wq5SQEPZ3jF8PBgjWpHrCZwZNGqtr5AkfLZiG5+T/pZxnrt5wPUdXfZFCBLcH
vxlzVwnr8EHvvFy58lZixdXrELRF+iU0H4GeStSpOlYEPfUDHcEZNfNV26F1mGi7
R2C5D1bLK/bf21txDU3K985RJQHVhR3vAFAlPGRTZXhXDO67XwKknJm6GJAR2Gce
ylgkrDKPVlMWnweQxwDDOujzyR+olrx9pD5/71QXh6wH/9VGsFX2PjfXuFu4rkdt
heAsnIeO8pmP29JJ4cfK9KF/inqN5Elw6H0sjaK7A88Buz0cweng/SNekgzRczD0
vxjh6sWy+GywZvdk3blGg3CjuUcQe3J6YXMnrTHJ4P8tvsmgF67UalOYcxdLZsp1
0tXWJpW84z3/jpsid4gqGybkg7qHMxJgGnpZDQhjIkMtrBf6q01JNV/8+EZvB1Ge
GnDMUWl9h59CY0t2Xf/UJW8ovgBKQSHy/Kgs+wDvw65hjtv9p6fJl8wAQlu3HQ/4
6L0a8IzAyOl1oule/xG0acuV4w+Vvx/vxxPJk8sJSZmUHVdeb+txPs9aupS9s7sn
ucEyHzhxrf2AGZjKsAQDVXGT/FzXNorahY1FCtLaExpEivbYdRXdrQUXaGbUfaPn
l5OM21dYmoyjXMS7qr2GP42XtJppE2CcV/SOBAAdMivm8/2V6xCDcs7IZ38SxxNh
l7aJwpdlDPEQNk/9uFLqEbPyONsr9gnbV3Ij9yMrNqrJmWc4y5H83FlkhGaU19Xq
QCenpkY3ozo7QlRq5Iq6vgd2Fafa3ciHWXHR3LgXO3yTvabu4QBwoRfeT4Ottcpp
xr3lINQcT30BpEtDCOemcAIzd9pTeJKc45ytydUk0nRpbqTQ7KllTKFefZGba/ZA
6NzxUBlnKgq+K6yE5dshxCicMVhxA3y9kkYrQy4oEAioTDbydF6LFLDGXUxIefvd
FJFAtckCKNfOvSn1yi6gBvswOuW1nbo++DkFjDPRYkUfrWE3/z/m+M9yKOnnfGm+
cfgnW0MIUgasvwIatUmlTrZuRtCxyJHUCGMjpFc/OPv/3V5RtQPX0wlsbKo4SgYu
3forkzCRrtpQq6Q8cgohHTnpTSpy2hcKVu3omXCDNtHXLly5bQh0Sh6fgUvBAm0X
d2gQ3KFGIhTk1benV2d6ybmn7VBcU8XsrLp3F+mVIBOpdKStnR0FFgM+x4o41Pu2
cAVNP444H63eqt3jkMXPN3FM1BsgljMhoqeGepdknQi9bn+7TZDeLvfk8azMqMSp
UPy6l7eGFIyrGVJZlgK5l1Hvk889VHuQWktVm71zrsVmz+ocl6V0vK0UEDC/BxLg
2W96JgurcIXZfQWlSsXrHa10/+JRzcXGHI3o6gnqyLHVIOKAeZX8FT6n9ckXL+ev
VnsNT6ZIe60V3GLaraVHMu4G6UEa46CI4JSH7si7CAXWFm8HgpJ555zNEL/Wmv1K
mF9u+yCNlWsVuysJ2XNMABkCqaSnKbLKSvhJ337bMKSCPrHdgS7ILUB9OZiH4Vof
d7PhX/NJRLrcxx6ZzMeYU4SSuNpV6+fqT3yaxGRDiQxDldsdBoXqL6+E7sCcnGle
JXGoRbErCeTFRtJl4Lt9Xzewb8hQEFcCMIPwx4mWcIAq1fTx0GN9HA4vGsk6QzPI
DBiy3KCKQNdFdsMoaSimZglmn+ThKUJacK1kIZrPysIGIDZBDq1r/V0qAXg85ego
fnrhP13wO4MO0I0dQIuFhPnJe7W+OptMJTEPwwevC/HegNkz8jcAiS1LbLGu4eLE
U4bM4oNDrxnWSjb8+tQoYP2tE14dLVokmACl3iEaUak0XCtSYF0IAtKWRiwBBxnS
lNd1qNMGJefsK3EvTncxZz+dFVSQS0woGj6My76onXQDSqjQcdKgU15FjSL+k1KA
mi4rt7nGj6XZDAWhZl3vpEqbL3VXFAnYJjcJB4UfEDmNPD23QLWvaNf+f4PYL9mS
jM7sd4XPDl4n+An7GN7KkOzuvfnOF5JDcSaKSxe/G+9zxBT8iGpgW9usXbl26UCZ
pZk61coRviyMSdhcKXpVj8mYP0fZzQ+YeCfi8sZyfoz/7WRmZ9KkMbPOgcfJINXQ
xf3BEd8E1GphMWabc7joaz8+HyiL5kiIOD6v3+4IUBbNwstUPci7DkFNWW/i08p5
LWNV3xh0BrQjo5XIGd0D0DzODoac1loXUfzGEkAfAzqyXgp2lltinplyCKkXHh9M
oEuEwDGtQbEikVMmE60qcHrgrfYWq6aCVUPyr9GaRPCpzJQDcvosOT5bA1c4PmLm
CKeMdhOgEbqi8g2TjcuTdiMS/TcjFDdmAwfzyYNuJ7A6KlV4iCbx/Ik7cm12U4AY
YbfjsNnX8tS1vkjfgGhzot8t0F/X8hz3/smMmy4EZP9Ma7nl/gSov3FMgQUhx0Sq
S2ZROCrjc6vJ4byE53REsplTfDvc8tWNAdg9iJzW8bYmi5OuVhgF0ichJc94sKAS
yutVkT5EAvT03+RUBvC9kmYo86pRnzgMkiDuQQ7fngDY897brjbyHCBr0DdHsJYI
gimtgp/izwOJy4rA5gRMbJ6n2nSvNg46Jqfwst0cssIyuRJGq63X6nRobsgGXRBu
EP2sW8CTDXnvP1l9BNg/b2yDIo9938WYaaPYkxoR0PjeSrzr/SH65dqswNTvWYaa
d05wHCiOVV1H0jg9NHwk6M5AFlcK2bZZFDKp23RwJvsMkELhwNEob3yJZSUHjPC5
LYcU/96escMbDz6jObIFw67IVeej8b4lIwz5ep45rhvvlNbCyferLhpBTiH08Tuu
cPFn9JR8WuAb9Bd5XSNCqZj0vhb0UbLRKDtizP6Qu5xzYD6rWOUyyzKybGWDaoZk
U0+R5epgTar3bX0zJm91lh2n4f1F3+ywul2ZeOOGmUn7XbtrEfNOG31z0Btafaoc
UvbgnYHaAM4WHnAICZ79ASmXmJB0y+OKT0TcxVYHD6vrUUxJmh06bYgEn9CIRlhJ
Dtq2cjvJSuZ34l4m8Z83C3a8wRqFJ2qESCJ36Hx1ICqRvcMYC+rH6lfvsBDTkCh/
N47stT8PKSGJQDjvUbO+768eVPWe6buPwVDRflyV8xEzusi0gJcsFIq8k6FFiSII
TeYkcGsK1klzDgM3wSy/0l2CAmUo9qPUmOzu+wyW+ZQPVvzJptGR1qLFtO+9Oeer
BHbDMi/8y+xKy4VW54J2fKBO9J/O0HIBPi8oWqQEDOsoYqfZiiptC/gFZ4F934bS
ZxkRF0VYLuJNE6AT9BWjyT+0KyaYMaYn+6pUesAsx28sEZ7XBJzTM9XntaVkSaq0
qQlK02Uuy15oqTbboziOpQZX3zNDCiJ+wIrdyaVQIGNPRj4J1cRVGjtU1ABS2Beo
slWvNSAngiMNf/o0lqh2rPFPPypPm2/hCLEqNKEXYgtrOokxwG9jxoJA2XZgvLmX
gVTNTmJ309jQa7lQz45S6rRhkwXXWktaGfFx4BrT0ZU1NbrYHLhCSIn8E0TKftZZ
r6nrDEE9+lJgijuSlLLTUmpT/6sEyPkZolcB1onE34GF8TxHM74Fr9MmEdR+Rvp0
X9mrDuMIE1t2rt61vLyVxjr+lOzZHPgGIgzK+wX9CAvfWjiiSGwCrKnKdPfdhiFf
MM7sVeTqpc9QCBZXNFmHlJTfpR04K5lx2vxAjm8Ljc+fhJoly8RaWPVu3Y3xK0Pd
Gz6qpVioruW3o043qeZUZL1UFmw5VubaKIRLXf1cpPcwP3prQu7BalMekjXnywcI
OX9EDVeRwDrNPzalJYzFfReZJ0n4dwChaerCmdLr81XiKpiINWjaVahceWFBJu+5
tQLvjBj9daZR5N49ATzCb1B8P9Sg2fa1rzpY4Y8FuVz09hOOzu9Yl2vEpTyz3i2I
zeNh9GkW1i/SvMDrfMNSZYskXTjGcdCDhnQnT7yVFTrCy5fuM/2qePsI6b+U+d8U
4AGJD9oM2wSfB7Ioic2kB7bAyuWSpMc+NU6Kc5B7Kd8Z058tH5ItlNhE77vdpA3x
6s6xsMJxEN/ne5K7pFlZyAjAlinMQX2IsSZOit0d3UKlNuKMTeOQ4Y5A12H/Pp8i
3vpiSHvnSaiU4/nwgKr5d/ttXWE3UxpMUmCW6oCITFGrs6ozoP+L4T/EqeCH5LlL
KTw8+ehl5z+gXpSY50qqQW/QW2vJMmW7t9+lBb6PLb00odVgYyVFpq2ynQLEnEpR
00zco7m2Y93IqqSNpS4o/Fp02u0alcC7RCGHnqZKWFtjnOQ0piVlUR/4DToBGvLH
qXhd3sb9uH/wSj1vB06MXZXd2WTZ0P3MR5nI2dkZxo3bKSHFz+qtagj3IjUvaOsd
6x9GXTm7boqu3HCpjvkDWluLGWhbzvsj6GmqRojKGMKKqdz6KmI3N6Qoec88uP8Q
ak6n4dvvUy2PBFaBv0Jgq8mto5swCiJd0+E4R1Yz6dDJurZQOsev2eupXzsx9AWg
AtFyRqJc9RKPkjucfiIqpCulAa57zvnm9U15840w9RGniTTJ/8eC/3iyFy6coBaB
Ph8kcDSqvbgIVpCXl3dVNdX7svVUCtOKLLO0VA41yHz4kyJHGP9t9Y2V76YxI4uZ
ffLrV0jZXuky6GrIb3XOjzB9LHmDMfv3WlzM1+GFxcfkJa9hFsBO0ggLLDxYBLoX
cSWLLsYGBuh8KpGWbKZoNtv+wPcNR9rnnHCTkBHZMUbxWbs53eEgYWX/nwsqBE3g
DWeWbeZKsg9du76FYkdnEA4rLOSmhwZ9k/6A9r2OxP5q617GpNGBE6Z5yzZQmT8P
9/BNuPW6W67H1l67aCUicgTtlWmuyazSxISXfyuJyvLEGWrMMYIskyARd10WeReW
ChqV8FXcVCnnhsG/P3fcSNRECXnm65kyepU8/6sXUSd6nRLWnelB1xx+4t49LsJ3
nHbyqHkVA3+paPdrjZTvBh2AVkVc2GfPQ+hx5ZJyz2ZQCCLGx/vlVZbRbp8exxSW
q3AndDyJlGJduRvOO0qVUL/9BlXpdMeKoVSSXV7wMpawDhK+cV6iBZZYqd+uZoUE
U2eT2lJkvcinakWYqTXa6O4GLIUGiD1t/VIogUZP2PAQUBn/bXhacJpznBLy80rk
Kh5n88TjuTW8+2xnFML31bsBqEW1ErTQDQgQG+Y3JjVmF2B+Yxg3yiMDQ1qaBUsB
hdHkX5sTapDyUhgZ76cBh2m1w1Y+Gujl1uXGnxrxQiDHCQBUb0T+faBEOOTb3bBp
oDAKWp/7xiLe7rbVYRyiyARoRc3Joq+ekWP6SvwKvZT+YQWOo8thpFppJBjIYZYj
d2kUEwrg7A7n+KExUK4h7K0xsRY7FhLpfumdHzn640Ztv2VSqRJiR6LZCJd8UaB5
OzQeFJniIG6haOZP5h0oSXoDMZ1OKs+RFhQQElNJjgsxLYp8gaP6lvXVam8v9dRy
YGx8GzpjXM4j+kPpYJZQFXrnHNYPlP49m2tpBJaIUcOEvrE8as1j1YhaDzC6ALkR
C7iLuajUMWLXEvkcfhN9rB8V8SdMhgnjKYzBy+tI9K9xI3uQf48PcqW01w/dHvlC
tNwpjKD3kO7jK7xRSkqkWWU3dRKfN+lC93mVWpXGDr0tYYaf171twIGMF5vDxtVE
jTA5EO0S8rXsKyiMHy/XfnyxPf1LQ9APZgsjhQBR12C3niXPeNc32xkkwX73fy1X
Dv6Nq+7rqC2l/jyDK7aBKJYG43tpaAbZLWXZFj7ykJ79JNZ6GE6j6r8GPJSg7ZFR
jWw1t1CZ0Gh+LPaBaKawJsYVwqeSi49dw/qJ92evHG8N73nu3mklgVBPkvQ0dLM0
76Mlr1LbVtHOX27pbks3P+6bXA7YbOCWBMvziqGWr39FvroZPs8uf3eDvAdU3Wac
7nk2tNhKsQ4GQz1nuXue4p2VerAjH9IO5zytW3BKegNy5lDsigRDF0xwJR+sf/RV
prkQ0weDhT6mpLZ/5UOo9LGNQElyqnzjlEAkAAGaPmwkct9U3DNJ0UWkZNCPxBAx
z/SkjTmLD11kTODuF2fz9SK19LUrxwUwIe3yyCEJ8OrjqayzsAtLb4jEPuBsEb7E
WNy5r3RREQo2qzCBXDtFAFYWxGSa/1s30DtEY02AYVcqpMHg252sVxehe/EjqK6Z
D+7Lab/oPyFX+DpVPZp22cvfPULw62ypeO1785yGjBDi9zME+vDvtq4dFW64xeF5
3JLZmxwBGtRFiwktysfwvTs+/jzMzW8lUzM850LgDa742Ufe2Kr6/lU5iYSxGSYm
Occ2RY8ZXMwNs68/VdZGhDfPJz3+VPI31jiyxRBFIjoc4SdjoqFK2CFLnR0d2d9Z
Abjt6mJJ0MeHGsdebCm4dsz2bx12CY0iIn48Q2LwnZq/FtZuHtOI8/MsfdUHvFoj
sxjo0Spr2ld9OQ4B5eyR8iH5QJ9ODZPo3ZMi0k4IA6YmQSVaK29JRAdbdwQ0HVFZ
uUZHY+UfSVu/ExnQ45uKot+lGb9whMCDKLD5jR+JhUtw6K5k+BGa0EkohovVfifN
IwCea867zfn7V9Q3dHHjDWXUsut6uLGNBWs1EqnpGkEIHXQvvrmDRg0aUa71zIRj
EjPtpMrbmhjP0yxeBTSr2k2WhHSdVezp2AG4LBSWzED1AdnLObQCPe3TCXCUhwUM
ZaZQtNmUSnDW39eEbqfaO03AEswiPcA+wVIgG0qUgBUOrtEf5gxB37HmEyRQa6Tj
lB0iMezurkx0X/tel1uOZ43SsLwp0bfgg55HFSqYpwFp0eiyJdIofyVyVLQjhkTu
vfjPQxYl0ZlLX2V/fOcA0D7lBeCR3CEiA2EJ0wCGhscGPpGrf54cRQUNKduwf2PE
5VlU1lgFalB2c8IAZuhR7X65EnNGZLt2YxZ+bSbxszwauyXCW/uEowr4BLZ4L567
rwrGyoIp8pPW6fmIK/dbPsRxQaOtmxkBlocb6PRvcmuncL71levkfcujoz0oxBlk
POkXQexQhyoU3iU9yHIEMLhVckOVwWD6W8MKOIgsRYzJ9YOB6Zp1XURDT+h6Bgko
xpWXlVg6HXGsAlBeszJYMlEzudqAZs66UC5DGv1meGYyvRr6alU40wXoq2Hi2W0w
KPxaFB2Dk9keN0P+pN+Qu8V/nKL0gM43mYfzJV1pvIpUDozRob6SjHb8vlZo1zvt
OW3qyF2rV+RZ+QsSnKWp0H4NlXy7z2WDau19bSnOaWlwI7qRbqy3Xe3dPuzoYMvg
1jjJC3XCcqU+L1TEs+hydxzeEJ0DhLVlIEFgcj/wvAaA2208k/i8+Vg5Tflpt9VX
DIZFRwJJy8Tsgopn1xfyHeXiK2nq437Jb3+hA5smFBY+39PFQm2gbptpHfPy/cLu
PDnC9lJSwuWbmr2Btv3VhirvfVY0JEwg7FijjBq0ZcdXp/tLQLSkbXgjWFtZUNy0
x+lkxHtgE0Id9rgno9mjy2uT3npwVp0sMMSUffw5nLJCrq2+HgWhnZ/Qor+9/8ph
mh1y+8C3MVz29trFA9vmxk+7H4Ik6unvc0D7vLKZHpQiE/X4CM/HVmXWwXbZ9rRH
TMxr12yzV619iIgEpCvcdt5YCakyZ3zWTE0U87XKDY5VJIIpSOw6rRuKrxKW0zEr
bi4QlLVsGdwZ4MGd9Zo2NaflsgJINcI7nXgSTHuoSlGEs00BMK9u/PAZ4ejOmWIU
tTpWOYIy3Rs6yzONPTJnz7qHTz5wYxcipkNz1g7sa6bKawXNg5EA/Kagso17qEfB
vqbspg883NpJpP3E8folNyOAIccqrJtVti3WJf2gu5UQJL6yK3LYlwezDZr67q46
G4Xo7dp/wry5S1vSkvJwhCHiKAtPFN1wxgnJuDb9+am5w+SSTw01qPnbIIH0vQs/
PDEer2ICCqjIdfOMsUvMVww+43pqX3lIX9gTw8FPP9WoZNcbZtrd4Rp5RqWLT1hf
zYyqkF/NsSIB7R/qNKsZ4t8/aEp7EEUq8EawUtyRHgeZkB3JYek1Wn7Z1QhFqXHH
5rVlEYk6dNmkKfazHZmkkhgKlVroUsX7KTxcNG/MCoo1l6iqIBGuXbIh6dhzyMKd
jsPB7aAkgXaOkKFIsegGUFGA+drpwHEKVaI+umyj0HcalErjuuxgVYW2UsoXaTpo
MzdSaIhJgzjIDPvY2ancEKB+Oi+yWunKJ2QrOi4iCA0WK18WBUyImIftBTd7MLml
sfmcR5a677OAE98Xmp4nKBQ3FsQd+HN2OyBp3B0/Q21YAOsRhjUjw8lMWx0MOZQs
L7cdPoWG5tfjshovHFzEEBiVGu/fbYUd/KGEPjGZyV55aHV6ZHFzzZU0b+leI40l
WMgLU8xqxu0MI4QXcMLCyqta+jHL7gY8duqMIk/ef65csNnAYecm0caeS7tX+HhD
YWS6PZitRJE/kk91Np6OKDO22rQ6GB/6nUJX0y6FQFT2twWERPc0ofJkSQ7Bg3NY
XzDQYL7iF73kVBtSbQQvaREGIBuie5IA148wYWudO1aUKHD9ZezHJ/U5AgfvgJ0T
wPq1R/coXivliJ7S3B2CqbWvSQDVPYAI2HmWa0ZUSjbeTcbnBYGPV3LmOnZh4/sO
gfjdSXIG4M/pMgqWA5bR4BFlHyglDyLG0kPPQfkOkPAe1kfjgVJRICK0DP+fhyzo
5gMMLX4w+kr4wyr0MUkFzYQ8nLAFsDx/QhbZ9/nQ4k5pw4UOV48i+icSLuSMirTS
Dw6eHHNPrTAoiBrrei5wBuD2In8GQpv3ZyajMuZpjELLWCVX4t4IpP5VuJHzho9N
i4DPVEwOgISRArkWvUOp+oL6Qqkx17vyHLvaZZksLK8ngox/CA15WEskYdNKfFGh
VfWgs1yGU0zvqK/Gq85Kid6XOzU0HL9Uao1GflCNb8PLML9Y9/0LdC8qepCfRcFK
E5L3Onq2r3/j0PFjYwzXfD5nDVT+x+ui8HY4Rya2JDPnYuLNSLJEu9rlJ4TuF14A
Cc9GrGiOzbmEo1pHMbMcBn5b182Ty18lJ4WWyQ+YIvk19D9er4lhCcJaN58eicag
YaMlCGev2IDnlpbEMo1YtzB7s6EV1EFrpGTgG9U1gNgvWzVEC7p8zMSwS2TaHF00
VQqC10+fXa0VvP6liKo2QTNcl7XeNE86dLXeM9H0CnQJo2Sxgi9bgWe8JL0n2HY8
o0GbVq+FWOslnvTo/RQu0NIJYG4oj8Rq1lDi9EWNkAh+jCvQm5d5fGrhu9Z1I25p
zaCH9S01zFAO09W+pCbdmTNHfEKEl334DWMVGHtZhDH4X8e3qNo7eb4Yipg/ZqlT
gUW+Eu5yXM86pPECJj2ixiVcjb0YOFyZJl+DIp4gxcIO3ZpPp7Y86f4/IM4QimnZ
Xz1UYUA37+1SLpPeqs20b1uEuatLZttDn77JC8ZaUDfLvL3tPpprfQyPO2KBr9KB
DEepbWOGug5tzS7vnUJWpJFyC8QIuEgxC7e+l3EjH6S+pBDN6KGlHi1JL3EtR4vD
MYpaY6XNF5DxJhCYN63sbsP735qCZSR5dxjsX/KJArcMv6+bv8Scdx5G/yos3S7o
ZPpzMfm3utA6Ifm4Viywp5rqDbTP6qK4RUC6iTU2oJZkoHrTr+8y0vJT7wFGOvu1
3tjRDLsDvmvmwLMN/pSHvMRxEV3rXa0t+s16VLMjOh1b46GKHxwymjuva3p4MXDu
L5yT6RFBxz09QwnGJVLOuoI2CankvKP4rL0NozgB/WBkkmir6817rnlcJFrT/Hc/
0FdQlByQ5eEmJufuzfEqaWCGR8va28/d9nJkvm1GHCNSJRO/czhvnKV676rUXAxJ
b4gydvor8uV7WlgPatxJN62zqikM0BTiKYJanX4YCwCgy0oN2ZzG0kL2+fqt70r3
6ra/9qxqzSOlW9c+9bN/JdbCgjTFmx3fgFU919DZd0IGuvbAQ2eLSWpMjrY72loe
SW9sIiJMVY7sLIa3FmKWUYgxFw7tpTZVx1qpdPQsThn9bL2ahEwqo209IVgDusFk
0UIqC6mtUkL1HFD4r37+JJV9mCdS58WqyuEWmzUBi939qjOEK53BFj9w+AhM1ikJ
Clg2JlEOUDVoJ/UsyeMZTHijKTbk3qxcwR8TPBzUZ5n6B5Z8av2nh8SQQUJrNAT6
5YJPy2Ett806t8BDirACpMqnDCe451/mza7qrrmgfVUNQ2eFLHHfwtpJSQp2inDz
QTWMCF4kKU/VdCYW8jqcTyQq9ldtqgc2dfpcccTfGtjRDQ/oizKxHNzfqB+XEr5H
dmWtjRXbHa6d+XLE7Plm79OLnf7KKZ1/Wjl8efauI5O5ywS1FCNDzJCTp89TAu+O
+WemvhpSi7ip0yX07GO1AYLWnQQ//5saw33G+sxq8j7aPwiTtGKP5AN2FVSysaHY
bXlMyi3xvni9OuUxXVGtfZXWBfNVZ2kqJXSCVdyQg1D7GVDUVyXliYZqL7A/1arY
sUqx04lWd9mKpYIQrYmAcD1iw5RM5xRivGkI78TaqUn4uZ3cXIibvtuAKOPU3DDp
xYxY7+uo5oFGKlPIHUFgYpaxabHVu8t71zvHton5rJX+vr0vHRG5aqz2g9FOSZqt
m1q6HQmqLqRlaxC0kfpASmgsqSL4JxvZHxFdMssqE8FFX1MPpfXmPwe6JRo9OXEm
iNZjfrcqWmyr9KkIC35l2j0iQW4cPXoWHH/mlXdXOmHo2U56SAJjk7DamrGV+BHU
d+PrrU1gAGJWRZAMkFbOV8Vv/jd+QxcEd3SAkSo/pBNbrcpeqiHsi5PRNeBpox/F
sOeJFlsWEHS2oCfbpOx/OWnkwOVVbr4is0El6bH9vTyGZvzvUWLWB55nvdFIg0iE
hSjKgrekMT4/DzRZhTXl9/MqFqJujFUHcaxATMkRlkx2fhFuYrTHDAidq2WT7BpG
8wo4/BwDD8FB7PTgHJeIhMgrAb7xyp2M2yT4ANPnueP/ehBcDvzMKppnIlN+dulw
2MNXx/o7G+j/lKkFEKn6NNp8eCUkG3/hbbTG8fMuKuS+wDqIm7n0keapsADvhUWv
AH4WKBO9/xUblha0LIkSjTbGw6vUtl3Y6X8Nk2yt6A9u3I3SQ3QdDmDyGmRSLkdU
ZD+CV5YQ/vWx5wR6BIsE7jHoS9Ox+d/44tJLpP5TdO1j6KuEykIMor0TPLPoQMpN
Lt9bCP/3HpnC5+nDoici9+0FWIBl2svelIQEK8ukfLreUwoMqoevzffGrlvwua9E
U8rA4HyxonVDXTh3qy+RBn8CaxyI9pxRDPvd2t9NkP+NKDV07g7nRNxDN/wt5gve
RAEGOkCFLeAoe2er4HjDMDd/b5ydNXtBAylIzgVGneur8f8GG2GP4vhsCDHvP+d+
KBjh3XdAYSbOSRJ3K7R/kL5SRUnddolVcx3VBbYcu7TbB+80jXrDJYLIOTKkFM4i
DeBR2mkxDWjPoLrYTBQv97bdumiZA1uHWN6E6CMrDXHmi3bpEScdxcS+Cn53X1XC
ILjkkFXdFbowjcso+B4ttLFoRoxZnKbbB1SqegesIzEMwSH1Ev9rZiMt23BfgIL8
7RJ5v16GFX7LDuRN23nvFxnykzCXXcJYneqf++roFmfuwTidg2RQXwGoQFLLZdQo
BhuGWYjp/I9t2NfdrW/EfW/SK8oF01eXGJzvW000E0SGrqU/1/8qsVP4PFuqTq+V
GIl5qTrtqXzhFL3kLN21oAQoSaXHK24PGLMuGmSIPGEGfFDF9FXrNBEY2OHCNuaD
siFxXfelYVpEhoucavOn5vKvWZ7RahMGnH9SXT446iG2B0trHjR+9oGeFsoVIR/H
zJmpaqM+AxwiNRZ21kwpS1MWqXRQVBE6YVHo1GGkNA5nuZZ7fs2gS1Xqk46iJRu5
SM+vZlw7O5v2WiPcRYK4y21cT6kAiKe3StHEJpdpzCvGS7Ryj5R0ZV6T5vrIQkbd
GoYvcV3N+zp6q4Rvib+DjSulLh3u8sB5A/O7+fcw9PHFppzw74Dyj93KvWfHpLOb
mWD9rPPLlLGTalXc4UmB2YL8F4A9O2Abbj4QqHPzTuRNQfD4jOhfDkT8rKJEbWwB
O23PKOyUHCEMRw8GP3eJCnVKjAVJQGw2/Upw6kyv5P0dqAjlDoRFhNL/YjOJYLwx
PfO7ondAn8mxCgF2QP4CXkwMmPdclyN9TgX9tlvHmChwEn7f7HZ/BdidJr7L3xrl
2g7tnXPrl6YuQznTpSRWMUHJwDSfeAWgTfUqUpsW39Cuv3j99UTiV/zSveSOfVwT
blRHcV8WPVMppM/dPs8Jd32zoEVcwGahl2qQNYDkI82k9Tt937xOoqUaWAyVg6YQ
0KbXYQdKwstmyPk2uubN8m7RzzzmxZRTY6ax84pEZ2Mg7h/Rv3BPIpYrwlUXC3UL
mG5OzQl9ijjpN9+qOJgi3i15O98aJfS1e5ikF5cgihnvZVml7NHXnAXB6ad38zFd
2tDQ8c5ZMVYg5B4DntyZC2eYRLXOlni1YWiVrn/08nWjKuTv7vKKbc/ZxOsjOfBN
+FTLdIh0z29VDQb7eBKVzf1mbA+XyphH+aUhcKAIDxtOs+zTmBrFWbm7kRBWoDrD
UqRc0Is35qI+2qfOE4P/7pT8hzWpWp/q2bh4lqQMBL1Hfi+AWB9xhnGXKM0yrOvP
wfCHlh2aXiwBAtQvM1udx/1XifgKkygQQvyEjAdVEFyxktiGr6m6Kpn83KgpO3l7
pewKAM4zFlQOjhVkAyp6KcGwI+NDbuqpsFeJFE0AhaMkOGkpMBU1438qM8UM4vAH
AFrARTKzbxWZvie8MpXb+pZ9QtQxvvkdXcVqiNqhnNuZkojcDt9Rlog/a5wNx1KU
R7476OPjaiVb98Kjpi6sfiJBxJMKLFm4VycCQIHKL4I4YYrfdUnWk90/6veN8dQO
MmJsI6/7lp1MRazIgvbPGhS6YNDmnLlq1MX/HKPqTk0SfQEYs9lMt7tNG4gqjT6K
fA1Yj9EyrD+2Z3/PtyF7/AxAuPPdNCjQ9cRCFgHRuMpFStvFiQQoFIQCUvUZmZr1
6CC3SdxsP/KynBOdIL5kYeSmsmSpFKWDa1Z818dwtRo3zd4k6RhVv/Fqil3JgklS
wuaw9zh5pWERaGq/t+4tddBbH0s+KfwDIcS4Pjx3hgiOp12ZksoeqBMsLKu0XgC1
lOz5RCVIurDvXuSaYG+Y2VAznquZnsaoyPiEguJNXPpo3iLJcC/XqKgBowC4t42C
pocETk2SoEpC52P1D5zBDcGia7Owes8Df/G/NCIeBPvfK6aaWhM5KQR58NwBz0kz
AFNWacM3QWrJak2LWqMhG3fqDQXJWRY07CQlucmfQM7crz4gSMS4eNscXIvq9RQu
uGg7Y3Q4x5NhuPa120z6eyq/GzAIVbPIhmSrzfZnyJHTuXJCKc+F9grHKI0DkDG1
lzENrxS2Nyd3Z8OSBGzhJhHKjwCu5w2U/MuRFa6HYkGt2aGLzY5j1ZRgyp+3vjsF
m2wDgDijF47emQnTF7Bk5sUdVxS0RDk8yytsK6KZF2T7Q4R5YFulaCbUiIASHql0
Yal/kebLD7cCiDbr6WQcR39pB4nRLo4n2MqgWnbOaDdXEXKXzwAyUMAtFzr7Lvki
AKcS/nmW14m82QFZ/o31VZUkC5BTgUuKJPwejqU38teDvvfOFh4ga9cW6/FRPlrN
9BN2aqFBl/Y++5rQJQaZuZEFs94gVf8X19chKjIYxWB+lEArHkBxnUAmHrlajOeL
8Wpd2CMAvbWl2kIjrYKlmO2toHUlMVxeI8ojFDXRizJOxFU5BS4qs3bYgSmNh8Om
GQwvbszbUCpzKayIKQJ83R6oQwMO2YodfvK6j26qfshxtHWLFEbzagJwwKDzMa6e
vIAnNy4at/WNbIR5X7buYkTpcocXGEgXatFRDNO++Kzwna9+nUvw+h4UiT9vTEPH
UI2YWt1kEurTxiQxQxDp5u6aFh1W2zHy9ohicfVTxw4IeQuYAWOMvUj3B6kAlhjj
o4wTgj5Hpyp+82nc3sCohx6yKRU5RBChchLgx+d1ngfJUS8lIk8fF5NI3eKeGDjP
9AvdPEk56fC4uub4ZqqOETtLlRFWVDjXo49Z0YScgOjgDvX4/DF+zc8TPL69sr7L
kOUip9dw7SxgwWcOkIuJfrYtZpvIq5CtkIxp0MZuh0g/vPRhVYytIcwKP3o51XxR
ogaWJ82vd4Us+V1KcvRtBShg+v3QzNWfXxnbdS1nHYwW7DzvDYJgiWq5RzXbVsdi
KeStuFcNHxObDqeqYSwsoimdR7CKXmP207XDvOCTTCoZITs3ITM+4JML18R0aDTP
JseIhRiq7EI8u3nCyZyl70vxMKRc+GPySoVFhLrVibIemduFGBpLHwxgHP1OVSMD
xhWwK1QKkb02EsbdPvdcFkdUnfMnnblWwi3JmwrailxuiogyCOXVmoq+yvjr2CYC
apqETu1S9YiFYrAQumG6Dg8Z3lCWj/3S9eg77QSvCbPiqh7BhPmTuH5j6kVZYwhN
0TDGuYrH1Sa82OuNvF1CQop/44gTiK4VEp+78cEHT3VFKoP2ASWpM9yHoeDI4IIs
DD6tox51jrXjN2tHWUOUst489vADaEjOeL4NtKfaefKiAwcT0x6csYYBQhA7ENAu
MABrK+KlhHCqOiuY5a2+brtlsMMjBQ8EWdtxFTKRpTyj6Iy2Vr6+17d2ZjZ2Zk2Z
v0MNybpRDV1gXaGUDNMqrCRm4MOQSSfxylqS5sftUuudb54RvzJWixqML6HTkxnr
i/MM4uEALb3GuNestR3xiIkqX4gSJNfuaTRPtrDDca0bYz7k61y5B1DA2ZTwAr+0
eBlcPiL4YMP+I+5HDzpxLaKtq5szfdT+r8SXOu1pUWCsEPYS3zR/ZLQ93uIgo1kN
3n0Swd7vRITx49p6Xd9oo0J0QNORw3l9zIg7Fxfz1erySFHIASYeMWG6QsBuyqw9
3i+nm9GzeQtKS7LAaU60S3+tfgaJvXXiuV0t3LicK5QSu6MTb3IeAciV79fGqm00
1eiQEzzacXDQwUstPhwshQ//9DGIpKL8U0xWRBlf3UC92VTAihCA4xEOWo86oS0f
iuA5F9oy8uTVgSSGVjyFtI9ebd1rejk+GowEyfBswENumxHaISkmUTwYhVffuSY4
Tje9nA7CIIx9pKPtalC2GLxj8NL62VQzvppw375iunbDWMy8dEW9IjvnWPNoICta
WG4rM33UDmXrLoAu7GPtAn+o6hyJBuTycGl0DSKiYsXebc2kqZ/Vcr0q7p/QvGXB
9OvCr/PK+g8sEA6zmPYCgXsXqa3yVNFkYlJIegmq8xtS7bgW9qcb9UXzTYXX/RmE
Du6NWqLHHEcxc4RAoerph/R+6GsOdqTZUOw3VPbDULY3GKkJtaxFFlCnJj6aZ2fn
WIArA7eICKuR++u0eCqEt3Ed72TSgRoxBWR70kE34lMhLUP7DSwKiC5uUMNSoWsY
irg5Ee5UEuJPM4TD6FUOHLQbss9KEJBJ3YFJkkYNfUSyMvNvHdQnyScsBPojAYvf
tWa/YRpv5wlBeE/Wg4UgovFVgU2FGgYs4KCUJNva6dQuszPLqTI8BjE+IQYsuoA/
wU86ZY55qgVlIaW3bokF1y3G8jbDFBIM+O65jmgemixIwAj5OeaKxA2POZMAGxDT
yo0JG1r2BMTaBO5Vn15xKhXhWVk+YHggWTd97LuBuIN8VkBWItgupn+04Q+E9b5b
UmCVEiIgml4cUlcdqO0QpioxRT938AnXEgklCmz3fppSNJ+d9XrV2+nICT4Q5UUw
PxE2TcbSdAuF3lB8kyebkz0ivuUMn0ywElt33NI5QDdmp/adDZtVrr45Hisaksut
aGdeU/jNluVWhtsYxliK29Rz/2LeUCIPrdzTMRCBP5G3HQVFM7Yf6YzrRSiTUZjb
9KoVmi16TEKsrLMrZn18x19hazWuisDOJfjE9mBHBml8ufnAfgE4E0BzuawucnX9
yf0RnyD7d4kTjkgjSwa5L0jcZ6bXn+jwLOluHATNRU+jjoXBRVh8z/zFZDFazaKA
I15Fk5MHvK70rny8iwdzlWGKfybNN27Ub0xLQ/iXENqS64RYTKEycaMXvyu/1AD/
tfh37xnFTpZo22D5TUWBcIZxDT8zQ8fp4g62s699bWOTmvbyFm6/h7PAsDZl4vrA
SdOrbENWS1yRuUxhc2J4aAOxhMc3nV/YTYNllT+9J5nFDM89IqQBqywnYqDVrTPT
+04u9hs5eUSktGcuCWKXw9ZP1FLnCOgFjBuDRG5x8zcfvWbh9TdP9jg1cUoebtQj
uyoFs4SNPvidUVSaTSh1ptgRmQCkYq2sCQKy1USZsBTxgx+CSpUFg0TBNg6xD53e
DNWssgBS4VD0pplyws3nzQT0+kXKBMeZKVn0mS6PJqYj11v0UQeOhELyeJZbP0AN
zEZFcBIdancpEfQY7dc+Xa3btYdhqxXMQc+8NyHEwQEzOq29Q6Dfv/mdJfeUqDU0
FwniMP/MEVr2peXpL2Wn15fhxufv1ERoLSt3Iwp0qoIAqz27qbRCUHDbxWbd3hus
A1KqsdpVWZ7Q2FSAjqFYkmjzuxULzLTgB6S5mm/CLefEPiMyNSkbrgkwtT/crWJM
OORY/Ln3eD4mLix3lSm2Bj59XMTGRpHBJ9MIGOYdOz0hzh/jBCfe5ljT1YY1E8an
MSsCozI0CIQHG7g5IqiatDGFMBnWKk6iqVReViaQeGASVdMUpn9vsUeFoyk3Ip8p
F/8ImmR+SGyXGFyZVA5nkFkQPUjamYUHJ9MMk15Wq/syTEEg/BATf3SZYWoBe2ww
iEZ1bW4+pr6ZTxgKsR5oyyO5pf4qr0FSEDPVWBmcBwbzAiyDCrVZeWEycZXcxwtd
w+mm61UBFdpp4e37lN/5aTo5MXbexborpCUyfXO4lRU/GNit1lEgPw4/oxACEj3D
tCywsz3S67F5tw477U53BASD5BWNOA1AI2E3oWoxgQranjz2KRpcAAtcoEu7OKMH
aFENHk87k4drKYclBVf811exVAU17AXk1C42ywwJmLSfcpB/RjK8C9u1pCpyyOVs
gHDqr/w/VghZu/kymw82mZiJkLcLgW+5OcRBkdAXl6PXGEzDuW7NHMwK/CZAVdiC
PspkXq0zs4XY0vYQaA4VzFDlZElBrNJIDeANXNVOkbFqeER+1Lt5sD5Zwd9f4TCJ
jRg6LH/8kcUG0UU5iLLMtng6wTef8S2YtaiOtBjI/pHA94y682u4N0NzZNSXZjHi
kTyGJ8t0aKDTzAkwq+TE6xAxK73lxtmmRa0Xi9kPqMrZ9RFvBw0CwOYiULw0Uk2N
G4Y6CcI/u/UJtBfw4Dc2MaY2gZL0BKIQCGHydU5tcryGdkT6AmK34HowTihNVV67
+83cVmm0iU3HCkCBaA2gn0sT4woXS29lIyeCj6BU4Fe8N2xQkPmAcBVhonYhJpOy
OpwXQ8dF8tZ+/FlrE+Hb3AHKbn060cXK5mTRrG1a99us2HUoN7fr1I44iF0dG7EJ
RJ95l/Mpn3IdiEXqDYiyadOLNK6MKZZ+DnIcxCHth1GRnatw0Owal5TCHTsCcLgg
Xf6zZ+wmGqfWuWqmjmWGaujFoI7cGHH+OZkiMzXPA0bm65n2yKvr3+t3m0Wi0Q7Q
5p+AEHFdt+2rUsRpoDG7T0brRKhnTCoypW3SA2UufovfV9GynVQ79qQ5Q1LNUhW0
tReQT7aEzKXV8SvQ1mqMwFshgYaGOyICiXvOLnaEvtY3PMl8g/X4Lex6n+2DSwGd
IIJEswTR5RVz/r7ImJtotx2vYFqThgbGlrSuy+gDZ//sNgiqOjWZOLr9QvqXkaTE
2+AHX+HPe9mkCFyd1YyGYXf6TOSfTsb61X6h0FdfECi+eZy1s/ql2kuTa6jDJO8x
jCUZ07fHdujl4HjZBMRq/R4OTgNXNYAmN15Dz0REMfAEXMoMndpj9u1t+XbvUu0J
SxUYCXU1WJnAkcK2KET7ND4IEdN5M5lI4184pgKhs4j+CUawLIZSiUTIevQq7Cvx
P6nzql0WxitxxvryyMSRHFs7XplKHdGI1Jsa66HsBjXAQ3ZBajRF5LibYferfte/
+9orWykLpcOkf7O1pAXgQOtzHZGzeKQa4AMBQLy2CgStx5iWhzho8abRHMbpVzC1
8VziuIPSB6kg00wmMxzbXSZOIlbqarvCymCJQHP52kiO68VnuQ+VZcy6p49BTJCy
H/uwaMwbZl8h6wq9bK9y39VqymC354s5oo3WqfCEpSND9Ci4l9daS75AcaxsLCTj
XsFRfgbykQAjthuolPBoiiPR+B9Htrm6O9wL28ewbxvpUSVa0Veho1tAZ74qCfwI
lED0RCuJsZodyxPuRfYrx5vDKBnLxoMAL0TLiOkt0uIVgO63Mtz1uH0ZXwy2OM+6
yrP9w3LVWaVVsmrin3K4kpnYaOK1JLxIhB9CNGFuldZ5U3QM4xXPMpi7PLlt3Bva
Y3ozsmNwzgvW98cEkseNg5DZEvOdlb6CB503DcDcxKfqCMrXpdqrz66WynGIi5BH
DYzpRq5GvNaUAGYgu/3PN/S8hY1jA0K9Z0ZWE366TO/lCGKRP64yldn1THd/3Fci
0asf7oQZps2rtEmZ4hxvj6/qQ8ulGzMNZmeS2cEqstMtJdAtsUG41Y6Tu3BLCXGG
+CA0VQgHzJdrPND0bqxHaTQt2rPk4TycqRaM2xY+FeSD3AM3rwGnIuNsxz7NdKoL
JCWCms94HxVGF9iPIRIFbpD+CABOXTZanM+8n47q4C/HcIZFD2Gmvi+FoB4hehAQ
fSwKjTrLWPE9XY3iWnGVYBtMDK04vXr2FjXEM+KO4zTrg6yGCZQzew4+iyDWXcZN
7oWPoLKBXLAh9hibo+z5UH1T9Jd1LcxRlhbIZCB7h8Q8RazFCo2iq8sDMMUc2zyN
vxe8gGf8DASdXcvKn2zU/n8aTz8x4F3OMTuyEqjvKFApVCUQLlPjHx7EA0s7LqGl
kdtrXEiFPuQwc2bv3DQeKoes+m0TshALqaBfpYRvVuH4QqShDdgth7HH0yZN6cJQ
qWirW4vj9W6WxTZ4xxnFocr7/4E6lICffPs0G6m/mJ6lfHsy3EVQHjBn2T1Iy3VV
OUuUsMrO8ZZAbEGLzgaC7zkTDskO3tSHWCKzHuvjVHn26jP2rSgTTx0ElGGgMz5R
TGN62pu1doQHWtxq34tdrl9q3jJobVMXkPL+b3qfBeXGY37R30u/fN0kpM5ODtU2
Q3CokKsY8TvYG0FEhG/0B8wIHukiZk1vhegLYaAQssq1dQxN6mc/i5qYojiDeL3M
hNmJm7gTJRwkZQLuciU3snDiohFZZ/Fb/22oPA7siFo92HttvePLq3yCj8gOeptT
9tiNrSqXa7zzc4LgWMGuxTYpu6BIQ9kCbO0FpF6xzvM6npVEIdLRX59kpM36gV2y
NGY/2lKF+k76laIedxBJAn5vExwf1SKukqNtSuXpLsitoCRk5pMi0gF70MXUF+S7
ApBZM0HLXn6TX6oO/1qYeUNFziMl2YvEJtqHVBkdOOBipLNOXxsUKV43TKrJQaCJ
ilvVGjjH1XFaP5NudfQyFccFosmPP45pWM+5umGAQst4yuy+HUPNkBMPz5ku/Np4
1qP0QL/GHhu/7vJfHrAomFNQxjqxWTiZAzCXBSoJoZUINw5zGbR0zK5gEJJDtLWo
ySEcGKg/TB10gA3z2ZDf3S+tjUxHbzpSl2UVyfgKmeI7X7eJ7pXgCElOjdQmYIbS
Z5Bgi4GWqVirOVnIC3q3KBSHSk2tS0aVMA16AkOuo2T1QuAB0GrImnbZevBZa7Tp
WPCPpRIraCCsEG7ZBdKr2ijaUhA24qSJ58/9Ndi0qKZynq8sK1xvNRrBLlRbvJvg
PeB/nNQIk6RJCmXxyoQ2+rnul5yaLH7YvT9TkS3j6NLYSjBVPGHWEL7/V0rJxT69
7vlyG2lVUe4BFy0jgAvv1a4AEkqEUZlivt0PiIDVGGOV1ictA2EkUJb5Rux8MKfo
MbSGd5sI2G59pMxVZBBVhnXf8eVqHQCJ16heTqoRbzrL5UMbLCLsGsiarfd7kG7g
xZu70c/92MHba3sDTHdbDxJC4C+nXXxFGjFdIQRrCHox4QiXqp7t7Y4jhQK5yQm7
nlfratwid0igCvOQHqKqscG7n1wP7uTP4nUeTshwgfWnr3Qkdek0czBlMjQwbjr+
VcXlxWjFWKBml8Ayx1inHH86mU54NBI2YTE7stVIiobZqM2zUOq2qR2d1vofNrW0
Kq1J9AVETErYTxGv2xbn/QZ+A4n3tRfb0Lvn82GT++nueRN3onZNFKxhPfw3TEQp
lxMxgzW//iaw56yX2FA74hA0VP5BGqXdwh5dSSMBNdSD4UOlKWVBE9wxBMp9mg7c
yF7mSa+zICHLXz+NjDCXgzB7/ZZ/j0wcGcs3M31MecZih6+pq/1/rl0weALnfCQl
VfqcjfJ4cpWWxZ5FuIypfDJKfbedK7pFmbyBKnQsO/DuuF4eSjEqVU4QarPZCAbF
b/dXBA7/za9dD3uwjKrKR/X5VS0SAEx6/Glu2+YK9SBAE9gedXLjCvKMuYxxHlVV
jAfEQYprncqNOpZgJ3ITIXvTIFq/QMATo3DwzPTP6QAaF7vz63+QbyfhNY8P7tqD
zg5VwVr+BrM8/PjHoLoDjfVwqzCxufvSHZB/QUqCsZ635eDDqpR+Q57mrkN54ycm
uIqv5BXkEK/f7ui7dOHhhvEJyrjVcjiq4GzVgZDcCZqtVcZjrF0B265SEYCVvRA2
Q5Im21X0nCzvi95InnjJEiTzXI5D/mL/8wWSfcxdh8ZiJKzk1q7jdZJYClfkG3Ls
bcYRb2Nqq/svN9e/Gl/CnpbjtMJGSz+ncBikkdAT4Yrg7WaviogRJaehpANljUGT
Cs9u1ZiNvueP5QVJDfPyhs68ma3zUpUS0zjwgJvIhAaOw3I4GBO4INMbIFRtlebR
5he/A3Yq2IcZjDFoXt/2eCFsl83sfhan4FGwyg4zIfymbUa9AAjZc4EOqBxIIRnh
ErV+y5p1Cqvd4mEKUsNLouvsdB23tmogbwEJZvFoWSeW6X1lUudv/S1c45/cpGxj
hKW6pSEPgJgtmsd4YzIqFCepHmvMHsOKZPEANw8xXsE1A7Q3+7ZTkHRs/AnR8tFK
QQr982ATw4UDLx+Z89xkA7agfNHU38gLijKmOmldH7nSdHCodOzrNF/3ekAHQMVS
BXfV8DIrNvvGV83fGlyYAE/Ej0Xvh8+rzVVlfozIDiw4kczxh9ccrjTkaRbFHl1t
qgwjPLlriRHmeFTRkSC/MfIJx9zSqZ/rW6O98Ol4WeqiPL5NXOju2otBa3jOiIPe
2VpYPXaaq/KtytyOju7lzo+mGUj+b/pGbCd7IECdNCIR/6XUo7Um1tkGbZRrBw+a
ccy1R5VfT1wC/v8j8o1eWF/k3ihcDhJW+77/fgnUzRQxGl0siQQ/71u2gQg0LNAO
YYkWP2q8MHQWKToi/W1W/Yq0JLp/usK1UFgBA63exT/TKY8Wy3YDXhGNwBgiNU/c
eRpCl17K8MzKqeTWhgjgkEaCMM0vHAjMJcZmoytA7KstP8ZRxe511Zcto+KR4Sio
ANjKFjzqp/CAf9gy9Df7/+/noVwRWwCLOK+A7W4+dgMW1PiW8NDj2iCFbItrHXmR
QmVk+GAALJlQ1POx37EmCUvPZFVn+e39uNNXjrEH6+KC93Y+8V7CWT0gQYZi049n
05OW5MEWnmUgkzbdSH8ql0on+mFLExmDns3b6ey5wu1bMu4pPbXd51m31rBUT81+
i4DOkgoozZUS/UfG8ETMF2ALkBOT+xcO4n323fOdzwyKkG665E9y+qrbG+RV3+yn
HzReZhL12hcYNcPTMOsaYFgOwfj6yD3Oa5JEePQVZ9MtO/HziyPvUFrs51/6k/OZ
p8KSFLfsfFnGqaueciQ3QmNTNt4FTbyLmcm254Qcx/hn5dgPsKhffa7sU9BT2XnD
NRLQ1wEacOHdv9BLxYly76fAdnwksGKxFT9vI3Twa0mNmnRLPfxyJtVr4NSIihh9
l8lKAudCXG6v+o/E8gQvaGWJmWGhPnzCUjYPl7AIQaEcYlhDHQOx24dlyiEJNNNe
vQxdbiMo3cn5u4AkaCBf4q0Ca1Feq8AOqYH1SSJKXpMJyTcTJTdKUmc3GUphWmMk
i+BBbdZQluJJ/HqT0weXDiHtlLtJbOnu57RUgjwFIh9lU3jTIQJB0u7dDbQgiNfJ
oqddar9bWDXWikBIIXd3nEfqxhDdOd6kZOwatx8XuZG3bhT+uDVUPbF7iAY/aE35
2/ndmYzi+sZNRN4rf1JKs35lQSlG0q/BrD3mKOZ8oYjScmQlmDFwyGzEntT569ur
5sWK79/yqdN98x+YdnaVKlv+0XZC9K9JATO/RPmp4YLbIdNGE6o2MwVtktUleUGU
AtunaoxR4aE9hVZgspQePSy+N6bjnJvBkFz1hw6e4Bioisa8nrZbucSGyirAhMZf
19iA/xgEsvgq1UgFyuq6cCvJFM5ba6KCFVn4YJIofXqn6BRRDfkfNQUC7JI851xx
6F9TyASpz2NEuagqI5wDwrMePlQuX6ePR8K3AyEgvdxfc2RCiiMO3Jyy010an9oi
+PyM0mKrpb5nXevlDa3rSXViYhxXOjwZunpJTsppAlwg+XRXSzXjRasp9588xT15
0BrREKypoRL+2IdhYATjOSSZEG25Hjbk4eOiGRRPalRC5MSMSHXtGLPrekK/xNr5
uKRyduoqFhLHMtHie+UmkUGoLL88/GnRWqOYjSXxqgWlkWj1BjvJmu3Fg+vwoRFT
gXXDxTx4SH8TzSQd5gGYnHl2b0/72yXKT/WQ4GlHWyrIFNlj3rXV6zfsrl/jrMwi
KynFyil0hGBYUiZt8tJSM4X2it94TzZjCz6ZqmRHL9CrhslidLwKktZ4V4mKq2uR
XQP3PRTpjajD8fL8+q3MiORcA3jGR3YoIFTvu7l3Jg7NhliXQikAvjqr+8mZceXs
O+ubM1qCcXr459dKsrgpQuSd5q6YVWJTwCjetbSFEC4a0VSiDLlM7xyaZ0wLvgET
Airdf9Bww8HV/1GY5bRkIhUfjbSU7nfW1hVSB6Eh6DHdfm5g2HfSnaftVHcjpM8G
y/MndEqiBipGYhTik0pAhIOirmld5SSIW/6UxOuBZy8k3xuaWOm0F7w8WQkdMn0p
RRqu7cEtvrwsfd3E4McppkmWfwDVaKmUT9iFUeShEkSEa1WZX9XHmWCheGWhFyIE
3mFIFgQD9h1ECwBJ+b7R0fgDq/+mz+VCoPNuLX2rYvBYNCXN9My61uEzOlwVHozG
P4YqJxlXernnc9ZhGxlR6elRJOc6U/oU4xFXVnyzw8yS5eD34NjT0FeJgyCxolDV
aLQ/kN8lrvkyp0oXvCUI9g+Kpqaia60apL5Kk5FUNgeFpGpPF0uHyMbEPyl10EhY
GF7f523O20WqbaxA1Z7r/hs7hQK/rnzlZH+ghSTt3fphLJRzoUZ54pYDCKf5vthb
QgIpHa4/Xv2OBcBMyMph3NHhrKCc9D2YQ6yqYasw5lGKmKzgiH3/iSPkskS9SSe7
tlxHMY23T3sgVtMB4pQ9DWhN3u/4TG8zBp4p9QpJelVsyyev2KGS1oYrHsqTa1l6
6Qn2ioaPJy2sj0lSIom5QN3fxPfcYPGokvWwK8DQxKCsGDYuEtoPy8Y7sFaABzVv
bn7uKHtdfdIMslxt7K/zruOLIfHXtHMe1gEs9sqbIrUdquc1remaDN7ybjnaPlUq
+TMmcdSYfeUnd1d7Zh08ZmhKM8HQD5rnIClGLJ7KLF9ENMSgRTB+dJNm6GTAX0G5
LnrLzZ+XiYHMopWASrLSf/678ipZ/ciQ95268ao7s5RN4IuMLd71oEr7Df5IaW6U
b32BNGNrJs8Xrrhq1+cDWkxz2Tj2XraYx+3LBpuoJUd+dGWq3ussy5bWrq01Iaku
HmJ4yx5LvwLyADhGlQq/8ICE5kLQHtzPSps14sYHiKmkp66US8For4rgfzCWD2AI
GbulKYOkqBmp3oqCFRMXEJ1dwD2gHxGl+cZXAvMhVsHceEQWgkw6v+o3BV0DCJIT
1J2R2T7E9K4oLNTSoNQp4D9btxX7mbuiMzfY+PnfT520hvdpOLH0K6k9thpCY4oW
gDfe2w5oUhN3fuFnn4/XKosyyeYnnZR2aXNQgt+XMRXXIeHTb22vOaSq/pRfBevL
l2zew1JzA01CxffL3xRvbiHLl3yrXz9gLKy2BYBmq6laxjzxKig0tydJWpElIL79
3DdFszk200/kBa8r/cpt0iMhkWHGvjWg28TJulSJgcMXLZA+j6o53s6wp9dpuq1y
ZsdQ7nJa++wvnpQMtit3jOVCRy5fcqRS5ko4j6G3lNG7+yO0ijMZUTbLoFSMABh+
+bbTZQWh4xBEH4DmQ9+uhHpq8EfBd2ymJniGcKtD/W8SbYRmADBst16Fh431kUe/
dP8cKk3KfziZbE1wtQf+YH6ehDtyWZKzeQeHo5oQVhx+KdhbN15vPaNnYbhu4fiW
77FJnpX3phi7PSPsBPIuI9KpOze4p4b7+0oUcUAsvh7Yp+QAQlJBRt+SHn1r/aLU
NYVbDA1hF22Hmp6tN99AKKgQe5gMtVWcp4uSY7EPBuN7Z2nZZKPINU5M+gONIK9f
BVuUuXeh98qI1dlB5caCOd3Egm3dzEG9jbI9Jk6eVtgDhQHh9ZWbeJvW+m2kCiG0
pDgd3nP3N+mOY/QXjA4GVoACIbRikWHo/ViasjagQ4O30MwHjrc/tWdHWgOY/XNt
1kFes8GZtrsEcy9C+CVWpLBXboUfax/S3j4HXerytCCm8P0run7hYcr6NPcM4BPY
9/W7lzXDmmSTx/9YnvifszofWLZH3pCGNL0yz9WSt4d8wkXZJ6Bb5JpESCLfP5Qg
H1dfRthVeSCW5HlSRRNeZ7h0oZRRlb8aDGRypHXJDeuw8UrXoKZl83OIQ9wIHzII
8v8AkJSDbWfYk6RMW5Tu+fkpemJa03Tym7Nzkl+TYSEnKHEJZFVaXmwMeR4mF9sp
siTL7EzQvMtqBwqFCEWIweD6Vkf8UE+8ZnaDvC08LTG2daDFqQEDXDp90lsQpPNO
ECELZYPulG/eMqgx4fw0u1oC5nbCv5ju6E4gn34p7VYd/IwQfL6hgduQQRHCfSkE
qg2iDGGPJ2cqq7+Li5JeX6yEnE+EmHIc7a9L/KtjHD2jrz+wn4zrYkyCjJeaLN+M
3B5CdpcuWcTdL39cqb6n8LD7jKkXGUbtFY//R9/3zBVPu96QuUBOGaKNUBs7SdVX
kyg9yGc0RpzS75fNBQlWudgkko3SiyXqBFX4jmgft3HbIvU2rSknBiV+SEV5sZ9q
AoVHkeI79iKAw7tql0dvm24IEywW3vI3qBmk8c1yFQ6zLCNlS7+GDTs9ySleXzD2
tRaRI7s49aoK4h4shG2cGMAA6Hcgl8LD3Dse0f1JmxAmTLLs+qMa6P5Acbpx6amv
I1+5e01HomX42bpCCx8pnfX2Uok9e/LywPjoaAauPpTpW5Qo0LgDALXMf81Cd1yN
pPCHOEACNtZM76oVe7Ib1ibAWlG2BjNcC2LZFve05P53UAnTdv7l3dC5eQ0DZdCh
fsCCtbtOFIRxtQPQ8d2wYzdgHzkOrFyYtocNuVea2ksXbOfZEvVLSSQf2Nzx6YBd
gzjFfp5vDEPNHB+gvfnLpIa4UV7Xbb6nUIdt29NyOWuEkIFv8ANBNBFnwrqho/W5
Q3Lg3hwangyslro4VCVVrbRrMFP63ftDaRgQBfocTjCBJq/I7ZpnkNwTh8N3xqSN
OYQFMi1VU1vWw9w7X5HFAl05ULBsvwsdPLN+3FPGvmT9ID++ay62k9y9vytzLYSu
mP5AYWadrBsFTKHHiXEbUrsKN/6t9c6jXeoyrDf+udr3JenrMTWFz8Ot4jNKVYfz
enAdfLkG7H32f6IsS1vKn9XbKfTAcVC6GJQHdfHoaYsAjzTCyaYdLvBVaR9j3VTq
ouOfi8IAXk3wXM1sEwHGb+4wLDvJHDY63kdphZAp1gLNNpAlOIToO4wkIBe4S3jc
5bTEfVo4vA9o4Ub766BOV4HMOX01ApBB1gMAXA8fFNvjFgtDCLrD2fej5//rsCe8
eChRkXK05qHwBnu2WCbpNjvbXloQdWWfaX+eMMTK9DviiBfp65XxwHC0gtTedb1e
VwPncerNNgCEICkkH9Ew4sYo7aa0rl9IPoJjJtYiqcTkIQDlMrUgSx/rcHt7kv9J
OrrGcuPpW6TpuyKgujArk8ppYoXO1k+f+5EmI/v6sV/eg0yselkLxqJXo3XcWLqX
k+3TP3X4mXBAnXutpCSwuFI/a/GT/QMsBmCmNH3wsJhz6b7gQq7FnmfDxljKmrEa
Ztx/ec6TJ/4+Ibs11jEPVkhR4kKYo66zHYAz/u5PqHcWR1/jzxmb4n8d1IM4c7X8
mH7ovkijDgrJCFKivxl5/gQ6axv9Vdfak5DNVE4W2hj+KojHDbEAKbZcjRMUOpmI
YZdPaPlCeUIrB7E1t6o7BMh1yCovNMEAubR9xz14Wo4kuIHgndDNd0wyYSt9VG+a
UA1wZq0stpZjn371I8Erye/3rlGZDgPEK4pRtnS+7Gc01VxAZrkhEVF1xS9PXZ87
OD33156/MEwAxLEQ9JPJt6UCi94nHy4nAVCPC2oawNpETcLd8WLbmeQfaN8VWkfF
nef9gO21Lg0V923LFVswXD8XTF1laEPTSPe0nQ3jeq7L6YegoctQE5BNDhCWxDIo
C5pKY5vEdIImYx6f0H1BNnBPG3M74ZkQYfphNzqRKk/+eJvLBF055HvROR4qJCpL
cYYle+BnV2sIOQt5ekLMTlXMOA0uF5xq3Mb/ILGGg/nNEPaVqsoEFvXeOx6HUtaH
DijTFrsAOVG60F9dlX5DNz6YxnoufxEFNGtZDfKddI7HhWV9zo89IKAHYL9KVIMy
6IPAqC0V9Gm/ku/NYSX1/ftYG+xGMmwOd+NM60N5Fwg+uwqsD55yDnvkXeKmi8Hc
ofDU/106HQaP8rSkvWFymEbzw17hgEbYp7oxzRqvzZCCegsU3qKKFCQuPEzE266W
O6+E7tHvHwhxrGomBcLmYL0p/IrJaW1fE41mbbP2f3+rTsd+NjmHLHtr1s2jiQMc
ruJLq8TYuYrbKEnYhRr0I0WWsxrGlJGZtcp7VW1C5/BMaTk49gfud8gvDaTCwsdy
ngbDaxpRMvAk8+yEi6XCufd3CgJg8NEzqZJzrQcZTGO/meMn4hdk3eRIfwEpPsJi
liBpVfHeoUJ2nJQymaRZeVTHfbtQ+J0EXZKy/rivZGgbnUJ5YKjDOwVpMIXW4oCj
7Bcs0yGrOa01Z13ered2b9ij2+Uk+hZhO6JRxnM3ywnFYEtkyS9GgdTEqFs6IwtA
ld7Mn5yXTw2FvY/3pnoR6M4vy3zwyQWhtM0TeonVQyd1fhGboJ5vm4hKx6Ccuhzw
JI/EQizXiNZiXBCHuPnBVWF7FPKoQGHRcCxuXZyE0cNcBkMgzgx+qN4StoFrrEqH
eTqIZkuu3cIa+va+6Quy/FiKO8raM9ChXN4d80q9NaAHvHM74n3JHxd5F2uBJvzE
4YZQf4yl7A6stRM2/szpKGivFU9EHx2MmzooJnNGWuq0TDHZvD32FZj5r/NN/YnE
fRUuGXm5m0rvMGJ7OgPwj133rSjXDKsJkBaNE6S2yjrwI02goQrs3iJuuvyBftym
J/56N0xUgCy8fNXAtwAf8E+Jq8tm0kVuIjlwVSncGXI73ozvb2UqQd9n2twfX5Q9
DfJuM/wyjS7BsVh3v4sbsI8Tmx7DY9ultigKkgJCGyCBOwm52fps4CD3ukJwx+Bt
NlpK5JKBnp1kpHBAgXpkKiWBoLhrE4mKWF9idDShPbe+vFRRENp4RQlB64fYHOGw
iGSs7WVHKojgoOl4lrh0gTL7hZDv2H0Kup7dg+Cuj2nj2lfobU2TvQhGRDFIqHIN
c9uCwDO5aIBcFBXwJexh31w5HvYmR822ZO87WDWvh8POmXYbhR8cb1wcVpIdSvuC
gPWMn11SPsX6NivbBBinLJs8fZmGFEon+MEuYVJ6LIPXfsyyGdSKckOGnpkuvZVZ
SWSKVnGIBfqR4dmQr5RhC/33H4THcOGhjwgm8ZTj2jygDmgVriMTrgEzglGd8gNR
q7oQ9XE0PG6N+Xu9+d352hcrBZxvO6zY3Y0MgysGLobUjFnNgGupXsF9Y9zYtEQs
lUXtuZmwgnIu4/y2BCns6bYasP488YObu3wetW98PV77G2qxP5KhGvdw3DpuaZZA
oYlYrtlwxSJMZja2PObCVrRPCBlmDHfshcHRaNLBvkG5g99Ae9sj756rP4pMtBiB
2VOhXICLqg5xEVP1JEZv0UQUVbXnMrp/9r9TWV3JUaFpjrZ8Pi942VZBrFkEMMEm
8/be778InuIwF9gRxOkEzmQHjsdjmz1alFOTjb8eAYEJ3wBDXLdzMup61WufN4YL
jz1g5iqo7pPfTGQHikWhtMlpZdp5eEC/23YQ9w9UW+/MEOyFjqHe9IPaxvT8H+A7
etD8cvSAM4iBxWPAvvYQ6vAmRaIGwmmue8tDmQ6UV5W58LDhUtkp3VimvcEtYLa8
uE2GxBzJ3CaK8ftQDrDiZuWo7R4TTtsFq9VynT6cVBEgKPGxH00uFlxxiTKxpI1C
LWAOma68Io+XsXfJMtNSfAmN1ked4t6qWMuc2V59dNATC4/fkeRUNg8wqJ1eOrAy
Kt2t1cNud0szHQOVkr3ce40Kg3wqEcW/Yq/pudH2dIwCCiCobvTBc44EehxIu5cZ
S+ZTYwhmNfXi5m752Fgw96MaTxdZ20PIU4nblndFtPQFWB+WCHqSsrwNIg7xUTpS
Euj9D9DqePgje52NSgKEeTGDuDfyhmF1jMgs11RozQfraG9ULtT6TktmUue0oBmD
TubTQrGBC7DMM5Q5R5K36DELTsq2oQHCIeyIuLMzbmgBQrRSCN0embDJEjOTAycO
koVsIeldXuu/iOPjB0w4ccpbOZdO90Nybk3Lp2tTEJpf61XJXXztkAU7b/43JKnb
/1Lbgp643Ke3dWbxfFWFaalII6zbnASCxfJnflHRlALsHaUzDZdGlcoFn5hCqJ5g
wGANacT113Uctr+4RgpYTo2zk4KDWkk0JQKxexuuvVQEiKim2qYGS086EUhsUSPM
D0IUmkqPAxLDc8CG7p0+j2kc1/wMlMYspwly6Bbv+BNMY4A2XWrJ9Jwk8nIzU9uM
xvq/SZ/PC2syIREGw6v7UdPrqZnMMLDe7VTaepRllLAwwEjvXCu9hdK6W/m73H78
1QG19lBPgRlhONR680lbctFq8MQrbANfjtkOLKeigD3qJIwIhQJuilwQVOhmik3r
YxUCaXzos86s12tjCySNFqP4AshijeZGjAK9mnTU6GcWCkt3NmksJAdKSh793RUv
hd/jaRAwxCI4A6JoGoCnz+qFBQoI5l2/t+Pps+MG639/vC5x0DF+vsy6cdrx8Kek
/VD4Oe/GmjpH/hyLjRLmgm4KpMkYqqdrFYuahLirIWUqfjBAfiJMpMyuFJ/do2pn
EZpIkRTTphSXwRpmVzugGeA4h2lKNp5/nEQkCwgCcx11N4el1e1diKsEPjy1rtQO
0L+JKQME8vSaLro8MdAgpbEemC9+Ij78V4+I/geKDHwPf2scL/+QPIMO/LgvnAx9
a1GLVGR6L/51lFpoOBr0+Ekfnzvcv+SWY/KlFrN4N+Pg51w7EU7TZ4QgmPRaytVy
5/Yl11uFQoK5fkswmmEs3FMgssQE6StaKUPfm0ZZVRLFleX/+qWIenlSUKrVH0hs
8UNQYFBJIyXK0wwZCPWvEZ7wfa94j7sVU4KUSPC9enux4/gF8zDWsEUBd0Ughv07
kACnssQAJg+045nMOR3JbE7Rp897LaqGQAS6P+JMh9dxEqi870kGwu8hw/ZxU7pY
VigrWNjUBCnoNYhDhswc7jMO/aE+uWJGvIdjdrPdfjFOOQdsaYzCzj6DAGEutxbd
25Uk/J3MgQVzwEm0F1Uzxv9Rxvx7kncf2Mki/wZ7CUAtRD+DBO+KugyMVAiYsACo
W9iA/x08THQ6CdleGbkCT4oFlggtdOv1xOaUb1aRTLzlc+sRJ51gDChWLhOusWAk
XJqSBEwLN3Wg3VOBhXlICEhYFHGBMWhypMmF8bPSqpNmKsipk2EHmerlhQ9e68qb
WQmgY/QG3SqDgqW5NcNB+2Ol0FWzAH8Oupg2FUfEGOmBtfACMcBj7JBMmusDwt4J
o0ZSX8M+xnxaLWddl7q0/ZPb9miY+BNbWBgzjcVf30PBf5r/wFGtncAZ+KN6MHI9
Qd5kc1NKRIuc9dgt2hj+d4UtbR0Uhyb6FsgkApK/IJNkwU99oKZhHMoOnc5msvPm
8x2YCl5Z5BeR8gdfCwKFnhN5VQspxKa8+HSss68RhUddZUctg/YnbNIgVRtFRWrY
fyy73TNYC4sx88/3l6DsfkEcTgiRk3LbOEG8bFWEGPA4YNnYoH0xl9Olrom2aWct
ePI+5WAjkdtevrNxcYUbndFr4Vilj/3V17HC03KcFj8UP8l1clQ5QXcJYCaan27D
7/LEANordM0kSdtSuB/fFuLAepSL6XQa9to7h2OyRLa5yEQVKsIOYvqT5zfdc3Sj
uRVIZAXTSUph9+aCzGBXRTj0vDPy5DYMwlmzVEz6pwGVYyTLPMKpqtLrohuVudDj
k/o0iV44MsIAJwI++7xEpp0O+eqBUUdXIDhYJG9AV0h9f14iZAHozd6cd+Zbbx8I
4rTPxsWJ0I9L5eHiIaJBeAWYxKH0JXBUEVJYCEEHM71XX34Xi7V2ZA/c33RfVQIL
1W7HWx2YLNawybOLXdrWTO+soUNz9HVRDspn7vSrIjxAZ5dZPapJH8W2YavMZ26i
yKZInJ2bQeC/NHGMT/tuToyiJDkKYcgsDtXLJvE40zGI5zcp5u3P/tcQFQZRYGVS
c3TfxCKPCkAy/3e7xWnDbY+wMJIIyIb3Em2HilFkBmO71rw84GYAAxkWqfj7FxPO
C2wzEry+RZfLqfvHJs4R+NOouchBCIm+Fb0RIPyiJJ1huLs01NMaV44Q/TiE8wfW
WYd4Y+Fnuwh7gSshusGACieyG50VJpSQS6pHDtOXf4o7WB11+I2780aBNFIQEcfM
aMH6dF4Jc4Jg47e5FfoSxaucaWD2B1AeBtDATv7wXs9O4DK71p2D9w8HQ6mGRM23
gLUBnbaCCNi8tc77v5fgoo6O2XQpnGM8lXEB+5KlodJ7NewPAT0puSLAt10ytxjW
Qcd1bcwMTH7XHOX9077N3IUX5jh9+2QsF4YRpnGgTKbKbwhu8lEzs5X0R3v36MQq
suoLHyInllSq+27IHti7bd4Ts9/4YGv6TUcn6b5tKaYx5jj0iH3CayoFTSr2lOTr
IgqL05+UKNfnNOvIcJ5CWn/iPkch0wr3jNJFNHHInFb+dy6DHidKK5yRFAO+lwLJ
Otq3u64ys2KDi1p2G02tGzdSIBp7qwcsE0xlMW0z24jL1t72bELsWvHXpUKQwMdx
aO8JOKARNMzoMITeukjWi/Hl7vKde4pWLW/tX49u89Sj7IJE852ouF/mDQrCmWOY
JpNhtf6D2p2yzP413EUFQ8JGjLNmijY0JTXupsqx5wo+/4E1prjXbSiRsP3t8lOE
UgOvJ0LD8xy+fIX4OXUHD5MjZxHuJeDSVI55a5aKiT9JtzmaBKHS6dnfthpDqIt8
Sv0/1pRzgaYCf/0BeTA+64Fg8BKgNfvVUYW0QZ9CUItYb08X9vSAgmqyCcDU8/0i
xdP7ZPRLViSI9wleENIcY3szprM0MOzKh2M1vJFyHGzb4mnV0CGRCs7PYwZlQmWt
Pi/OjaioFbsmZUtupp2TusSL1xiD9rTT7wDaCnkKCl65ERuO/Z9bwcCM/NlcCynp
gLW1+kkY8LZCWFN8vxbJ+GNCTMxeKmi2NSMmQcDJ4r/YssA8mGH+4NxSZ6khJoDJ
iEPND9gIZyKeY2j19dFQlsfNtyzR60dXXRz2HWjwB9/LwvUykqxMxGILHnjv2jSC
+Z7WvB+SW/nBhn6/jLTCWZelCghRu0CfeQcNchRxEa/OYCOuLwJuIIKHKVmOABqb
9/ifJ60aC2BEjZ1FH83iAaEnj+Pf/KSnWtLmpSO2LglbZGpCm2QtPBaxyF90KSYW
5eJTiqzYGAzYc+aKElsFWxUMMsjJhcbmnog6feROGh48ChwniJxqdY+EGsJyXrwm
WEzJLYxcnXr1YSy4Po1mWxSxiyrlD1/ZMYBbiyyoLmds5pFTmo1HFzry8VFp9uuL
WTd09AZvT+zPKrGDR2q87PXyxh+8UrHk91QrKz6U2vqv3bvi3xnl4vRFljZZ9CSb
7JkCgFbOvKHZkX6JW2EwcCXRVh7ErGibeQulURliAW6lGJSD4OZGM/SAqFKg04YE
3nnXkkXGhK8srL4JbAuyWS7zrdV6asq1np6atZ8H+xGqrmcOQECWQzqKkT+x6KWu
eqX6DV6PiBAZ7evzCTGd1uMjhbCGOmn+JPGNQWpFZhNtzFpBjq83GvXTf6lWjORD
obhL24nVCx0E0Obnyyw8q5awwLuIMWAItYpNPOHMqrCV5DIiWVDgitPZ2CB9xWvz
3mRGNsDJ+B5RLE+VpndaAM3SAibayL5eHXDeKfSW8BLzx8ihalzjk//dUYYzt99y
3vDjiCVBxGikB19aUr6+I0NFTuIWhdLlHVxmfLaGks3m9dXw/vL+MSt5cYebH8LB
xIcO0/01b485KYK/nxX2Pzx0bIoSPR+NYuA+FGls3Cz69Rr2r/ldWBdgY+2o0OmQ
U8VIkOBZNlzb8GoaWIj/JsgehPMHXD77LUXULyfu5ERuUjvo9aFofhQ2OwHTEeS/
RKtmMzDeCy4D36Fs6/uck/y4cNNYihm4qmtxy/B6p6Jo0inqFHFjkd7QGdA0ODsv
+4AxYgHYfgqXBoiaP+kai4l+52XPBaW66fmutnoD8o7s7oOtur7Wk/lW/FTmx5ep
g85ujATwy4bR5Qf/4Lr9fRwGV9jWvYKKvnI6rfS5RKbgMxe2eg1H1NSnbGufiHts
J3Jc/xN5bmg/TvUzO7GO7u7jGDiDTBXw9oO3z9p8YKLo6/xes9eRk34zdM+QkJIi
W/cPEkrEWGV9c/q+KwAmRLQO4hB6+mJpgXB3E3HDdtV6K3buLZjBElLauJv08H2l
Z8JQJUAn8eR8SINVstCeao4fo9i1q68Examz2mNNuUvDEA+inESOzXIrkuvucpDs
YTItpjjNPhw5CO1J+j5l3oxCSb5Ta8mjZTKLUU++cmLcQcnyP1cF6jEy/s2hms9O
U4n0ZC3NkDlkQEdul+2rrh3qgTgMErd6QRlsWx4hzX+uRtuRsi3y7kuvILhFAV2q
GG31ofqw+s+ORcHA5iswebhjlaL2mosQ/CkVz04ICfYLsIeRY16MeDZ4Vh6s/oAC
QeLE45hCDbqkzwhF/vFui+aHaOGAd10hdNSrUc8QBCPjrs9EtXbxwngBm54A9P0z
oBCTOsadqcnj8VTGtqDF3i0NlJ0RcftK5ZfMvWdWQI0j1ggAOy51bibfuqdrmopx
hXm5+EM4omaJSGayGQEaaDUTY3QeUob7E1dZdHrKbgt8qg1m0H+4oelufe7mWbha
3+3zPJHYR0nh0p5abcbIjB3xldhEAdCHNG/FajoelXY2cyDSs0HQvJg+y1jPwWCF
EiT2PfntKufbRA1MWnfXn3/RkZvMi5R3q3t8qhluHvuZq9rUG4ln8pNbgCpPR0Te
GntP6U/+voejom6+ED6vgJjkuwhmyNF3HhZErb1hyR3KoXGbe1EM4YxszCfnWft1
35MZnFxz/jcTsNfghFmRvPvgDBEWtf9QHUPK8KZNc+gTBHJUL+LRrpFkJG3JGWZQ
1FwKRm0ChAoscOMP8aYVKgD76ee/xk1df6XqVdvjVx5Jnc3oYowRFMKtbZTQlizR
w/FVbvwnd0X90jc3SRZifMVcff7ZJ3vVt75uuY34QFbwv59nbsMdLbsWFsLTwNdU
e0UkpixRjegMcj8w4Pq/hFdbY0DEc5t7PyeJTu1yMpY+xZV2kzmiktWKr8IfgB5U
cRrZWI9Yr8tgs5kdk6Tb7dOn/40qIsxKlJ09uJ/XSV16fT7FvSGSaI2CJnTMYB0F
CaqDEaU0ZXysAFBeM4sEydiEz+FF0Chk1ZNRdcVCJdqJbYkurtSKTGq+q7L7rzlf
rOBon/QNE7ZHK99MpCVif7xIIo3xFC0fjHol93mFpgIenEI/QmlHED2rc5B0o+GI
HrPXIAorO8s8tqGdiPG60qMyESUgiFl8IDnz4KqtnBF5AQBsf/AwlgN0crQNbsKZ
aZI6ozk8Ax+dEnZ1p00vnTu2KIVALYSF1g3UkkZbjrPFTiXGhCYa9vQ5uwoP1Lfs
CLlsZ38qRksyGjOsNow2kf0PwTwG5li8CXh2YT3RFPo6GdquNKFhWXiggHIIsagW
9sI0bF0V4lrru6BFxPN3Xkmh17a6xYfZqWUTp/CwtUK4SuklQdr3W9TdqqGW6Ahg
YxEEI9aNaSq2jnPKChCj5lFcZ22NFNoy13UGqIjjdv00Kx0VZDOxmXbhBmLvWHHx
MpDKn6KLmwF1TAenbBU0jDYZ+PfwcWZQ2q83kBodSrvbn/VrGzcqcARKo7cMENS8
1Zz4kRKW3jFjzwensSD1q2dQmDsjRWEbq2/YFt1QUB213zpOmhuZa1C5Tz0XHOMA
TbD0qWkZtbZueb6egz4njKW0mCSC8tvmykg/zDltVjrMeUXJGRo6Z1SgciOHEJEn
dn7kadKpDVnyt5/ka+/5p9o6kvfREOxJjfqH4HCUTKK2pLfhmMTF6/PcI0IfRomB
RHp8fnMh2pYrRx0lSQLaQIknzW/aYgwAfbVLeGZCbr3VKb6hq74vjAJwC/Fh+Kls
78WtHHYxPIEOkj1VrHOzRSPmZJ7J6IHL1qCxx0O8UHxIpnAuLMiINZUqeOm9D/vI
LcJd19fNue9vrruqv26NMIhwNUupIumL+reFo7GBAn/onvwbjz0IHVGL895EaoOn
M8GhWOrVasFf/2tfLXjX+ygTeAganbskW+BKjrgLpEG+FkhyHbEK/TAuzBA75EOj
eUw8gWCcMwAzQ6kyJ07OQNLYhq2M4pHO3SkE0Wu9qJ3usbVKP1+bN3K8/DLOkGRu
E5C65e+6G1LyXPSw205wn7GaoskDcAFwBFAOYtGajcNItO+dxylUWNYlDl8G/glw
r3Wf2peTFP8dxrr1OqYE1ena0q+jkiuLOZEkbGZlHgEeAO+PvAzKA++frUzBEkPa
AqFxArsJfiR2F1y2Nq5wXmUBKUjOaYWo+zH5c+442GX937+ET+N2Yalt1g2FfoNt
700hSpYk9qvWNPkMO0PGg/jIZNsr4/38hYYQqw9BOSEZkzw7675AuimwAbwXbUPS
h0cEToyJFqGqJTuEHJuJDBlB//HB4WOsjUAljJKT3cBXuS0gbywNawAkSkI7P0KD
rakcjVN773FLe0b0sBVy6m4C7S+nkM98w4jZp/p3lHzL0Z2G9rLyhHuyPkW5WQDQ
dzLuZPMC2E77+GgpzOUk1KD8gRq+d3USRsU7JOTqye/jHSHIEXKbgtfQGSwSFQo+
dJRgmb1rO6L+wibWDGSrO25s9eS4Ha9cN1BNAL03tUYxIamP2sPgJSwcZl/9LGPo
ywhRgANS/Duamx6hPg0OKbebstImI415/I/J4C9fneiqrE7pcUYSjc8E9Fcgg5wl
2FAx+Iq0xwbl/gdXKOF4R7iZobPupQL7ysjZ+FhlHIGiUYBajPNma7ou1mywDvCf
dtz01nqUPzD7VFFnb1h74Lf8FALW+BFnLBi5LTFAeGBPJigWs2VW3YdxjJL6hvmm
44t5FjyD64YAu5b5wM6b487qsIrzND3XFFhFQ4KUzUPLHknRMF56lFUtbe24KhRc
7UXgfi5Wg808JmnfJc8T7e1iVe316V3IY+Lln6OD28Lu34YgatVwRnjfh5erlcSJ
gKdBdZQbbJqwVzeke+vIG3xC3FdnB8E3XTX+UFz8NaPWT9ckQFPARb88GP5ErkBL
7p7NNNMDdFcDBwdPKQHZCI9nj5U1XpdsJfEwe4jKPYU5Sq0c1m+G3edi+WpupFEd
127Nxqaf8opwmzCHK3lREzvWPhplSLYKicZbs0A20ln+SjygkzHrkt8iMcmodaLX
xTNC3CLQ4geikiAFCe7wmuCUlutffqayuUajoLgfFL8JDsNqfBPAdzF/nWpJponj
gPmcdM2xh4QCGGpiI8Sg4k0LLUbw91WD6FTQYLHrsfw4CDN0ejKVhvO0PVrYsWd+
tT6wWTolY11abzHBGGCJNA9Cc8ANHpq7P97c/fnsZskKxHo0lhDDTq1kagYhZ75/
/CKEcHFt3b8IJO9YqG+flS8NeKQ4XlmVfhDPo6MDHQPmRXrX36SLIryFwj78pP5b
Pr/zRE6nQHTkZ11Qc+/8WyPsE2ugmaz4m8R7X9A0FORs1mt6j+bKIXHx+KQJ5sPC
lXF3sV+lAKWZIWrurqfFz7hTmOs5C4w3Dn+GL26dqQOzLt4gct6LFmts+WXOihYJ
ubLlGxu7gCQ8VrlAEx4jkaxOjPEjgxOlH+uHbazY6siQ+3S5ASdQ013r+Zh3h/WQ
KMza6ldoq0KmZBLFsDn3aPsmwA3TEpmdr1u2yrNTJCYuL3GcWMXxs7u6tcj02GNR
NtMVTzNIlKvcqqO7bTeAwUMzTgw+CBxUCVZUZWL7oga3j0L7SY7q1wjWIR7b4I5X
m1+VxGo4BVN7yQyEl7w/SgoKQKsBLHPmlQGxVhN1tgTQHNDCuZpFf4UFrmNPDRGm
ZvsOK3D02Fs0/n/44riVtZDQlx5Akn+rsFKr6lHfi/BlQtEP/O4cgXD+e+5BhGoW
8Sa7D3ekuT8XkWNZfL5tRBQ+cZFzy/KnDWbL3ftouAcA/Ay6hUGq7oowTxQ0iHdW
KjaJeyxDqoElLV3PqnI3kmnXKKGj0c46Bz74J5hzcfEB6mfg20GwNMzV4MXthtZv
2lNi2j7O/Fbg6EUMquvKrQc02GfKh+DdeVW1r+JMQ72GyjD3TpWAt17S8wQkXlmY
J62fKMNnKVzRcs97QVgdMcH+jDQTEoORD8Nm4ywsm5FRGM9oAqqA2C6nCQRSrQtF
7GmrlvnwHWozMfDbcqwV5KSIaW3dtpEFjfNRgza8PQp34HUdEjxKtebcY5k38+gx
e2y+OxAKU+FR+5S9BZ5PR9hyVxBykqTDxF4e4O19HLihWNLXaDiUGiKeGG7oXra9
9WHm+1U9vbZZpInajTMPDmEBChYcd5dzNpgDderfh2co9ScgL1ltlbQydT3yW4aC
dt1xO/IPEsptB7jY23G3yKiimoFhaqzlplscMuvd0gQzEjuRryuMfWzf/eRWcFhN
9mxRnODQpaw/uGvymN6Kv1CgZPgC624mmzL3UpwPYPE1Odhk+ncf7ZaLVSOGhsWA
KCgnQHWQ+ItL2fGUnCBHvSp6/seRKxO41cEArVMWpE9Vy3h+WD8xnoF4lThfMgCA
toBruYvq29aBR6VoyBql0cNYCiRV9DdBUNZMtOXFhgoNfroCz+hCqKeN8ycSHKiR
glpmjMLLBpIm7duJ+/Yo41VyDFnCMfnOfTDhLqRMUDW2QjdSRyaWO6sewBpsmZ6G
ryVL9J2ju8UmPY1pCV3xbiHwNrWxVfNo6hmFXaPMivGA0tIYIK3Grsh1z7LeEz25
MZCzGNLDep41mRt+uwf5ijAscSH1+3L4xqG/zaBBCQMLjrTTJw3EaTEm5f6OQBKr
e3BN14HvPaXbAcTjSU5zlnNYYHD/RzhZzOJNZHZN5UV5bRg1eoyMthQ9zgNrJV0/
N0uE5IPvsyG5JCYrUbMDVUA8QeOj46AWJPjDxFd+JDajRBBQ/Vths3VhMXfpKrZF
r2nOjvr96ojuxZvQndHD5vIhJkiXhZfAJcYGMe9zDQDfUJCBZD/gU6h8NItIFCge
LNeZZfQ6QFGQpvobzz2YFY2+KURLHUnW3jrz62s1gDv+Mo2yrKrfswhKy4K5KoUq
QIaYsmTfb6SLAyvT3THab0U/ezXU0uW8lIH0TNWinBOq01+m4WBMnGwhJjlhgkno
GZ64UB1dWb8LrxnKCA9rMG0x0gLaKFPR6EkVGbLYa9gAe1A/icgZkg1aGE15zrHi
w0CT5gyU2i9WARbuKxYew7/SXV2IH55JD/Ptr+AkohOU52EZbeS4tEGIYoKSet9H
4tcTZF23CZddwwxcJfwWExdSozY6TQCDNA2xtCskyGm4L84bS1WjyfyWMYFCea9L
H2OEpyhn+OUxxKcZtE8Gm5sSKLPK9QZ9k+SQ+okY98zOFkKLqWwbO4zQwIumB09w
YjrmWVoJmH9vmOFBCYPEMHgXasltHst6da/BaeSc9NNQphX/ZW1yjh8ZNenaCHNl
KYp1X/bAIxUAzJJ5FOUy9hztBfuE5iUnn7D5DiuQGZjTIYXVGTuDwesyUU/yjf9u
QVUN3VZ3NB99Jnrw4A0cJR8QeSfw0TMZWkGmYS9Wdul1dqhpGw4KiOseDyI+hbmt
gZr97IrayQAy+Gz+E9K3OVj/TObOZJvbdGkThNVvFkA4gcMsqWzPz1toLpVe1KA8
pJtXU/Uj/wGwfrmEaz5q/6Eqg6nNAZQQ72ZKPLhnKV0jdzNMOLvBRKW0p3sJmhBG
Zj7PcBMvmcrg8ghIh2IEmIsBOBmSGd05BqGmEmHVfPAhBKIdoAvuJzTqH2gdVnNr
8A0C7QFmfSugT2ZzcOe++72aMrVvMmbkDNqqtPxJJuKfDW7438s0g83En4rFO2P2
FKquvPA1XNpvzoqqc1jMucC5gJAjQOCJ2qWBKuq4r70STJIYvXMGIkTuFGoA3r56
K1TNuyhuJNLTpNcT5VQS3Oy7QUQ8vn3wsYHtpEiXvIb943Htcdr5Klr8qJ+vlz+1
fRxn++sro7folnjghRbLVW/7DlRk753wGud90Plemyi3pSdHVv/hexNniaBi/PqG
SiwkwDUogBlsb57X8rMSEoJ44Tpw+7RBiHt77u3PSyfkNmZUTYjD9UfeogDonE1Q
gcAUkoY45Me8yh1AEjK/FqwKveEZjoiQPxizKhaE+AoelGm/7zzVTstYTYXYujmK
x8BDvcB1oaSdQg1XFIhtNelN2o8LmbS6LkYLGVEh/9bQrj5O5ZCe9AShoVRjVCkg
TJn+POpGCcIXJOmI5hV2Z9icdqfXnRuysI5iwpanmuQ1lqIk975X1NI1WZ+8QZ0h
qSP7yrflXudPLz8XekJ6ANrERwlT8ucoNFCAy18bs33dm2RFlUu1kI/jJKcKRQ7n
RQxDD5uYTNFYXhG8rYxwR5S3zDR05L4Zk1p0qL3JYNEqgL3AG8fvYvZxQuCfeCh/
uWHRPdFa9S22ywyxOiSB0Gzeu4tA+7S+lPnV87WoL2A7zrPpP85whOCUJyCLvbba
Gh6BI8LAPIPru3gr+ho0MCUgJbR6w387+uprlsLQnkpEjXZxwFHt+o8eJdzE5CyD
ux9U6JJjHiZSVCnQszvXjxB5eMwN6Oda1ZGS1LirZ7NyL8P0fmX5LQsoODxQykhy
W65FMCvlD1V9Nvy6S0kWWI8Fn8HSAwK03gBgLBO05eUra6IPkvbaTDmNRE88EYM3
WUY72Q4TZdY5Y99dwLvnTIQwWXof+LjTfBUnfRJtAEkyEnv0B39BCQy8qfMhjMn1
Ydr44wn8dg232tYNMJ9nuDmYw0KciLWwinq4YQdQkJ2pskc64sBnQWfXNMiC+Cc2
QMsQlU00Lp3Z0UBc7IRnKBlOMO65E5ts9lser7pZ4L2WLlewgKepXOcT6x4VS6tl
VVMkuBxm0QptR3d3x5fR14vdQYZVv6Yi8t1gcpBGuOfj2Bf5rhNfcLtrBoSRiTP1
AxckNmCs3kwjFun30XkhqPT4ikoIbNC0Tco2vCT9BBicpIK77apltkjKEKOM2+rl
Et7KCf8xj8vsb3hqm6uSTV7NWSY8DL78RFdLQ9rlVOX1AtO0uoDK7w2jq4ElJhm5
Xlwzr+X7cP6tVpT2YSUyO/XP5ebd/xomRSBuWgEKJZhQgNbjekERvzfJ4kcxz84a
BzrmVN0zyX0ccKBdX4lQ77KdsToQBDpbPjpf92Bup9CD8aq8HFnyQ9zv4yW0/v7G
nsAcF//V8oVVQMLiz6C7idMuiJ1cuvSZKhBJAP6EVzITh0TKpMcBY1v62ubBcfNw
vwTgmDIQD3dFCeLnZzHnNdk9PsvOTkUr/8vskwzEgE5DhU2LL/6PASW7oa0j/1PV
bxHhKimpxd3+uDcJWz70HiTNd0y3bjxGrxwce4FZt7Vc0o2nXe0NcbMDLt4XO55R
AywEM+4YdomVfJgJoZaTuh3FqJjEP2aEAltM1YBAOlcxb6hJp09kxk37wcaR0794
1Tj6QqzY3lxzwlo7XkojTjkfHT0hMPtY95GU8219spMo718hN/Hx9rWlLLXd9WuG
uIQX8fjG99C9oaCp5YxfLcE4MzxpYJGSIjcgVP7k1ytz3W44fgE97aanprhwkN+s
r2ji9cnALMsXBhtmY5luv66msfIxgRKB0rUBzD+41ZllsqrqKvy3kyE4V67x0CFa
47s8UBEiOlsKzzJIX3Q8IJWMlCshXGKFeuUTX1m4LtmTmZadQ1xSfbM8Ku4ATpi+
oOY8FIQVDDATG8PesKM3g1a8RW73uxTgQzBqzV7s0T1L9Yf61aweUObAX0DkYxXh
5O86pB8Qdgpb/hrK++M5lllDm7qa+XFOVSwI95Ds7Q/oBmoL4TgzwGQ+NLf/GcsD
oE3z8iy46B0gKI6+SjEcsQe4tOM7gnXkEk2hDpOWLx10/1izyWfPwBZQrGvqVRc8
eUdPisQmse/UyWLwT4T5Rw0HP8ODYE0LRhsfDk2QDfi/eaavG2JVzHA6G3XUcL3P
wTRJJYrInCApuWvoBMGS49hh7FimM96FWY5p0kiad0DeMDDZGhT8iFUJJg+VFvZg
riCS421TSF148AYD0hH7NHTJd4HSfslJ4LwhyhmxhrCZrJskZJa9g2PZ/1+G8YHl
vfGA0cs6XxHsB+lWBZC+B4PuuYKlsAhx74XrY+6tcqwYaNiHmRkbh1yxd/PgIO46
4UUzh5XY4LHnHRt2uCzAdUHt3iE42F9fQ5hbsAigSwsFYMEKobA6aw66BxJWT8Fc
I1/uAH6+yiAehzT64zNbOKZOZGA042YxDb0XV17jfH/g7Ysa4gmuz5YH9cWSYB6g
I28F+iY1pdrDOA3WG/y7lDwZYydismjKooPH+Bx8bSD43odBWO4AZGOEAHCabfdL
uY1KW3xLeUmrqxbPVfc0P1utbQS7h4qDfHODO+IsZzRpnCqWVajWMX+ZS7oxAEG3
KnUdWZovwup7xXji19vcWa1Nv/2lEVGvtkzSZqDPLaxJfeRB+49S/w8XCeDeiK4n
0CwOdMG0hvtgt4H2HQu5cKx7TEFZnS4C3L6xAIFijnUCFb0DiuHAgHUAr/5Tu4NP
74FGx45CXB8nrUQG0lSvZJDYfQuJT66PMbf9k8VLesWVV9RgwYNTw7WK1y36lnnu
PKeQZyg+cgJC4lLobba2lewskCVXg+uoOfl7HVtH+N0uY5pn0GYa1II/cnd/fleU
YhuSp7UAnE3BLkFCrNItQpEDy1Rfj+JphWL+J4Zc8/AENJziTlEkAufpjEZAAo2/
K6JNDuoyMuxDYu7E6d1xR4Tvm+tWAJVMSjjGGMXWh13+rkDjrhKwEWSez4hvixyS
l8VCEOcPQdUfrQf/gulX3iNxPxGGCbqJ6/8b+6pSYQnMTK1UthA8yl2KB8rV3U2j
qNDmhQfZnDifqNL7nXOSrLhA33LdFAWYkLsKI6RROiN717vTEHKT8LxEpdckxrC8
TSORQMUlQGzKkmDuG4P77N1nVUp7KwJ8dfkagKccZte+NyT0npyZvvQ/3WOXyi5a
ZrUH2Lblconc9RnGt9eOQzJrvrXya2Z48PdKxZmI+u4mjHifG+QAKi0J0Z8Iptms
3L01CDYs9JOX96Ug/eh+9MpwvCTJHDzCcr+MnH1wiadgydbJUlAdYv3TSNEcB/4B
hbxap7zkXb7rKdUCgQ+19ilmot4eDBSVYhVzBfWU1jnqiNV8OGe51XJjyIJ2kisY
fkqgNexiJaViKro0mfGsHJ4OCiYLgNOnLaBldZ87YVF3uUHpzKla6m4rgdFxAWXB
PJ4MQFDxHtTbxxQ5AzWMmVCcvpuRb2qHOMKrc9BlQy9W6Cbn3MaiJL1I395fzpZX
KBIhCENFwt2rRdr9iTIY5YYIjORxLCk2LaZUB9xujPQ5f8u3RbgjpMhlsizRC250
PjvffennWQdfsRqagFc3Eu997eLygYtp2NuCFi54XAC0+3eI9c3BcxwvmVjQMErW
Yec3WGrcqD2f4t38oujNYaL3wZRyddDEuPVBskGYzzEmpYMEy+5+rzafiKNgFr6I
7FRrGibs3wHHz4fDQprWmJ58gutq9iGpEuwOZYiZllVGv5jscYt0SJutcs6GmJ3r
qxJJ9Zwq7/I1yKWRXm+6vV5Icf/iBNxKNvqmuwpbzN3wDL4H9Q0YQOymgEVtlEE5
K94zAUwAhheSLbN7bZ8ESGGUeae0WSZQE2zijzUrIuZL/GGFRR37zG943fs5ydfZ
ZVUsXvCWB9kC+xgBwaZy3pxCH7dwONZ3He4DmRPcPGqlQuutCdK54kM2xb98WsLO
IcvGfTxYqg+0Hu/LvYHlGWiQ+ZTvt42+O9MWHuppIxAbkV6ZnMMy018usewceKOl
3RKqV6nhD+UIgHNoNAlvxWO/rsBFPx1AqWS1BgddeXILd484Cmdtor64PJJiv/a1
PQ/pHvWtti4mc4kYos/9lD+Mop0yqKVKT4CPlaMuGC0OJZBJscoLJbaPxDQmstq+
RyWifTmrBpYJpcthsIh2YY4PS31K+0r8hLhD6KGAjKFF+k5ChYlbHrSLxZ53br9X
e+2MT0H0eeqInkFfTLternf1x2h73+Cu9mW2T0hGKldwz8BTn6qZrdTRzRy6HKab
ROFOTIGndJ7muC87D/kxYTkGuzLtbwFw369Ze80LFI2yFlPPJU+1Gllfv8Q5ttQ0
fqF7MaMg4YdFwkMaOAVXbeM4YMNZgh1d4gbw0X//ooWoEMtn8Ih3i70sRvou1dWh
uBmlI8XYt1Ee3WcoDXFTDB1eVuIrwOhFmI9yaQf5qXSErkqKBvx9IiPDCW11Swxb
rwe1T3RBNRZPNFUNk9L34YjuyKaFzIBF/8GEbXzboL5eTCKChltPISDejUJEITOV
QIK1G6nY6d2uOU32b9CPjpRVoB4C4Eop8UUOm5l9IuTB/GmQTE6ipWeh73cIYrct
1vyKtn+jPWeSpNoxryISXhb8HpS26VQTUr/VRGKl8sCqxcBet5fI4SRKL9R82Mcd
bjDiLNU7up5qQJyJ9zImKa3JuqvdGntFcJstNrhZPq5J7DIWYmbLjlyHpG1Bw/oH
wuhl40ukeguyZEXHcpWe904o+kn+My5lEcQaEprhXStFQg667mTqNhq1wPxRxjtA
8lWHvqGv1/gHWIxZSnt7NvRUo1qBAsm8qAL9H4XNDvYGODiNt0v24MGDZGBHc0AQ
INDiDouVxsHPaeRaFv+V8yUZXmTimhJiNjj2w9wI0+YyKRzVDd+29vPlAMfT7+lK
rHZVp1VX/mv0xA9B2qGimogTpMQTm/6KGaXEZq8xKDXfkbsGAlV1jr3oPzqWKMze
QvcZjz57IqBN1P3PyCwHyWqM61oH6V4MWEYztTUGoC0YpoNPYjCfDQkQQXtu2sT3
wavl/h4U4mk5AWZk7Y8AMreEixflolhtLHeNgIIVECwRnwiUvieZLuREcIKDGQDl
3av176UrIm+kHtR65vHcqHgCwyFLLM3sbUieDDBBm6HI4AHlLcyWV/ba6GhDf2sG
MZ3xJ0HfHp6chXq7xSZuE6Fy4HrZEVHCGZ4Znks+mLWw9vdK+gEKXNC17mQXP+tX
O07iBSg+L2vlBA6axU4xoXXY1Fxt5HicrhVpPpQfCsu/BMxllg7gC8JYyUPqqD6E
D61R6MqZl+mfyQ213UcxDxGzTI0VBtkBGJvqDL8HCEa3KW2IlWIoHWDTjFH/jv8/
fWIX9e8yaWPvZJFK5qvb4s4w0LOSueXKfJ+gyMaSXGaQV2cLuGO0qssgi6pGndfQ
D7FQkath71nPLGONLP14+IUR3y7BwpYJx2FOPfdpNuT7NrBEq9KU0zkpqT1iY+2V
9s+g7ZPl9aWp34CsRTC849m9hqDtJNZz7vNgu4ueupb/E7xPnDgW+SINwjug22DU
0L/ENSEIlJL2PIsdS5fGtgsrNwX9w2J26z8eKuNYD03lutalJ3MENUrVa8YoqJST
xpKTRjFQDRRwEiJD6exeCg745hsIRPpBQKbe/fcU9/0ZSPWj1ud7mjtlKe50Ri6c
Q52y65y8jYxpm0sMPDGIogfzxFs0gE0O6wTrT6Z0EWGtNBx0bBgmjfC3FbTbUeeB
JZwqUmvSNO4PT36kWM+YcCHtlFDf1eaAW1uu/K5L/ARdcGoHXj6k96oNXRuWGPTx
DqzEPI5hQo3lABSa25coBojQjwh//NLpSqSG+ZG25xwhNtyP9Q+dlZjMyso2geUS
+KqwTmG8hmb15XNkmfFnHBtIehjkkaJ42n5oqkPMRm4V8c7YucmKHpy6f5/wxMzL
bjqIXo8d4MijLNvRzYsna0rgzfbCZnPe4lzbA7qEaedhLRtGjfTy53York4mOU7Z
HfjmgMcIgJUWYhyKAJWHRIndcCuMkFrX6tZoDHWGa8pUJps/SALv94l8UVqRvzhy
3+cFqwUFkpd33C7A6yF1qRIg9Ssl7Ihe14fYDFE+2Kei07gTb4iHRocwqhsTLnoD
QcqCEgIsXZlhMo4HSxSZWM/r/+stSF1W65I0BNMYTdHL8XXr/U5XDnRbaer4PD5C
KxiH/16OaHNSXmTuc3wEfwp9XAx9VhRqQtc2FtIjFHAK+n1Jr4k7lmUw/XGk9ghB
q4loLmSQTmFja4RFyrgti7r/VPBkSjhHhFnZt5OUw0weHFQHWtFKtSHKRjgFL7J0
QbMrwQOe2Z8BGzk08PSLecEFyKDcdtRSDApYSO20fUyvh8J5kT3bIcaS92v1yOwY
B82e+7lAQyHbdZN2Uwzxz8wRUEwnA65nysvZms9OBatwyuHYOfuxSa5oFjKaeRBk
ysBjE6vHi9Yga4+tXhujqRhPILcyfZWAeeZeou9tsqBO5AQCYsvTup8bcQ3VfHel
Qaal5REwWzopNudFKivlogQLNRy2zHBu12/OvPMLpp4bzBGLMuiYY9m2fsHK8m3S
1vvD9GHQgYCs6SDQRw9d9z/lueAm0AS2D9U5vdObLcn6qlYkW0jXe4m6s3l8VoGv
UVfo+fp530I9n/3H+yaYiWRj34wL4lRRtJ2Mkzswlk2WK1hnAhJx9+rqky/aXm9t
3H2ei7mZqCnYfARvV3NLy5LNFEUqZcvfjwmvaGcXsw0IUtahVF4FY04EW3AbyQeD
G3igDrJxsPZuCPtUvp1J7gzV848Wyiz5XbOEbkfShad0DbwiqcHA48b0DQxO9iGy
RS0Jzt9PY9w+WEfrhifD6ohKZA5LPmpaf2hzJ3D3HBRRnmTkuhdGqGJxd72EPq2F
Pde6/gEHhm1Wf2WmxjUT2INJdK6ejBpwnbyF4W+lnTFWxkvvTZuXbjT5kFg0egA7
E2env6CXjlVcLWsUeYIyC2MUY6ic6Qom5l6VRDGQBStNMi+mV2l7vBWYF1Q+5ix/
lvp0l7fX8T5zLSz7gJ+rD4citj0vFSJ4h9z00wqm4c35uOx7rywrTm3Z4KKtIHdv
dAiEMTFweNna3d6A4TEuRWHjYh6+YqWWGQ8Cs3rii86FNKUiby9eIn4CpUuG5lrg
FSsLl9Dw7qMRSeH88Tiqipi87SouhuXxoj3fsMcK0qoCMkVsywT+r2FFy4PbCtW1
JW8ZLQPhTjnKz8ONQUDvJBo1GPBlUoArt7L0BQ/0AUTOhAng+1/Rc++DzLL+qg+C
xKto0qepuNKMnVDzir51puXqAJDfvb9Dw8wlI+xxjdicyoLQK4OgrCkDXkjeD/iD
1Ds8MIrEL4gjMebkpBhd4S4fZr0Mu/PSC+hSJSOB+/FVAqI1e1mFMFd6x5m1VJRe
5Lbenq61kwACs901EIAA20X9c8B9X77R6I/S2twgT5yFS5BHkdVsmzW6uK7LcZUV
Jcd5vTXd7Eo+ffewGWjYLHaZvQ8oqwPUth9b+xbmwwCmSqbB1z7vAZQ3Y0uhPgk5
l8/5VgMqE4ayvbb7YwsU1egPzYUbcDHOCRzYKhOt4VsTbmspDW7Athg8UNR5WYzV
7Pa9lOpJ2WkvoN5jWrFseqF4CLvMocLSTiIWT7WwRSv3hUykHwjYJGqYNEPqKS0y
SbKq9tkJ0jBPhqd/VaHl8MlZepMKeCpNHNljeWcuRTS5iN3HaPMvDQf73rRVgL8N
5QvHmrB5lhnqajfPHlbaK8VtWVdlQ0eIzfAT4DqtPmzbjzLrn3Y2TDaZ+sC5F/hr
wIkCxDba6xB+otZsshKAKtgCHhaVHdoWoSmXJdU4ZryKYY61qdzWQpQ91QzuDoHw
IC+5Vrh+Jn9FSKQY3mJnWna3mZOU2Aqq84cZS9Eh/0vg4Xs2XZVcaXiyyziBXsT7
KN8S7XMCE0Ga6r2VE5OiwKazG7wlxGSjasJVMoBu1rFuGnnS58DOJOKxzQXfgxuF
3DxAB2qEpwzHWlkxbfAp2gpPKSweHS0rYOSLM/kWWkblChJZZqYPx0m4mdCzwx2Q
xjivA3IiQRrbcW6THOl7VO3wEoUhEHrAg4B7LPs5sJMEzktLWox/Y0yin/Xi6W/L
jB5ovHXc70hqKpIi/5raaG+D7O+0KfkXjzOddMwb1CJ9ijotLqIC5IlyVC3rv8en
5C4gDYuyrEIWJlaxaQQBM3nXR2/GfXRfs+nRLhDYhrKwZdNZ1+bUDdtzirTPETbS
VUz106Vb4JsA0VPdTg8YkT5FJD3m+bCV2hfEkE3cxq6edzTU//n+0FWCCxcjOPbu
uDWQQFVsswcM+NefX5kkaPa6M0OYWqwEYyvTe9rABBjV4gHIY41sxxlbd8zsLvho
nEA8uSKVcmlKJHwlMtav2hbwEO9L5TkcTMQL/w/24G9R9aTPJVkaX5V18n9MYkSM
uyTl6kDIrzvBjHW4VkV0DDhxwtUExp9PyY1QF8EaHa9VO9idxyd4S8z6IIz3uePS
73jcPD6xY7uTaUok3JqnvwJQhE828hBO5Da7DSyqGFgNEsIIGIhNAy/EoatOhQC6
N1dUgB5cxOax7FKDk1wlZPBcUmi2JQh+VzjVwLNNzxMvxUYMaIY1y/o85EE8KUDQ
8HWfK6rmDsnLdTYNW+UTXcoWQ863kcZyObCOLiGTAomkQHu+ucrN+MuUP5H4UzLL
q9hT+bmIDL2vsxlv1UqIVyDgO4tiSAP7eaEvklkabvrSE6JxNSFztLHGqmdVL4Ns
gh4DSxmpb3Lg9alHXtwOO4G/ONJNoN/YJ71XgDNxvEUQjFkPgaKyrraqNDdVYxCI
yDLpwY3kgGPhPDU5QnwKWb6U7S7xwn5miG5WrlAR2tzFeQRyNcahv5B2B/OQBJqX
BBLmaNQsWv71X0MUH6vmaeAPSrLZyXIQK0w1+WWJdGgIUTMfy2EoU50d1EnB9ip7
P+9Clm8cNNRFdB3rPSbzJKYKJHwDqy7nPj+bhOFBYufIohDV2mLgrITlV4A8epD6
BcFStLi6MsldoCDdEmfFEdQnZRSZoHKxvWUplXs8Z12l/zjiQhj/4aXdIYuTQODE
X1frF4O6ifFtewKDgkcgGdR2aDha3z2wCKISHBaysgFYiDWaNyc9DF+bzkKlAhfq
f3IDTu7njFyFG573n0F6GCXgOWBPzTirvrPqyF3xVYXRcRLiNdZx+JZosnQZLW83
VI42We07fJCx3GVNYe/HwKZPUYZC0HnTd5Rbo4gA3fDh8v7dfew6Ni2l9y9VpuLl
XbJpZewFQevuYom/VE4gCYtABCJvk27XHXm71WolZYmwkPalDizXvUog64fPY1QF
ozWe3FK0sckEwfdqPo7KDsOwRrvQA/XQU3lSjSvWc71Lv8EBp3E3TrHCrYws/S3S
ybGcYrb3xsAAHDtTRwmowNBcy/ExZv5TDQYgCltaDEK+MeFeb5tONVmYfxvDbIlz
RZ1gbIpzcbbbHDHh/YouS5AowYdNhlanCfgQySZdpgDw/PoyzzC29n45MbcjShPl
Ggc+5LToRjHLMCTx9CJKURNRFM6Ky5cYatnEP/Uh6jgyfsDTObgWxbCEhB2pyuzk
Pov/cLDw/YNr726JLo0/wADit7PZF7eXLRhKnd+XMMHWkFpfa7dZ7pdCB6sxpjv5
yEjzGI0gbfJKCXsjwNcSGZGhLqA5pJAeCIpcvWsIF2Pt5OJzdjQgyykipN9wBL6U
avJaYTCeF3v5jlYGglU8zQdD6MMGwTEcqfS34TOVM0qdpZUk15NKqdgIU6MqRd8M
NB5O0Ymb3547rJWPorhqr77ascgT3LN6/NUwujA2VHU9rRoOPXcIrlJWVY4CT+pb
vv9u6ZjpijE/JAXyaQrGjMpfa2G3LBk1x3MRN+UoJuEXzDIF7us2k4UMmXCITH6X
hzNWWax/P0Y8cApCPF3MXifYKq927O/gicb4cgAnTWRJkhrg2U+wklQrrXPBm144
rFRxn9sFdKhO7NwZBNfWD1iK9M9i/+oq8rUtNEuf1E80itVajvPjczj+idLaSXMX
SWQDPvIEF8Hw1IL4dmj+GgccREMFz8fKzyRWhX5AzvTPaIx1xPT+SPVMGplOoTsN
kA9KzFX4klN6IrINgddW4oJna76s6SbP8MYReMOPERUnSm/Gav/IfWS/cBGvlY7T
fawFuT1kQFy+ZhW4p3c/8sdcshwkfFURbghtB+bH3FB/+z+KUFEkC2skwfiqK3jb
TmbrdYa6M3CyjdoPXHUwqbKfMCEiR+ZAD7Gz5En34Y2QvdPa5l1IOMrTUt0IojLZ
zTQk/eadGt2ndNLbFCxc12oGdmESVsWanyUaBGHZP6Yzq9+4SsqBqbC8k2xqLBmH
OtQqNHlzdBr6kOHVh0AWhN4MPG0WdSVQbm4Orbkg4n445S5r3j7/g8bui61kpT6p
LhTrncI9IHP2Aheiobur4kU4FmRajtz8UmGvoBf120BGs+VsIKFO7GLj3tevPK89
onqilpjHGmxzUOY3OKavbEfUzKLedVc52bUB/IeHizT5uS7EchtX88yPjIAtST6c
VbBQcwe8DVtqZgr5MMT9s7vWqaGIS1ar9rP5gy5B2X9ZqhXJnwPl1Kw8zuc/m113
FhRAf8/TiXO4IAow8Wf4yhbYMKh8NXJ7ySxLdaUYSakXidGz0Q2egNtpZJPZCzfG
j/+kmh5uytXQhwwDJJRcj+Tqp4zz+RRdBDlu2fy9t1mDgVNvzaiSTxmDxhNPL9oB
ONQdjUXdw2crsVx+8tUc1hgn+W7e4qw9utPbtm+4D96nxm8tDdBfZF5PIHpmUe+X
QfautxkrOBcxZyKrmC65C33a2DP0Lp2+dtw9ZCa+84xtH79KIP9Xw+jfjFMV2Wl6
Zeoup7PKsy9Fjw3bIqVruEL+6Tr9QphavxjCRKl5y8xpOzQqx4RXUVuG0e+2f2/c
7QxoTbc2SxIPyqD/clcPzI3YWHSBJCIIHSUOCZjAp5nVdwXZPj3vVvGII68Fvb+z
nS4RJ4efe1QHcBIBUtiLADFMll1B/0gSI0DaDa1G4e8SJlkRGqSGKEP1ZY2OWHbo
b0aN8oEjzLmdlETuUgXdXQz35imaekQYdxTdbsYRBdZc5KctP5+UM4xMrniAQwWj
CARwvR5zHWqNmcnWHS2UqzGh3MlFzd4SQuPtgJH3HXLO9nmsd624UW8ubcVRaD25
tGN1cs08vsyHHPB2c38SGMt3fAc8IUVqzbUvWEjdyf+H8/C6JOWXIBJO9gjq9VM9
aAEZ8jjQyfZmy3t4MFq7t1mpw2mFmROCQGJgoVvCWZPCluf7wdJN7LAlnHwi6+xh
6NgFkde41BAJvjA94/hwZQEGn6j0Gf+5wuqCJUJwR/FxAM8rpqYPAVyQYLBF9/hT
jYqKMkM2mItKTXsGc6630qngBMTvVAbyPYn3sts9ary3hWpqw3dyK/jE0anT9+lo
1MZY3GWuO79Yl68KmfTR9DCJwItxS27xibFwwKE5Xxo6BZ7T0fEdXTZmD1paPQBS
Jsfc588+QKLm8YxoIUGdKdd0jqxFxaZEXQLGIcM7tJ2aPSni85Tj5dvpsBv8KA43
dnEBPdEtkvG3pCNZO/txjWzn3Er6xnyalRSiLmwWIEgw1YFn30Lns0vvRGSx/bpC
eSYIOp72f5RBXMdB6WWivhHVlCG7j9aGDBJo0CFRRgeJJ34z/vVAdMx+Du89Q2kA
LDiO0uhet0jZtaFG/E4H3R2SX1SshSJLZ0htaULrFC5tyZBeSFKxVALSVWStTG38
p8CA1czvEGNd0+Dusj4m1o0NQmAllZSFZ5qVehCYRe5SHK8J5YZQHrFglWxRWww/
0O7LCger5+n3JEHzXrmupTvUThZvyc0DKTXfLnLvhPEiRVd1VX+XMcu48Vo6Ebct
kVMECh1Eomyxt1pDsee+c+e58GkboO2oPO4we2mzEkYqM0QU7TVvfk0mOX6JVJuX
SKlGf92VMEDN7ZMv3SKcyasvm6ssx3iwNj2OlBikN2TJJpOYX5bg7ySJNzFWp6bJ
yYwqVxoH1Q3sXdnDtDDemgWPFrjS1ZlBPyyk69EvxmJlyuH5VYncOeKIDT1BxSiU
Nz28u2PZt4tIQX8QwWtqpwKMeYlvQSLiWwxNTTsNkSF8hjHP+5KAlmi5DJM+2Ujb
pN+LmaGauvL135MWr8D3qeAi3feHYtyj1jomhi29y3tjMKyxzzMuYj1U3TpIWUdD
mBQc8Hy2bjJjYY1gN3fqvsR1HWBoYxXPRIn02FM7M/7B5Bmj274k9K/HnszGmkED
GSs1x/ffE67RFpCd4Pa+kQ4cRCXFwcAjr+jD7pOy/ADNVJkKgT6VQTQpmiaotITX
ttF2UL0wEwmHVuaEPdfx/V5I7+ndtxeKgSX2caTC1CMu3bNxEJQXkYuPoYv4526b
A0WuNsI0phH0eTuTfQ0WNp3xT1BEsX9WrVGh4xT44sy2X9Q6xIv3rk/lKNArG4Do
OU7LEujv5rzOyMu2Q0YeZtSTxB6sHQonPBDovP04YA4H9KvOMRAUo4NeuOsRlVjp
NAo83jFAlWo9wXW79TtRiSbHUZonGWYPiEQS/iEdwo7yCSUdddIrxAw01OiDPzV7
Z136se1bCpdzn1rhphO4gIAHzEnmtWshg5Opw/kH6nWtA1iiIPC2DyJdI+lr7kP4
mRZZfnDF6r3ipOPfMu6gd113QiGPwm3Ug6MmGEYUK0Avoc22WIZThimM87YD6ti+
vsyVlJIIqCftz5D4ArUQgz5IhuMiYa0aUxfM1iYpF1fIsWAZ6Oh50Eyv9+X4PWlN
/9w2+n153pdcI3RWtVoiTJ6bz+tkqOBgGMV+N4LP5VzqIiRorHc8J3B0ALtD4b3A
+We6MbKCS0pEFNXpkr9WqQVRPu/jpEUpVaEwZkJAUo0SY1LiclN1eglOZIEYv1mR
YxOr4c8zkGLGHWMghtaWUM6dFdssyT6Tg0AjiS1Y3AOAfMJmwzFlpKLELP0Rj5NB
P8uDNA/F//UrZaDB1J+RHDWDBsVm3fllPNeMLBOm+kqlj198d4ybA0vf4GRpKCrM
Zw1X3GSXNmynl4IbBhIYQLehjtGcS/zkKF3mKhDqZe5DaAIzIZXznYYQAXdXVst/
O0FaLXXgUDklqiZ/nO0rlacV/AzH5cMw3GzGbtptpM9Lejgz+MVORSvRVtrzjbGU
j8KOzEfUxG8wZHctZhqhO1bokE2/suKitGBN8ROuJ/quB1lqsXBwn98hS/8aEDa+
zDHzIyPpQYZKt/zLd0Jmf9hrscSkfeH2XCm+m/mp8L6YpPaQyucmupEIKpjvhESr
kx9cCvaoEyHAKGpTgJWTgVi1gcMuQtUqDNU0OM8O6/nsDGsGoocZz4Svum7dSwZH
7064+nYwXX+DujTNi2mSqA4UocQUlco17iWN5FWLGDIZYlfZXO7Pd+QUTr0Amxle
0ltM6KEeVJa1uVWXwfbIdhT95SIIR19TygQSmUvCpM2x/Pbqa6J2NsZfr+JeXZX/
pZ9nhcjgw9MzznXMTrCDOQKoCqygY6acHJRRdkMqP9qbOaIdx4u5GDrOb6C0nAHm
RWLWOpPLTOdPvBIizveWG3lnwI2UAcGflMT3j0aaC6yAuu220qFoShqt4x3strAr
l161DzOmXJocH7oF2zphGm2YyauiO9XvexeTwjSixxJe+ojeU/cx2CyS1gIfMl/M
1/M/CdTqLkt/WZR1aRVkAhNX9Nu17QZyxlda6IhduwfzvI6P5i/LduHMWVnfHPQq
cKvu9WCek/Eswum3+HmOuPBSj9TAtQhDoU+bDqYGZZGOwT2E95nrf+xjP2XlppYx
VdPtRT/kpX4+eWtI0ECV2sU5svvGvNJBgcJIx+rP7HE97fSxMbeRohmYzHwwFkll
GVSFrJw6CgzWhWVaM+7SwckDbfKoZYEpcwzr7X5zCkGnjflxxBRiNcjVlrgHja0s
EUGUpVmMXPdUO0cUjqTkuEIdr0pDu1euSG16r6cdmFUcq7NHgdv8bMmWUFtCyJkh
c4NYNgbMcu/vD479+UaZ0/ftxHxijsmj/Zl0U0eCLWRlzvmtPlZwgsWzYJYAMb9g
gWzoBs8Addx4LXhjFAE3QJ2Gcq8F42P37tHgs2ahTavbzC92CRvxcqz4sdq2ZFtJ
5GBy1UnywWQ5+tj/5qHxwbruBOmtK4jaawEQHUtXcH180y45tLXFz2TBGC7C5ncY
B4wdAz4DpmrFOudCcKOXjmHnXfuxPqVl/m5qUInSYdiaQqEaawArI/BKxkOSrIlJ
DV/jZErlJsi/UFDYs/OVlutc1pycasBQHnpy8wVMF2zvUGbYrxSCX03ig5UYPk62
vG7dXdWfTcrWyl8zFcymwqj4/gXGu5G+b+UO4gjjSvrk6XNcKqxUEK2k78tMHqx3
++dQkux2nf9Aem+262GpGaAoebWk3vDA/si0LvnMjgfeH1dGrZx/8RqJyxg0AWNp
F4jXJKiUVWOaKJM21Q36A+xhv1NwwBW3kc+YMCk2I/llPN+0tcWWJsviR3crl5BC
Wj+FXiNdd58R5c2kz1+J7AC7Z/LMxmO/OyADsecIg3Fhs1V5mhugn1wRFvgIZFoy
lsXVnMKXmnLiqpJsda0NXuiw2sdw0tIKH7SuNw58xq71Q/QyDBHOuQVDhrKSe2Rr
5VlvA5W7ou9gW7OL19zvZfup88PTAX6kUFsn6A+hAXXwPwCSFfUxMo8Vwjk98vAo
Dsja22MKvqo0cippUcCV3hOWBPl9v73UFdEQz2J4gH3uWZ9CBjPgzEU2tkcj1n4N
s/E+fRxQjv+1EGLg7wKRNyUYX2vL0mbqvQbIrIXNRy3Av8wGJ46/KqVAwxQ+68yP
yFYO1TGPBNyzaZJ4pVx3g7xILbRohOvQohUaFioeaXgDbhK0od3Sz/0O/xC1+9rb
DQLm3FjNkXGjp6uqDYeCCgLMmCSko5dWw//97JZ2KGoaJHT6MJTXFcIL8lbYSi8V
YPcZlcVnuxCXm/wGi7AqNwpqJHFlY9tYp+AMrU4LGPsW1m/suRZCAJePdzVv5rvb
c3FYDkNBqFwYqVjELeWIlmdg26pnHjEw+y++rPd76cYW2sSt4LTp0+IZlrm3CF/a
Iy4iBMTerokdKMmXFT0yFt/gpdlONaG9WlPkgmMRChki9jQNjLbJbDnXpIMEz4kG
HfIfPG3Ivm30NlXtzkKoOdwtMDzzPVR8ZVzj0piQug13Rhp24mrTOVvelmm48Uui
Q6i32c2dXBZKOgbiV3gPUCamyQ6qvLYUaeNxeMEe00U+YmX1p3djtWFpEBDY5z4v
wy1rFthNKnA8GzGnQ4G6HE05FjTsA6n6WfqQt+rjL0Sz4V8yJTMo4w/o6v2vZMxv
rBw44haMQPmaiUS04IU+WkirNsD/jKHVYuQGQn5uklc4o3vdKBBoBxpsg7VXF0Em
tz5eAWrh/crx96pr/JQekfFTbstLk9QVBc/cRv+VPgHqUypxpPhHQO8AD6Afg27q
3NVQal19bxxP8jRBcHQWKJAkDY2Eovi5rURpRyWTAshE3maa+TIDQKUrSAOfcNvy
TkkgFQz0A4OuvxjuLHa58qf6mn+ldzzquHzJcgXgZRUQRhl63gP0A0ltPtmRLLY6
pVHohxz4TZ5vWgdG02zehaygFKmYtuaVQahcs+BtlL2ve4xT5Bx6b0XxTCYLkua2
WSnGLhvtdXFk4/7bAAUm/CLpNuV5Ml2nWxFcJb/an1nMxf1ExsL1s5trrvsgxMqI
Dr5RwctdPvHoWsFFOqdKpA1fYH8iO/x89MlZpe+sTMzxlFikSQT2eXHvLIpix1b6
9wXj5cZ9fmA63oKCHAQmb3EFzIlJ3kXz5qe2rc9YGnJvmhE0zmxB6m94FKR627Oc
s1/RIKGTmn5oAmLmRvK/8ct9CkuUUJx9Rkp7yy3MlHgA0o4xNZGH+KKAn6jV+Wy0
6+SOwkMZt+tkL6OUIVMJwJOUGLoMWXudvkEszxcq1hpnRabC/aadgjRAh3Zkzo3U
11aMUsRCDQXE19CGm+XWkp+W2S6H6bPh2A/y/dFIslopob6ALW2WKsfBt7/53mKb
s8+ph5cnZn1VI9vPzWImsHIeSwS2veOKzt68EjcNfd+ieiPP4iB3ujk+CjjHMBQF
XmizXyyhx+CUubjAaizqYza19k+ItYhx/SuTfGBqXGi7JC8a5rdCbAJMQRI86RF3
AbS11FyWqfIu9iyUEx4ICUwmnPLdyXljp0yG6SqB1z5gOmtHwR1D0uhHg8Cc1sW3
s3xij0Zoc4eePlQLogg75wb5KDZtd3lHN4jRpjxEasffKby4IJCofdtQNDDXsQne
Xtwh2ooDgaBnwubKnaJrmKz0/8OS11UGZXoagRkQWqxWbprb5PeAh8TkrCg4sZ6A
w/lzOdvXy6Mj+QWR+17jv5qlq2c+clKod/WkkBugMFtEzy878bfdD1906GHmOErO
iaIbBE7j0/8lItX4v02i3eDSfqT6fXyi/h7pfmtvgU6z0htyE35qa9bvA0g5yerv
Ko6UsuVgGBArmwEf97kun2RqdTFAGdFHYIvG1BubZ/ptRHUI2OvaBhp3tlBgim1V
1zkAStLOyuPNJOv7BIjNB1cCtKTvN7ZiWkrdmOfKEfq0x7GuX1lXpdcM6yzmZnSE
TGII5gPOtM3KVA2PTIafTcxdj9w+o3WOgfOehGdBf6rZh0in7444NMXxdeLDD4df
LH3qgMiB7YSRxrG5wcz+VTsucA6mBBUTFeI7nCf1oLs0xoQBb2kYf3P4xrr23xwY
1ZcborXrgw7745TBcHpMkMPAZWmF4XyGWTMvMkx5oTjMpevLmjm5U6KFIp5nFmet
siXC/i1KyXx0nJbclFd7Oa/2/nsmn0aGIfGeNC6pEQV7GhQj7PVYZUD4H9Mcx+CU
+FhUhslkXusG+VYO4dp/2VwDhh3Jk8HJ0tFflyZGyLIb64f529on6AWMTeeWkNYm
zC35FNVjpQXmNgaRD2+ca9ynWsTjMbEQ8ByYsCbLLlt7wsy7BonBQ5CEvp4w29RX
r6KRlhqo38a5oYH7YhpwrSqrh//Ck0KW0VHA32bCav1i/FYrs1luqQcpYC1HlbzX
lDUPm0oQ+wSwAqfK/yNGiqEhO+GweUDM+/Req7PkVqGUfjoUwui2rlc5dbn8YTWw
lPti+zlKzTI/6sGvpOEVQiugQ5ElRkf1UhmKLHab3usrXn4MiEyAps2EMctXxcU5
1msNoS910zOy/YxY8dT904t+jvN2z1PUbuAFDzCB6r/SnFMNJrScmEAewl/gaJTf
MNx7cwPcj3uuyz9CG9B87jxp3zhaP7p3QVxXMOWdpZ2ZSyPIg49PSlSMDt86Uvfa
sfV9UpZ65cQDxllgmgIHZvN9cF9by0nDvjglWK6CGpVThL3BY3eSQ2W61LK2GY6F
q6Ugt6ttxuvkM+xLHJBourllV2ubU9PMr+Xohnbbg7GWcA3M05dt3gqtBtWLfiU4
xQmVv95R45OPNWlQYciYf99eyO3lM8oo8ej94g0VBfqHkVMtqCr8GS8VQEF1WzGf
QsSi71zIUXle++Ug1beD9X5+4i3r6bh4lvsGzHQ+7FK1M3CyruYVVJMJMk0iC5fX
Wpv8FuBAZfHf9VYa+VbWuaB64fjNIONdiQ7Kq4iX3OhyRGsalvOMooTVS4CtNvA/
pgqZxHKNlLpiaq0Ee3EHBPIX+tcHTAT8d1dxoMcEql+GcjYEXGuKnfrO0Te6TxYj
m6rq4A0IoRym2FgVdoXtqQPEUbNUwfK13ACmfe0iSx/IQq7snlUCeoqtbvpsEHu4
JvS8RPucYVN+EVv8XNFWX//VBK0K6me5pzr7NVTBcNr7poLEF+N2R7tKbM0NYyfM
gzldOhT/qb54pyWH6sa0/mxFCRRB11S6Urjl+fcY0x1iDLnVaQlJn2jLAIBNYq7O
FbTZ7NlFDQiZ8/wwUyS6DUJXW/yCFmr3QNWVyBAGC25yFT3XDEW4EJsS2Y4G3j+c
ZMMPbPozDdm4jAhbsxvUIlQRXznjLcKO34j/cCMrhIPLCO4KBmCUOHiwScQBCsos
d09f4ezImLOfmw0MYSceteS6hSQXdFyj0ZsA8XCb3zTTsXbZ4ooVt/WKLUQ21kqr
x9cRVcVNHyEQufJ107YmH88jBofWm7qlOxTn57DITt2V+zEXND7oWJZuFd4wCoEV
nJIhKzRbuRglFavwRQz2OFBBhH7it0bfyIIG90Aczi469uLHzKUbJyb7518bnUGp
8Ez7sK1LxKh44pa/Acjxd1ClYUxhRhXbSx44wN3FuW5p38CpOI4RRlqTyAnYnR7E
buw0xrt9iacCSQLt+kEI/F4gFLI81t4p/Gyfn1EXybe29iVAbuQsLFGmE77p3LO7
yYQCx4LUmJ09kbT9Jn8vV8umPbZtjBh01ns2mr61DpHM0adi44tLInCgZCPSaZvq
tVU2CkD1lyhgSyurGd/+kUOG396/d5OzF2u0yYjMxJUvnqTna5D8u029HPXJFkPh
DlbMm3i8mQKjP4+M5/fpNsqoljCX3vxCIcXWo1/3tN7YIKXsSx2gUbI1q7QbhfNB
sEl58YW9iq7KDhe0U619coGSX9sngaptsAI8WA4ToAru9SmEaIj/HDj0JRFqqz/l
lTLGRvi1Zb8BXMjPte2y37bpmFWIPPO/9bEhrP257YOxHQYCwdIEMytWaiNYs4Vw
ZwdQWs/8qhVQixlHyLUELYT949D5S7BCcFhSX7Yy63ne/xPW5shVPn2247/pBx2q
rqtFkfP/mm4Gu8txwl71OgGD93RSD9XJVlkbOGgBv1QS7GSEViJXD+bPHVwYIdR1
/fQn9rvRt90HJYdmrQraUE/LI2ik6SBRaNw3LWuUnadzAS8Ms0ui5HLh0pGQekpc
chXVTr3Il46QyU9Fn9Ws9lLFz8Qn7nqjuR7HsIYoPngfeIShWAcrGA/o2s/ZYrxX
LXxPLeClieoZHMCdk0i1kQZWeuKikQHt7Wp0ClfdNFLMfpBLLVx8+gOKXrRahM9G
paUiD4VaZfIPyEaAPDCbf/8YShlbPZ8tJW88mCjkLo7jZBGWafwLRIb4svg3EOk2
3i3Gn70jtSRdtuo3t6Lg/WsuwsqwhV7O+rxeTqOQetxtSnmwMGuJUaneyxUKNstx
Umo5Y12R8hiQTDuDjT7Y/VH38Boce5Dfu/1wj7TsJl7PtXlLv7/AGCVNryk3BPfF
gNwapRegIdfDdBmZiNAwvcPFvAno73SeNuz+dzs8WIgQ0wQ1eDBwbuRUSdcKHjE4
CvF1yfM4w70bk0SlK3G+Nftk3ECrApjhHdtXP6nIeukTwd1D7H/MoF3lLFJZRyVm
hxiHfgkOLZ9Ua/q4bGvWATI4NrgB4+6V6BEZ8Wvh9ZsfRG1J2bGiGO9KKId6tPFx
IC8MJ/SjwQX/VAwdV304GZWbcxNBf8a0HhQOQKqgpbt6tfLvFA7NeMvowCFHkfWs
dcFxGH/cIj6aGQCSPzsqqmyonto9Na4PWN+yCgWPDcr0vqS+i80y/primXVkT7QW
kGhGkkq2QTxtR+S+NbS06STJgWANIJCPahWoegzf3V1XcTx3Z22AomWLr3E7hZh0
9qcvosjG84d+Tf2lyVj5Oke8/s2ac/ocblX4sBKM6SVEw17iDz2vztI+naFjNz1R
cQ5gJtgVG6RCpdy9cL3Jguo2cOg1gYANZ2JW5S47S0duhSqLucmzo9oCIqSkTT1L
2WvNdbJwD39izJ3ROmKb112FrFozthunz6FzCXlSvGPBxjFtxECmzULzIR+x2fpU
8xsQdpDhccUcD9P/i/2Mk+pbY7OBvdyCU5bti6Oew9JQdSDEROpW9YS3dEISiZ4J
AkVQL+KDseF00Bvw04AXbbSef5F0UN/J6+OQUr86J9bztetwMAQFZrqtqx0uDy1a
/d22OMatI0c5BnomRF47r7UjI8l9w3OzvfZ5E6/EG0xwSTO/36r0lh8JdcciRdt6
1fn0sgAAiPlBXt8EAntgSjLZENvyclnrAuO+psN9qpvx45cIil/4T5hkoRYJlU4h
2RGzzmeE+OTzWBFGwW8cbEwPyDdNzvqpDKZZuQjztBoubC4tM6Kb6B25/Id8PVTZ
TSlf4vyf9dRa4p9AWLT9sL3wGV1U7FpvIVwa9j0eZkKbXWiF/9sHLh4CF5BQN+u3
m52x90Rikt83VNyFO6SuWA1wcv/qIKrm1xn8j2DWcSTdeESn1kCPTmSZWKMQ/xF7
hxKeoTazrbrn8ATr6u2BbTgU0pQIGS/5vcv5D5yA70hwSB1N818ntFebvUbnSR4a
eTPWudFm8a98Bj3UXXVW7mWDtoBbhPVLyFUeOX7CHxHK5070HDsK59b141b9f51u
Lv2b5SlCe+MRzEaElS5shD1zLK7ds9MEKuZLb3qHfHKYcQdLZiYgLmLCfWnkTmMs
hTgQIZdURhoGh5bXITonAOvvTTbbrBnYvXFjO1JSlDvPmiX6duaFiPX32PmcmDzE
NfhpHTg5bpBbM7Gm/Wv2nIADMnrubDFe3woc+EpD12JUlcloZE3jTP/UpZ8p2AnJ
BypvLG880hQwnYOHoB+Q+pVECN3+GouKhDRYC/GEta/pQyN+f6ydvspfX6OiBg2j
6gLLZX4fLJvKnFDXRZ+o019hutKU6A6XgLrhlMNcUDH+qmBviSuCCkbXYLn+sD2J
qkFocTIcStOaZj9qpegxmFcL8Q2Fe3mppyKBwKHryp8/5gERybU3bu8EbsMXqCl5
QisqOVon6pblYsUaY6XbswD910ytvlS0PYAuvZmVWynp0BKV56dW4hDgccDgR3XJ
ZGXlRFmUOzsEbe8HykTsETTgCAlzG+mnTIY3E6FO3rVqFy25y1aZ5PlZkPpgcRWh
1MWZWqJXBNQehJ8gLmdGYm2Axn6jY9FjVLaV5NE/qtx2HWvlzB6mof2bZhQOiteC
y+0Ag7D/4RYOjfp2HhlCd21g4cej4dZDWYCheeOBXrAhiezSMT1K0NjOfvNhBX7k
WKdhi4vEk9N288x9Zfl8q7DR2onVz02sfLmEeENE5dz3rptXY3GwOlzVw5dis9dQ
DrYIVrhvHtUHisO1PTQTeJLBtHkpdRi9uuNiSFptzDD0tacWKUFbopyoayZOKHVL
sfnc2ySiJrENzYdC4S8CmBjjUrstbHoFxFtEF0cSfVB6wrxNwAFCH2K8B+FVXXB5
WqiB9PokFabVDzWPOSlFy1+lBTnzy/6l2Z7sN1M4S4skLL/6NvPPA8RH+C0mR/er
L6cZiCDsSsSjr8Bakex+g2qZAjDmqXZHA6XHNnhVqrMlXMQ9f5xUyMfddMNOj2Vl
ZDA+kOgTp3qTWYubt48Mn3LNaMjsAufbN2Y+oDtA/KNF/gIMJQzd5anbtrzhKY12
VMZBvDsyxtiqEzXuasV/P/TwW61oO8+Tr/YMUwOkWoUwhi0DXSnSFX3Ek0+ABiG+
6sRHSxRJwrgEFb8X+Pp6zZggVYZtfFL4WWSrZYQHDqoH/Q1M8XtpoW9RKKYqLd24
icgIAbjN7JtKdRy/vB+BDpmNZ+KWYwuQ1kvuXdlg0JsaE5mBuP2s4IKGnSnbduOH
VsSeLd+v937prK/pCyxS69yWdcRLYX7vO5yPFTTAKKvz3Gpa0fds0/tT+WmJfBcd
Ispd1kAF8woZ1AVdiFh0iPZDTH4xhnyWtruVDNU+ybyYbU7EJwcGLbkHxGmXa0F3
ZKjhn3AdZJyS01GB41DDOsUAdHuWGdDW/j3JBrU2it2RxivrbLyC3GoZaAuSkTfa
OjI+Zv42yir4TLFAn95wX4LJZsgpBd3d+FPQPKA5xtwwXwil3Vk8PhVw7pQMXVC4
jtqzR/Q6MTPUPlsq+mQevY/m8OSSiS2TJU8m3LUZmF/eWjx23rCtDY1dAb6KDEC6
SA5I4bP19vpqc9ygHfDXHnZXJ7M7BI4712YNrt5caFJQDsHilX8S+WBxz08NEK02
ZlGh8KID2hvMBf7Yu6E8vhp6EvY6pmt+i2wY2cODnDt3RYP4gmFUSIeAlPagujJy
NqRMrIFFkjtk+WNrW7Tho3wOxqYeNMXEXmm7ZxpszMPXDKk5u1znNwI5OcG6E3J6
uqhpKv4gDbQuH/SjP1ocPwmlZlQVpUNtRXTJ0DLJIHyo7vScJ6kfgytpBpFrYaMh
TYhu6TyYRFtUBfhG2FaG0qt+HIaU6Q4P3jeb+hMo+Ssl1bQO0Lofn6t0PZon3BmQ
nGql5PzD9CTbiEqVBTqNMNchiUm4faZ08XaF+L5Uo0FsR0Wm9+dtVGvowwyZ13iD
qa9pgMm4Y9w1Uo4cpCLp1fvVsxF5D3oybCNLaS9w0gz7yC7VZX18D3Rr1tb2gUhj
4Q+xxOyhE7hITSJjWwgAIzWhnIWWq5Luscmvk0ZMvCJW5x9krrP2Km6duevqX35l
4LkqpE+AztBYA9uTJr+JcU93hcvflCiUFZLr5BUiByeFS6aBrghKkROBddLoODsA
46aJlnZxdP8S31EYl3km9oiktNdRXm7dxxXD8l8bmDUNrPJyMBW5rkv0rr+N4ntS
dl2edrlyaGu6Cl+tI5MjnWJhoOgLUCRJQyIVMBNNSUbXvFZKf4aHdCrTuawa2qgb
q+7/xb8bWHvKlSQT7Mbq0QP7ffpAzUpodj6xhOHqG7FdCBFwKuXv8hivPqNS9Wvg
vMReKePydXUQe2cEiOH4XcFdPsZMIXpHn5RsnEfCzxRe1LfbaA6YVD0TZbWd7Pom
GmttGM/8JpSmNGW2YROSamzNPQ3Hc+UjDmh9na2V1owsDDv63RlWFjCw7iYRuZnt
4uUdJKQHcj83tWEx4uJHjAaarkVFLdWHGTOTkQk7AQO232vt2Ii2udLjiUeYm25v
6Rox/R89heRVFTpFq8V4pddTCmKLt3EVT/CMb0w0c5uT2iXV7nbTAkqyOYeNrRIc
w42NuTQb02IMMag40iaCgUYRm4QQCOx0QRMKrUQ0dmpkXgShGaZLXbqkqKAJAfqq
gG+QQJ1EtY/YAVcXPbX9gBb4LfO5N1k0y4lfZhegQXgmb48fRnflcg8DjzxehX1W
Y0mocHEAtw+RfqX6siXQ7GxpnkxWS8KmzKv73FXeYeUQSX8V7RG+wGsQPA8RVufK
EcrfimRKeqZ5F5lLIQoDWAta3UoeB0yfZgqpcct+6wyNd+2PRzr786vc9fZgTbCs
x9u01YaECCUgjCPrQ5YayeidieRs7mamgIAlT+17cUghGJqKDDAYAZRyDAniKwxW
Jv/MP1aW4t/yvN1Q5/Ua6zoqaZBVFH4rBSa5KQMGbZOw4RLnv49O+xcQ2J1nUn9K
LC9wDZ71zV02F/o2VXiDXueWYmQQX/edh0LVSvVDb2m9RWIhCUTyb03fqph7PF+Q
pf78z95mI5WW7Te0SwUXpacA7blcNyqrMVkYKgx/mn6U4iqLtXEj5mVK6ppjGLpH
latwafZWjP72vwsxDZShSQQZqfhVnXadEB4grefkTLMiOH5Kv0QoDwHI1hTPhSXU
NN517xy3e+j1FENz4d5TG4XOLA2ZUGt5L7RGErqoxs6UUtfkSR1PbCldbO7m3qh/
YNkTCftROraCMqbrjIUoLWyK3JnImYndi78Epl5LxOYx1WQjVwtgRd5mGG0eEdcz
MaswHU6jnUvJjfsrv5dBQrYJT7t/M48zWP51FthPulPHLSOAtWc9HqFY6Dv15NEG
dvl/GSiBZ4bbssNtodN0SKi47iClLqPnzrnZUUAHEPQQsQyC93bcsAzM6LMOzXuL
sqHiwIef+ezxR/7GMHrE20VHZ3I3zhTlN72Rk7fyxs9eNZtOD+PUu/HX8GAszDsM
GSM3CuDVfCLG1kvAv17jtri0jAOis4Em6iwZ3+xj1PYSu1RsBH7yRigqYce6blS4
2GWdbxrLJjVKW6eY/HVAY8+xZx2L0ho324Mv9uRdeTp6IaKBbAfTwxCDcJg1A0AO
PtPyo6Mrr/V8rjZoOUCEj7GZ9TxCiXaBXUFkOuUO7Smf3igPFGC9buSOiOcpgRfY
L9vSKZcma73ChBeGZwOctm1EhyKsPXLV1/X20lDpKXWjQJ+GNORFfmPnJphxnDVd
gQayY8ISn/tGC3DAnNr+3T2UFLdbMgoQDpUZOOzPxEZATHGvkubPG6XiSsyi8Od0
aM8FT3eef6cxpP3pavg+qkTo/agkbc+3Rp9WgrPzrkTDUjFYW0Wr0d/GIqylecZj
ZGP4GlP1u0+hqW0HudmqbyRUdHPD0+EKjQI/lT+MPhUz1Kl8KzLqHfNsKM2C9v8Z
v5ExWfwaOP3BrVnAwhsGYf/6V8S7+s5UJ5uf8/PtNWkOV0ude0ltvP5MQNERiP0P
Z0EWs72qY7wLgbIsWxmyZp5So0n3VKjIqibsBqAkFJwyL/JY0vpsgg5QRxm15EXJ
kSylzzUlEo9se97xQwVmi5DAJonNMX6gieSKf4Inx7mFsk3TvoOv+kqTf0S3CdyS
AXAV33W6X0NdZ0izk0n6+dMyCJ1jxM0F5+99wxU2YsYusJDo2dHWR0jFTsGIaJEL
Uo6chYKE91Stjaac23Jk9C/vEqPjZI6e9EVSyE7totbOGT+vlZtha7MTHNMBoQQP
Q7ZEQ/H9RtDLRHha4NhD7neyRq9kktRt+9P4SUT+eBPigF/osjdx75K3/5nvBxsT
IwEhejjnENMvkHQbthKpPoiCWVdOEISasVjAtTI6LFxK0hXpvJuavZLa4HYCkmQ0
8V3TsLDX6sIsqruedu1jcdhF3D03Xbeji8wFEGEm27UZobdEafxP+VqU943p5+no
JMKHgy6CU+xXqdU4tsck/U8mRiNVbffn2tjh/cuDbyOfi9HwKldrxSUSTtdYJTjt
VavocgT6yltrZNk6h7zY4PrlP5pmmMDtQ4rypq0q7OZISY0ei6C8J7740DqO8JqF
hjDswFEnUA3+c/Sfq5CG/TUmvE8b4+vJhRFblC4S3PwGWR5ivIEVIdbMlLHO4DI5
PpZZhDgVET5a3veLx86l+Tc+oZxjpQSxLB4Gm+M95QcPa5zTujRLykPRRjC0wwm6
GatGx/LvO1OrNdhX3noinIOLziab0XRDUBVRQUmP4WomrNebsf8g68yDKyNUnQvw
7fQl1Gau7/4wYSPrEDHxyD8e7BI4kgaxkazI5sfAKnSsZSQb0ut4Esih/gI1hIRA
THy2QrtPHe2B2xoM+93QQ/4mFOK0tqf5OukYFDmI60hnA4/O6aKs/DogsMmQW/qt
czgz/7oNEwRsJoGqyyXzsgT1rjHZbenWtn+NsG0f+E66jbXvJqZiSvL7+LptGM9U
2ZDqVUVFWU4NPc4OAaocA7LTaJircML7vRi2MQdZ6S7pEvyPs58pSmbI3GwXvfhv
Yo0A1J4GinfShjYD25bdpmm9Ikjes0U8tPmBqrscz7DklQoEKcp7O4uMazKyxNeR
8+r5OJnvibwR9/RzjPUqrcW2RJUJ70WT2UJpot3g6STIqpN/vDOY2RSy86x3tBJA
FbYv7UKd055ttj+dRiEOibyxN9BKXZQiifk0XxBBNBabqNy3yDDx00pgkWGzi491
o3AzLFp6Vi7jB2wZpMm4oWU3/uahuYzOQnH287xX7JalMkCV54hXfcuzjZbqnEw2
Hj9VcmEJXMZRHodrdxFBnUecnOEbodzvrXm7OSjwS5PJDmYtrI+OU5MdZYGWl98t
BZEqSFCy+IoE4UnPqDuHLftdfoT1Tc2SO8y9ea/nDZcIzS69JbCU198IZrDnAJYC
cRm/z9sDUO4Zv/J4enhdJtPJN7AnhIl7axywslOwYKQEU/3DnP5ZRRqUQUQNo7Yz
3r4LVWFEZWIYdkm44XWHjr3wVrRK7AbtUc/lo3LMkNwG1xhsIIipRMX41rRbZU2C
u/hnqmtCdF6+JG+54g++wCXARpvmp3WSdyh/lrIn6pNQWra98bHi2fRXX1epuu36
DQsg7frjmpkt8VNXbbWmdjjXwms/XDdZR5NHFo9Oh4gSFiGhZUYWfH59VDRwHvD3
KEN6YH8O+iic7kkNZSZyxSONIIYrBArNF3sNMtDeXrVJcAX4K9+kD+txh2sz7WSn
i7wFLpcHBKmUKokIsGxa1wqTtifOyDpwrpxVUmipy+4S6wEvaSB2sy53zRirFSAr
rqXB3jsf6RAkeZfGEnEnTKKdM09j+SNyZ7J/VTGm2FZNWXHYqQHD4gXf133Cwyf/
sZ7TYOjS2Bri9N/cUc/SGbh5O3jtau5BfHOW/VnlzbINaxiANhb4Av/mJmJzC+Dt
OvgZrR8kfNZRhbwc9/CP5SewTvyLSCEuj8xjHY/eByP3KM5obcmyy9JnZI4NtWrD
O3GZKUWB2MRbuSXjOWwK2/RYdzH6X78vocMj7uVhNyoWOsavv3xRloa5jhfpGGRS
ZEg/ehTtFYbKea2TB5eDjZM+rwBVPeidzFWvBqSxGmKRxNjn5yQFlDlnpLTQOHN+
fTu6lLsqzfk/H9wI4bl2k5nAYo9M9rvmU/JldWBOi8RH4m/1042vRGNw0dbyzt0C
6uQbh12BfNAupqF/NIOVzlH7og7bFDEADnQy9hR1oPdNodkAYlc5E52JGboa9c47
UKlziBJgwbREJ9SazsgDgacnu5s+6Y7Ek9sI5k+JLfc98inQBkuzxOAfT5z6tZav
VMcYJ5H05hzt25xKJ6knfwHkUrPjopqsIZKCY4ATNdL9uq0ZJ4b1qydESL8PD3MZ
h9OV0Ko6dH9tzXmeVPoU17ijIoQfVJEC3QTOVeReuy/yppdBrjcIO1fDiP3Znq5A
isR7OEj0PxX5F4+4qeMmMXfui91bFX+PY7sLZYXgyO0+u+UnBbv9YZGvOMA7tMNW
B1toIJRSx0Pll/GWFp/s5TL6L9FKvRB8JKzn4CXr4YNS6oXbsn52ULSLW+wAGW4v
7pV73mg5BKMRjN4bNIkLfBi8Z0lobpfNla5Icnw7khgCWepfwJDV7jEeuj1VNtCg
+C+vFKOBfvti2o73G0kyatdZrUzNU6kdV6gagBF3lVwSTz+EuZT6vKnzSysM31XI
XQS0gzsrMSNzZ7rouCbgAHbw/0JY9Zu+6Q7BfDKuCWq5JC6l9Aat7yUwIlKI7pbp
rBauq0CKlAENUfHiu0jDL98qI7aCr/gIFwWh79uO1Le7Clh0qZCtsG9J4Iuhpix5
Rr0feunGZpoBVYP/7BvIdQakW/dwxDatwTBbhn4+xNaWfo4Bnhs7PKtiKDUbvtTO
BJH0yQ0r47zbvUh4h1sLEjZO5QpK7dqeoP8/0ohQv2h52I6IhQdp6tnqpVK4sBTo
Ppq6BskVr3sJEUy/QVkA3lsIUOqedFkuqAcWjYliiQa780G32+GACBxubHBfOdi/
CwjF6rItXhekB7y0r0mf6Q7mtWSBCTfTnXOmxBSY4iYTIkCnonBgNtJ5xlKHqVBe
spzOBNYgndhGag/MXNLInGhCKj/T1G30u2awnFXHtKrDIZ0e1Vheqo8rXU7vb4Zn
qXONYJnbZzPyFwvrtc9djHP/7cpnSJaaVi9oC1NG0nm8mNbBf3bV41ksR4wNdvgJ
x5Dx+v+DHmSwsUQTYnnY+AxLaRhVpccjELX27T1kPOnErQqvEUbdOIc6JT+8QCCI
+LzJr8ENDO3lOq7t2zIPYxSPGjYPFq2LUTog7is+0MJ3hw4k/d2W5WUIH4dfEKfP
gaxAqR7U8wAVRlPDu/3kAoldGXDr3bvbruqe25iohvHl/NMTUKvktavTr+4YAtK1
CIE3Qet2CjtyAh+eOaVvtOD9Q3zZ8pC1Frzb+14irmu6saUD1oemf8dkqaxAFYjW
BjXecWfh6nQAmMxCeFhjgqjbJ4KU5zNEcm7+KnEnfdRpNW4uc7ANjId6wD/eQPYP
WmwIxWoDBAfRli7sGC/gnlPX306glXYaZlTdajhVZK/U8ZjZglDYl+Jtjqo6CRz2
rxAgqfBpCGTWuHLAsiTEYWDcCUmyXOGQ9va3M8j7Y58rM8YfdkRrEV3ebQq0M9uw
vjFuCIFphj/r3RGkUZX5GSDuOL463CO9WD2r04aPQGt8NnAfnQvVv/npJpPQSJWD
8fRdnnvVvwWsqPNsPKTtftpo3f97UwnaleYDW5/gFztE1nUSSS0puuzARqD9jHER
lHDSmH2OUsrGUnCYuynQ14PAQ8TXhRak2PrgYOzBNDi7Bw5I8DkMuMHYqQ1KJ/ho
NCQdJG9sJNdqK+nJzOfzrzBdOTPMUOJha1lEKNTj2Tvd0Tj4ZuyoLSteUcDnqEsK
2Q1xKF523KYIHVHZX+bHDGfPWL0KMR7CCRqPxioB8oJyNPfsRnPqHva8cnMkSaqh
swxjxZZye7URHBdhbW+xI/8R7dovfBgqzZGvJxv6O7wapnIfAmHGhGTQscsN5gRR
fVXpi65SULfC68AkjgUT5V5B961cXkJVGVypQk2A8ymBuY8yIg/zoqQT78ffd5we
uhBLC4ltAvLqMEgWXrI5TrJjK1gEoVsVsYj9MN4VcWx2Ado+qhcxQcT1szUYr+TU
qplFbjw6/nDMKvhbL25gDT4O3VuJmSEYIDfqvpuYH/uWUNRUprh9ePPc/HzCGf6m
qD17QW9+s1yRJqnkqUlcri/Ua0aUUkuI3aEk90igHzZAS17tTaKvOXBsVdH1lDjv
lXStpUbqUTlA2l1P0AoOZGZ1QoF9f2YJr3SjULDwy34xb4i/PqTbdgc9RGJiXoUr
TZGjCywYJvd5HSl/4MbHAK2FjsQG7nUdssDfTEtvmHJJSN4ALwIhIop/eXQZbtXY
dA3wUvxxgmThDK0lbp7vgN4DQdNQZyfMEdIjlBoGKCx5kY2KIXup48cxkWMYgqFw
a40HKsB7iBBmG4nJMicspu10Iv3x/H5UtehYgwlwrfYB5jhCMF7ZDubMFF0vMmVw
p+2UesH515yuFEYD7UBrq68njrZaZRXPnB2lI9FhSzdOjlu+sEEjj01LRIGJoNR7
w4EE7EEEa4JjLw0qXkbDJr+ipZ2hKeA8EthKMS+buA0A9XbKgxdmdSY9+e+mqn0x
SFwxol2PhsbKvBukJEkP8E8PPfqwUV0809hNSe6d59eogCfHHyYX2gHXZ2HICWqp
sYzFYJ3+Cwiq+svYFq02DFeQr7y+jUNNHzf3kt70nToBwJIkSMmH7cGk7FCb9JRm
dDCgSq2qBwWj3jeTZLFUqpr1KA3fhS0C4gaEnDoBpIGj2PzHfdCfV1dmN0a0eaUv
t2RlTA+BqvfkCxheOYvlrk4U9b+C1TKzgbkSsPyk1Y0JA7tVM5U1qy50sLqQT33R
Z/mahVmtZ39n+Q2PZeqM49QUqXN2KX8puPNeeRapLG0f82dvTM2hzGW/ZuuKvrke
Xy2ZjMxk2AXRY3RqnBd2nrWMpTmjsFm6nfBNEoWeTIuYJqrp1dohu5BUtjavuAXc
CXWIaLXTWQDDPjQ6FVX4i8qXQho81vDca+LY6TwXLJjuSMq4EYvt/wfxhxR246uU
MnlO/ZAKrmJZEkGk3JRUdQoarZliWg/Kjy5Ymrkbj5pK+hpyiKW86syu5uMi+oes
gnHKpAUseqvVbbgz/9xeuFZnxa+ATnWGTtiogJdHSjMd/FyJDTmBt41ENwh6CIwQ
M4hhW911cNpMqJ+LwzyvPUjQEpLHJe7JwRKBvJGsKyKUTCByMMotJE35TiZZsO7Q
lBDcUv7h7i1BDKO+PiqUf+wg+rxlp9M0svElmVXRItw6VHOCMo0+AUF+us3h/X7o
3tONaFM/FlS3RKuxY/sYrGF93DQIZElUTw4QWI7zRlxnW52iX1TNJPiRXpjf+Lu0
HZdN4cqaHnkO2silYrc6hNk4yMqA5C/Ae6Unb1mvcWi70XFdSj7kBaxzaJ95hDJp
a+eyfYkJJ0R1aiB3T3/0WM1xp9QRc59QFKKGNYmg8w17+VolwQ3sTua0iElwmYAg
o1hMYGIcruqkWDNZOU81w1cHcfVQQ7ry9rIOXfK9FaYZjizKyNW2RUAppul2WkeL
IwfLT1DYtoxL/tUyb7+jGrk8BYzrROyXEU4i1r8f2es8yhLg98RgKZZiUKrCgrWz
4aCalJY6KePE7hK2LQZrM1SRIIVgWiFUKqDRVcI1MkqzrRTG4tCPUBEFi3qUZSIH
mHOrDn4gWD06eAKbgq0OcQCl8B3axMCcZaHkdBUIPMjHatXd+JcGQgDcSESwY1ib
RiDLrRkprTSPlq8yntHzWcZoDzZOwQAJb9XgeJ1UaUp/h2qz2NCi9MsRM4UJDgJh
WvwtCqQQoQl8nKy9UFBfOBBnjnkH+NcIQQzHiKInDhaVH+Os6jBGWsprxTre71p0
La5IMrtIZNFqLKFiKJI7k05GLZNX6Ev+CqM9WwZGxgKmfAqchb4FKd6RRgcL4g2N
lbafyOuXL7+ENWcidBxG8VugoFLJO+d7kKb5LGoUion0irXnSyrtLCY2pMZL+AUV
pbEZzSWnUuQ8vbAhAL+xMCNgQiv5kPBZ+oqNq5lW1ODpK5gdjFKKc0VMfjMXXbxb
1Vdyj2CsWrcu5sLzAQrL/9cW9wb2tXXSUGhtzEhk83EouYHSJd4wVK5EHoNpAAC7
+m0Hki4peSIbdIoNWJvSPT91uhbL1olCCoB8+FAHLij6pNZIzS+uCDv7zMo61nBv
lixz9fi2XDr7OBdJcdO6vGtY+5AX1DQ6JBAG/yfffe5MWf4HvlNhhUEerBvarsXm
wXQQ/3GWqzeF8+pYvR2fuacsD5yK7dpe2yUuZZJAQWDYpJoRb8+CEJEIFIouP0cz
PIWaJND0jN9l5ysq0UXmilZHLnLqsuznDqhC6s59DF1QqvQtjW8OoIJtv41tzTQX
wrIIxa7m4qBoz2IT7/fGEgAGoHCt08abM7Cw0Dkz5KoXgXx0dWUt1FW8/o3Jwknz
o5NsNAvbwWtC6MMm2jyvHAAmwpWi6PzH/qdLEkQuAGwrYBbQGTp0Zcjz3VUeDmjx
2Z0tAvf3w42s5Qq9+3ZqhtiNtP1BXJ8QQlOomkOYZ9T+awg8FBa1YOgHSrAI8EZO
+8liQOF3SBS+xGQDTpeptzhZPXoUXQjNb/AeN6qxmuDzThsX1/tSgzsLrTwPmIGH
/7hdpUKYJbJSQWcSWkn42pOcVd9h11lMKJTqNc1evR9E63GCSeuRTxDK2q8u32qU
kH4+aZ3KCD8wghI030bG4BDdL5W3saumyPzv1kl8gwNI103YFIuAmZWdWqDZXOD0
s6InIaF+VSmtAZQhTqhSFuAzbXJSFW4k2j33sZWiCHYSVvMUkEa+CdoRqfSIB2Rb
M5GPIzB88kJFBuHMm2dWT4+/CNHqywde/e/TSLyhPdLSV3ND2Y8mBvKfheazK2Ni
uz56JT5lQvNkclZFsUT5O5I6b7l14mkd8rtK+BAqvUNlzpT5fxcECrRy6Wa4G8ar
WVZp6dk0/uE0o/TShj+34/Y7CyYcYOkqmvR73/q/Jaj2onWNo0eN+DTqNX/4W6Yu
ktmIGFmaeLZfNdknwuBPhYfS7qr0jYRG5IRk+bSKMU/sVNK9fdKCCjSYDds2aHhI
q83yJ9pHrYIntt5VXQgXurqO830oLQHAKB72GGtmAkWn50EVU+FSfUK3iH744y0r
QSnq3mMZoX7iieguHYhQjmn4ttQqsmPcHX7oLsmniW+3bfXng3PN4rQsmFq2jw9e
5fW1mFowRKriFjh/nmOw9yOBfsVuwXdjQBa6Hi/w7ycmvSzYBurxxYYxw6VnMazX
sKnuVVRUtNfAN/pxl6VuVG6awgyOcb0Qj0nh7ptYkgiIkiEaGIm2EsSDxkdfTvYI
cP2gQfnJtgIvWZ8W6Rew3T4XYPqmdXc3CSt4n93etU2mUdVM1q9QnREh/mID1F94
TDsEU+d4SlzSGxHJpOcarT0P2cS5q6GsYX5ugilcp3nzUCIGJ8TeT00qJ8ro6e8N
w62d6Fi5PecamPpDKH8IXinWuWvzG/7elUTMdtj4/ZSkQ/5JL8I+H7og3YX4IolZ
mEbKNfVSzzHojyCi+A7MkXP8MFGBkGHRgYDaI9laqQ32gH8lakHY2ZIRhyV9LQBt
ulwZyQv8e8VrVWO4kVHen0mmuqj6mc7aM3TEyMGb3OmkU5pcCDMpM5yZwg+C09GF
QHXObWZ70T109flPdOkQFpe1Hmp0ekQTjdvp94qYKM8aw3e3g/my6enweQLPPKKY
Sex089vTg6Vg5MtSNKMY6SarzX+Op8H11U1gqsjBKfngO/OXV/+WIQbNhTiCcZdR
lapNwabxtzlRrnYDGGnFRSOOUXbjTBhnB0hVAx0FUQwoSNbhf3Pr44pt7U/A0Wdl
4m2MB7TEjgpD2HaNlCTivqqHOQZ87kY2omOo/R8ay3t7fKBhy5Q1Kn9ZbN493fB/
pb/02hbQRQyHJKGJtBHheZGVOTBBEUkX+awCv9TmYoYqeZ2GghmK/HQSvX9sfBjb
uuIjln4LCxLekC0TzzFecXfdy8e29TF8oSSSW3ftI6DfIxXM8X4uu2TMVtD30MHs
c2w09ADhb6Cfut1qPki4ncdvVzT5Xy20bIMkNBH3pjAqXpQQXJu5F0WkXxCvDkLU
sb/S0nssb6dXEbtDE35ScvQuejZUba51mR2rZwOp8l+PJrXzGqFKZa7zRVrYNtWl
dE66tUNTJ5b7cvofJ5pFoGFpwAcpAZlJT7Yhl+/meZ6/f+AStUXPa0MJe7e7+GCj
GJG6qmVRKZ6Cmxgfk+9H/cBNiW3ZVKFfQRk8hdbmeL+J8lt1Qh02dUdhuKAv/sAl
OGahNN0CGOfLrFwwOg0AVeHmvf+SgEZWxzSKZdoPZ9OprM689peQv+zmYUNIxh7+
3IBSOKiazmIuKxRT0x1j2wuxqviRaB0gDjOMMX1GtvdwXEssx9fgk9xzRB7BcTLa
Ggb6qkLXLXwjhATk6JDe0LkXp+l2vYcHitoY6UY3fXvPtqKsUvK5VycKWwSQGWX6
1AjdZ6jp00VYuEG2QOkluuHdapeaDnyrRJO52BLMrhicGwi/Tiu4Ux4OPirzHsmD
908QdAhBf2jeML4BaFdZbA1hrJSlWt5i9gmVgy6NOPpO6MgcXYMQHpY1tzf3UtEZ
QFa9UKikyn7th24EIQ/N9FDB9J5sS5xijPZPYA1y7Xc4MyoUc/jf8qS1eLTYDjkt
zcPGO/KqgDg6K2GwgRVvyHUQOStQ9iaRQQDAtUfGVNSgC7UjqT902ruoLRJxapFx
l9ox3DYN0z9Y/XCNX/b8J/uHNQhqyTdKYvmja2BHzi2bnguz8uRW87fDjuWe0xdB
4si4riTWy+UcXnbCpAWY5ZJJ1CF1wgSP03itwaMeVogOVKSnZsWPmW+qn7psN8zW
F9zCDg/Y8whRUyFrZ8J1Gimkg5pot0mTfFTQho1mX+x3gE7ArX+cyanZOk68HJbe
yKTf1jjfMiSg05S4Bihl3l2Ssw67vZUFxG/DJVnslTEcLBq8+0WsBNHEraG1Ft+b
cmC4tSpZImJb5gG8wZYPgBj5XxAlgMoq4Zi0fmdgXOvj0ZgnGeqkH7IiKXSPum+i
3FbCkv2TdW+7CSQDrZMq/81ynbEXN223mdeIPcbXJYYss0JeU5LN/WQ7mpjgj5rL
wLypFvBfVN4CYiTXb0xLEvWOkJwe+Pm9sZ92NfQxTtUfxbbijsFXDcBdapdCBmCK
ByiQUCVZonF7dq6bZI/ajmEkX6aFdUzXPrrRlZPbCvm7ZLzcWYJqrPK20aFLnacw
PAhP3mXIfrS58o8uwldqpVXEDYJ6Qn3Z70gVwCKd67Trp0/kngWRRbBMM9W7krQA
uGkxTT71K2hUOhtoHu7c6+ugHyDE6LfZ0CRtAX89BdGWRljLrfdhrSVlmbWMVjQw
D/GtuqWTOd4gZOjqSCPxqVW0bMsRQn9dN8IEtGGNXJydtN2Q3JyB2MYtdoEm6SwO
r5Wk3HXzeJrIMaL/6JDlWEb7JGygjVlVldYWNH/d6iF9uF0NqzsszVo54fzLeRGG
no4LgoHMyka9kCN+j0YJweqka2jFJ/P8IcdjNhayv78/7PXnw4bGEr1RxoLbvpuP
iTnfGj7h7KHCm/quMJXJewbuY1LfZA0KuyWIcwcKEyLTpl1iZLyGMMqNq/SRFRU0
hS58oY3N63kiv6FiGXPqtiOkJOLB8Wq7og2jFB0trr8g689nJTAx5Qlyx968HjXv
DsrYF9OwPuGQqNpA+kESTLuIYkXCxj0I4vvH9yfUYjOKV8rQEwBiqM2jARCQrFNk
OUgs1+on4msLC7K3G9PmLHQ/unLNiudXmgDwlwngRaXtPmJE/ggZmRtmQnZsDcDj
XjDkVxwiM/umNUp9GDMeByc6JGa3jUmfveDWQgGzxZ4p/cNoPH1F0wBSv9mqy/mv
BWytiBkHB1fOVyxwOFB9YkIYf7my9Ybm0IX320v6jxHiArsuLmCEuhARHympYQNm
0kr4Isi5KRLJXlm9R5TGOIhk/XrbtQZHAU3k7ZnO6arZjN9S+At0Mta2/Cxdcxq2
9/Zh5cFYJC9efMEiLTfXRc+oTXVcv2Z8xk3W4sZrAUdNNhiirU3t2Yn931V8G1Q/
cmH5COQ/GIvzU+IBjnNI20OTEJlE67nDcDyhzTqM/Sl9X7+dLDid6opfDboQv5mX
saju72twnvZENQUtixPOL4NePNggiUZ+FpmAe8K2puGuU6h8GnTGUEdeVXlXOXqi
BjlwwfgI9wNorjOq55u7PvqOvcySotR8rbEYxlePmuZiXMFuD7PHaYKIGRaxmY5y
/Cs1BrM3Ec74je8grIrlaKncNYf3W3T1sTOZrMZTqZ4zmfASAFH1eKbG5aoRnkYM
NhMyMx0njVf5Fd4+h4SiIY3cFWPyngVUMd/gjXO1IJ/yvW4nZ51TW/IAVjK/KqsN
zl2Rb/Nvme0aFoehgNS6+2QGmiBC5/hDH+QQi3GxEG6+A5MxC/RwdNI3uLAm+s17
ihoMdca7OqdPeqnp65PDcp0ap0wOCpoFJm3ecug5VA/SvfzN1fbhbRZEXWdn2FMq
4v6Iq0IuiH+B4MTAmcDsPFiDSa+VniccJepq0Qe8GWaeDnTkd+gh6HQuNOhCwpEJ
RtyIq7bjAY4V71/ehmhLvdaAOfDRMrHJAE05Plg4hVY4pcljBpPEfYSZaY3r2WrW
UKUnQIrmM3btGAkDxAXK/kCmYPOoTeRgOogZZBHy3GBOls5Ehmiq/1iWt7+OWfxH
baLfhB7sZSMwoxFoTOJRykTlCozFzZVeazPc0W34q62vicwBVA/eGQ3g9UKe1fI9
OszG8NHKKffbAdVTTf4XdLXFA6TJFhb+WP2Pcv8Qxiqtr62FK2j0vg0eTM08jjrF
xTTUdapHeoT/0FDCX4H41F9dEHqRTFJSg2Oi/Ye2PfxuzjExnsORAZjeTcF7f9eT
5aJVm+xaVAs5jab0E4/80qmh7n0hdKr1Ngq2C0qh/gDl1QcrJwR3ECCF1v2mqJdS
1PwA822ONcMzsP3FKoMbozJzzZKiwmDPSP3JsXFu7nmg8so4LxaZXPaJv9O/NhFI
DXuz8g6ib11kAbZcXOeO9C8DXosI86HLL6mHatuIetS5tEVHUlvNYPt/yszbv81p
1bli+OrPaXxKsdYyJ8Ensi3U7scn7m85vceHrpS6wQ94XeMe0LaJKspzVSt4Ox10
2d+pxL7exTREnhX9afUmmbOk/Ns6c2o03zaLTDAPwt5pM4hFB/MSIqWp7tv35ZuS
DlDFeLqiDRLj0qs1bI5MXCEMioyDzFWCLol6aMmUr8Tm114UlQ2jAqIP+/s8Ws2Y
FvPF3CDXAnf0uem+7SR6MSKSeDun2ayLG49PMTlkGA8Mz8z4Y3dKPMhUY+Zuhlkg
RkDjGyje50ECxDLP6B1LhujHO6imCipdbdOUr93w7VeBANqXpSroqdQW8N6+wSpe
6CJMCsgRGQYlv561PdXlB2t4LkQKXYmcvBgxk/XSbJSyKPxVwNdWAq7WQsfpjWda
nEjZg5LI50DaElNShB3w78xRN870oZd0lc971a9itC4se0MmFqWj6gwDGlwD1cg3
MtPpVqNDWEz6PE/iJFR8Z/QX09pxcERFt5z2HJ8prtDGNd/ceW53/XU1veJIRoKf
MUDAFklFuwChkijMMex5KIqS/azTGsPg/sfbZVT+x9Xmbugw90hFscZVRMCZFJvX
HktHYQ6G5Afmx1Y357KcYu2q4q81fSeWhuQg74OOmKhg0o3vv8/uhqpHH2y+rKZC
8hHQCBPWlRFhXLisamVAMs0Q4W5d/Ny65clehYv9cjfzrCkfXaHUIsreV19EHVGn
VroNnA/4ElgJAM+d3pogFxdIyP09r2OlcHQ2BVrl2GDtnxQNNLgDPZUDJBRTHbQo
1QK13NqXDqCV9dMW1Ja5KOWTgxQTv2BiKgGNPWQH0kHBCwld2AiLhUx9nLc2XB1e
aS8xp8wbSYxzfThJDL/PUx4kPsDSxHzAWqr3NkVTPONO9XX0aGGZ2J4JbvhIXMHs
bxFtEK9WLJQ2UXuQoHcbS3Iqz1kQ1cuQZE8o0p9M0Q51vBFDlxtAECqdyZg7Vsq+
i0CLEl4ftt58/42vlpwf0xV7RKr5wdhxFswC2WWYFqp/SpCFsv/WfifSk0HohInt
HZaEaV0Y60gKqhPZpz9laWq/i1KS8TXSdDk31zn7wj5Hey8nkBaSAAYq3d31k4dO
G3+PVaS4C73TCoGB9K2ubwnUr+nTv/Mfxkew21P5wh3gpCg3lH89mGWstncuz/Rv
lxR0VFeSjnX3wv+UZubdke8uMM5CKNLcXT/JExOgy2UyV+jvscVsqMWupw2+bUmI
WJXfasPtISFibsang9qZ1NBdkR/lOAx62sHc54+5zAD/KYhbsojK/tftFlyJNh3q
QEPjTpQJZGsFtlHpeJkZFzYBvREuKNS9c8O+4fYFszf6VP5NFcrhaxfRItzhrMso
YZs8v2TYlxHwgAhlS2s4IblxwTqgO3WjjO2fvC6Fsu1HApBeSU+IypgTvDy5FWR6
PZBxuNk9FS2AopiIIosYjYCSb0FYhxk29FNTWsktIIVRGO1lGfIehIwG0yKVX5ek
AzwNmtW8BWtl0FL4iInDQUPhPG3czqd2+IWi220TkZE/A8Gcrg0vn1qkMAhOkrrv
aViXl/DpPwpSvLoQMu3MEnpB6QeEoaEgXmWcnSR8dFM1ZwbwaT6chFD1P+QBKY6L
60Qw5rQAKdGqVSxm4F0BxPB+NViz7ZMArnD35wLn7M07onCU2uqn68CjVLIDtlUW
eBln5hua+FpXkQOZW3fj8hwKcHFudFDDJ9b1E1f9isvAvbPz3DSt60gEJczurluF
LSs2GLyPTrTh/ERsWCeYeZa0eq4iZf/WFCY8ztj1aGj91NtvoV74miIKTvQzSPug
ngo4TiBylOPCaA5PImwjHo9ApZazjn/IzxHL5urEgyrZQZxsGKyTgn0UYvHMxe8R
JLAwF1c4r0mKN7NVYnf5hWGaEipO2bMRrC7nHgrKkbA4r6/HFwNGl0r9+JI95kPS
2QGRbRhVTeoXaY3vcat9wD9uUbyls6KfoHTVm2XwxOchHL+qPBHh8TIxV933rkK/
Q3BevHLI9JQa+PGXFu9yJJ3vd6qbdor7ZKP2w2ll45+dWMPjtPJ/Cesjra2kpJIY
oryDZG1cWDhBmcUlmbI+K2n3ucXAeL19g8ylrkjmgtztU898brwm0D59sUgbwIq1
zyu2NFziQ7JWdmCC4UOr8hJhSMWDcnq6iofgdHtW8JIMcXKLomuha98RAO/Dxepx
QVLYT3nXjPuhyRt0cJ0CtMMBKvwr8qZW5Ub5AD72up0kgXNf68dyYnYufvMb+Kkq
2Juqpd/j1kLF9F6WgoM3GFGzSkQMcP9N6lpa3lw/lrYNZgNkWCw6TNrRXEMZsUZO
xFhCfgrZfiPJ6rKEbrr4nHLQcolaVD2aTNC/1SCwewNfVzA1m+qV0n+LLHBnLSP4
lhamtjnfaO94xHlQ95SzlaWnchItdQLBwQmI1JG+s0ahEeF1C3A0U1Yqec4ZOMES
EgafF8efkcfnhpciuNzCz4L69o01K3Po485x92KJvyhSucuc8gjQPCDeFx2gzHH9
/vuXYw0r1M4igLAfn0WI0YALcthDoffPrPMLNJgzbMLhWDGlO7RIgKn7dcCr0Fos
mVJXFmdqn+XvvG3wN30TE5LYqr6tnAU7oobHFCXPSEFKU5au8Qo5YHzdGXNTpJPF
+LDGACVwZnpYyEHdidMuPVlEOlF+NwSqXV5aKyvquRLPLYslfczZ24OLX4PAZMmj
8SnEncXyh/K/SgTKDPQdUizLTgbcu9Z6OsZjpQu365Via1SWiynUqt08Xt9PPDEc
keNx1UFXKKDVYbDyxayVSKQ0qW0bKutlCm3h2yg+n40KcTpFc4rYE7IdeeLVcWT3
xzx8wvkDR+LhmobYfj4IfGjC6S9/aYqqLHcKgQDwPTDQ8d87/BZA1Myvavkbf0xD
5HgnSwcjf8OBb79LBzFQV4GwKQuevHt4GqzaNKFN3jNBHeoO0Cow82nuh4hNOY2R
QSZtAtzMV3AnltjYIv5nyazDqBBMrQfZNRbZF5YpX9AqN/1h8U181NqtwT956c3R
D4QpuxU+lBsjk4zggysimcyHkmEtc63FQ68vAoX3xSgz4tcJq47Ug6D/EGRQ6Pxk
BWOesWg/Pz4rJyYTBKIsk4UDFMGuAo2QoeLyp81C0AoNtXcw/kvbCGUajlBcMbQ7
PXa3844rfPJayYuZ/YvzfaG9EjeCq4wrtbp5io4fNHsx7TwnzoBx1B6HEZRRxzNt
FnN3xmv46S7sJE8LRLqHXg1hJkd98nBA1MsFjg7hxZYkeJ8TB3VwCfwdPZt5bg6q
E4IiYYBdzjHP6wdvI9ELnkd/sUYzyC1ADpfI1m2DRdxqSLKB/1jUnFa0qJCU5N0+
qxfBBqUuLrs3z6uTNeiXdxpuWdqE8Ban3NP41HdLEtZA4T2mIv+hzSL7Yzkinoq8
bW+89LzfbJLXKI8I/JlQYn6+YxPQFFD+DkMb8Rba4hY2s4AWjKeVY/lHrT0QBoaf
Mr7ltMMcO/nFCOtEF0DCCXt3ZiN5LQesl3SaErUYtVgCkien4+cpju4O0c2H6oua
kJ6lqeD/YcGRsMS7rJEPR3Q9qjrjBwULGUSJqscZwPYDshBVbYFDB4NeVkNOoAhY
nRJzD9S/ScIrVwLcKcDieoe9jIa6Zf+gE13on1GKWOZ7RQIVOttnNQvgj3B3ZkNF
3CFhst3VjdxvFgbwdoKzDlUj0AvmpUpGEi/LYBrF4FCBW9HU+gEPneTHXzpzSMPk
erKnBhDixVaXJ/vETfcRVf9K8BhTSDN2g7eg0iBDBdkfpbDXEqsG4wSUHeidBeu9
WU8vkMDFFXQxs2tJ3S2/HjQLHWPfrZrrJKaUTZ198G0n5h9timqRTtt+bttmV9LP
tCbTqwP5qKkkO/THTKnKrfHN/XjVTsXq5Tyv0fYx2rO3FlaykxDiDZDXMgDN44NO
yMnvexRVekAZUtxaFzjLXQs5pC/2jY9G+b6DTVUUjov20B17juWphVPvBvcOn931
6sTDRUeJIyzcnwvXwWlJJIfsh0BM2V1qXkX25zADpzXjxmPsqP4JbrvhULSp83+1
Kqi2yviYp5NPGwO7CjoKMNlts8CtEI0hmVgHv3gzP7v5qhHOOujmY4xSwn6Bn2fP
qVSfTMQ6bAS/bePnZIST0J2EcuOaA3p97+HAlU8IFwUouzPWrXgx/nq0H3Vk8zxg
cLr8EMnTsOykmIgDENkTO0Y9OMBxriShMonKq38O5xtPjhwuYDZyb76swcsbjvZ7
cPsc/e8XvbDRWweUVNu4BpdO8CUbJSwfcm2cP7+qjanjbt8dE67z1y2kOl7Y+mwv
SldgetG2WfAlZmJnocTkfAdnlCRlz/Nsrserc8rsRY23Q5qrV/ns+ot+mxDZNYZu
88TLgI/DNjVBusI+FASUbJeW0XHxCsyC+wrn1MPlrwOlo+L9oC+IkxYHrHQLc1eI
CPlmPzo/6EqLllIQmmiTACRybgpbk2TWaOjhzP89Hm7i6wV/gILOKXUWCQo1EZTH
iV4ph24Ui+cNvLcJ+N3vfk+l0yB3WQN3ldelGYDwlvzVVfWMPMc/h71iPi7fYQsf
zOZCY+NeAP3nZ6Akw8xaj6mOwm95HsXKnAYegutTuzCbKQLmDgpHFj6mohKjObYh
qDwdGYh+l7zAyjsUT+jnUAUvwEwCkblGk3B0BpLS0pchVQT8OtcF4TlRyX7V2CWS
wJmUr+DCDkV5KB3WEnfiSP44p2D2Q5MLxBv/RasbvS+tAAIh5MFwnZoqn1hvteEz
kPsGylkYhN9Ib7YxrZ8nuePuP3YCXKDIEjsmURQBRyeqKSgTgXbvSpcHNMCzFW1h
KlAmEVP4KeGlwAhd51mecCzZZK9tzLYfU6nqagom+gTmPn3io+Yuz2A300HqdFVj
KUDb2TKlT9HAEpFuEFoQBYzROR+GBnePfAWBISuPERDqgjOS3xRgSMHwosgDW1i3
QEI1RPN+46IoM0/tBqeyGqHsVePRtOE/2qMzaws8FrcgjMj0Gnt7GfMGcDbOfBXB
YLUM4peNKJWLI+e1RdV6FKe5USKScMhPXRSqYqdDFXNe9jtCF2cWwyI3LtdaYBh1
mjv/2BC7zbBGS2uGN0kZb2kKNvABtDnEVDfX+hdo4BlITwFwkwLpwFFGGgTw9QEa
eJi/ywaZBWR/PkOtANdVp105BliqFra7yUH92kw2RpGufWaUaHEV6BXKERoKhQfD
qg+m33IA42nW1bYMWcwJqs7yx9ZeKUP1CE8S7mD0aH3/uutPyHsvomeSjLhrDrnz
6M+LyppAjTBo7WrEOe5YDg99Ls4l0wmDnMx61GbJDbpmb3bD5fOtTrR10y+DL+gu
P0fcXu8R/DPIXzRaxaSPKIZG2Q84zIa7hMfyC62DUlrmyjlxkq/QbMtnvo6PqbI2
6nwX+lDt+xhvAt2UVrI1IBjHsaVxxOY1/zjpRlzTJxQjsGankvcDMCw8rqB0n4In
dpIsyQsfqMZoKAVPsON3x1chk8xegKOPlSyABUn9EO9uUpmJ4CxxOHaLvzrnlX0a
DG5vMj3TStEtN/qBWe1M7UMd+4f+y6PiMftncgpHFjSFkxpuNv+LwtygWg6cnpJp
GTem9UG3CIq8k2059RXVzT7NlJtxyBlryC0jakdf+Y8Y7d/RT5yakeb24Qd9vprl
onliT62H48kmBEEdLxJ4uAuYyPF+ajvbz+7Z5rOy2pTczAa7pQa9jf4AtGv1aaHT
MvDSnUGCE4Gd/RXyvN7sj6rLQ2Cq1LYVICpnHNNM+aZP4lcxmFqX+kk7gj2RUxfI
Kpdfli4Tvci1SxCsj9mb0Na78UlELcHM8arNdSWQMpe9wjJAe73/F1dftZ+gBmUp
/rd/VYXfFmBivQuGpPUi2WVbVwTc3BthkkGockm4Kiak3W/qi0iA2b2pbjvzodt8
N6eAinP73RStZ9muL6Gz8N7Xu6wTtFTs6qdagOPIGP4+jM1WrGi/Ns88OLudlbz4
sMjxiDhaZQm2rhD3PPhJ/7OOuhGkrUPzAOWF54eAgFT2wyNPHixQykc50ae7xOqG
LI+23FU0M1djvy4u8qn68V0Zqh4FHrF/5kELBr5uAr1kA/7sGqz8ZAFdWs64IVFN
xtWmIpMbvSP4TwFcTBrCDe/avKxwaFkaWzbXfEp3pF7FhH9UdNV5jLcmSDg/JPQj
jcStD21+QvFx58brS6sqN4SAcHjE28iOgtUxJsYdmmBr2JQB0AEBBCpype2OIGrF
fMMWPp66+CVAQ7lcT5AgAZZ+7H6XrMb1hWwyS0FS9idaccLKDwkoXhE8sFINtB9Q
WZ0BwJw3s2F+uB5sq1H1seWPFgMHgyu/r2gqTHMs4TK3hMtZL6GaOscZkHposwwH
plVBzqvNAbl4m/YT3NF8zzzj/g/tdInk7WZyjKZEubffoxad0RuQM7gmpUzPZk3I
AGgU5q3ZbVxB7JYqMw72ANG0EzGr9Ztk5WV/dOARE777hsPtOEuSmkyt52tnps33
p8I1enC/XZyHwwatsbwZ/+zHXX1FdaCFyr9xmFYSs3FbtcuTBXtI49wK3i7A/Pys
J9ZaQ04JjhJjlTD949zyjzy40uiWubAbkjUuvn1hSFUPFbkIdnEJi4Fi29yZYnBR
+WdffwDfxLeQS8szzGlmC+mRS8pgN3A6u1LQlKma2sL9WSvGkmNb5HmGKLqj05pX
tjmHQjHzLv6zlXi4gvrzRAgDNEAnY0vPHlTno46mPd2oo9HTNxyHiHicp4UKLwLZ
C9jHxOWwLHBEi7yRawjdgQduGFYQ2VtVZL3OlWxe4+Tn4wjC5+8jTvapJ9t1SJhs
iywYbuCG/AcHyr0b7yujxs4uWmv/UVwgPtZCqftJxaPV+FkzG7Z6x3Y/4sfbyG7Y
EGmfgCPm0aAggYGwpDZPW9dVFDqfzqZoLuyz0r5S78ZUdpOxjEhs2kfW2AZXuzRH
zy1pzk+wDGNAazkL4nMt9w7Cp1BZ8Iz/imjTtwHHLKXq8S0bNOdp1EpxyJbZMWBg
/CJnbY+n36k92n3H1eSpkXpJ8V9lBKmm1xuXTEnfxJqnob/7IMBJCEkAu5diAMcR
OBZ/nACuenVWZKeWabxhKtuNS+CXM7oGNXUU+Vu2pfUAWn0lI7HzBV9Rsu6XROwH
FHs+QgQ4xVwnHElPKpgdwsDevMIjEmRZM3y4EjxWxU5LSXAhqCTr2wDY6boOK30X
JsvddkcJZZA2kTGrqPMystWZ9ynhpcmci34Vwg/hNCrwrYaNFJlzApMroJS6cdfS
i5BOX+ljBRXzxVormaqb/CUHJlNNLNb7zk4q3/8dyJ/QOMzZk0zNcIvnRG5jDnRA
XGbHHeeFq0C0SoO7lvw1vFgF3IWA4QpNlGTj9/OuoBTGieIpBfBqUEh67kM6TXQg
O3oUHba+azUewdRqF5tsNCOU6IurXqek9Bfk5zKJOFjTcc7FDwfHEq3i1vcIVLMd
L6Jt8o4ZTmCBxoLxYObQuC5o4aUL+WNr6oihXlR7MmYMS0DwsO2JGhBiV/kGciEO
vd5O+WqYOBeghtozkZhJ5zBFnamRvIs3BNGn+5atdKSgmqrRj7DFDFmJbxzpT0tN
FnMZUcB3wbxBTknozcYek2NLgzVfYUdy0dNfXiT/dHvDGyUOLn1E9A33KXHnwocb
Qxsg3qX+hTDbpW+dJKnjDgTPuA+INJXeomiKCN98XKXdWB7CwtZbmHmeBCEF29DR
S5RIIn1UEEEanvagDDdMV6H+W6vCU1qy8zW1LBPiqM2ETagQ+QCOA1FiIv4+60Bv
pDql4JkolW3ki5nCLIjIkyGdBAKQYSnVl4fsqpbod6H9Z6+1q4zAXotDohpmYWbP
1ZoWovMVeZptm/xNWi40lhONdOyyI97gCMS1PyVNoCpareibeEdb6zRYkzoGEziN
wiVHzyfcbxmE7Ej5mgTfnb0wtYh+Xgb/5fvu5m9Bmu7SwyZMSBoELA2zzgAzZXqa
qxVaFsRjk1/dA1ZTxwmnx1Bi8EYqgTVjLFbWjhf8oP/yEC8X6RMnUBuaLL+1Or5H
SRYulyO3xYo71rmIKLFmUxVqDr2z6EthSewYgj5HVMropTAjhgnPE+3OUzPNduh4
f77jeup8dSkfa+wY1v6tibOTBoQQBKmUzHGGBUAtYGSoz0XtYZaA9pGKmmoZ9R05
pxmkQioP7ZXbUXk21Nh415xNZBeEu+RbNPLhjtI2vc0vRSk8ievY9+pPCERYjRzN
+2YoTP4rypdNUB/yOW2M7j+BeW1AiVcRrEL44CXB6qm1FF98r5wIre/ysGTJ92CX
Kj/zuE5luGyB52K9y8QSWPHHe3rYuqzbNUPRHNH9heYJBQbga9WE6u1XV9KU6OvN
gR5v81imeIxxwZg6CqU5ki2QCqUVGsmOc4xvkokuu3XrM35m97pNGRDOylH8WdTn
Dp2uHq9k5RnJjtTJIwhlXNoVkYXZ1Wuc1lZ2ytp242ZrQB/8orq0j1LoDH4kxRt7
CLctf8OMqqocSYPrjNwbG0Xg6saW9jhWZ/u9vOnC+iedYqqIa/cDowYIb9AV7qae
pRYNEtbzpMx5931CZ8yeWPMTR86ynBw0vVGHZZiOpfnlBCFSo0QC9x2BD8F1kyV6
Udd6NcGwJIsf4PYiyX1HuQ4kPBv6+1skZwMtnG4Yuyy13IbD3Q6+IIvEEPUqm9as
8bkZOyRCP8nhCIIyPwUUAuL++fLXt7V4RRd4092rKryyOkRw9S6JfzeSE5MO1/Lc
NSN2QOy5eEOJX2LumwHJs+Nu8taCMMjcN2aYxH6Ydfgkx3mWMdD1BkzjIOpc6X31
NbpzptwV5KUotq4rm+fFlrG4b2M7S7V9qGrrNv/OSeiLYmQ50jLkFJZZx2EEaI7I
M1TtySXFiSiw7XL5C50z+fP+pK/0IWkMEc7BKGhVAH2arfcmcIM42AkJC/dA4k3P
U34Qc9Qa4a1+2rMCbt6j/XKo5qGoAKXmsPUrR/JogZ13UPhjOgetXTx2zRQ6YVtV
Ak+2BvUMTWkTgLcngPU1faU0l5B3/wpweXlioydF54UDF8Q911pXi9I62PLlP8ad
gpixEhm1I6g5CMQHt79lMyd9fHKwylg31IElrR+ln5DBe9r/guYZ4YZ0eVHy//o6
h1sjbP1Yh1SDVAdif2vIRoz2ZTnBjQYWugTA9iKNgxvBvB2Zjr7x3dHo1iG6XG5u
GEUc37JCNO2CBuTA4H3LGDdUxwEHNEhzawIICzSHTt3qvrw4nDgAxBNYXa/W21ec
pl9A0NlOwo62LgUjqA/eDHHjRCzjG395ToDCnYijotRtQZeEwlgd6zfZrgZYD2IW
9RSgfkOsVYDvdgen1QaztYhLQeNtGbg35WlPhVwpfceVqHV9CgAoiNXN8WVaUZwz
6MkO3bHghlOObGLT5/vQwihFR/8Z9W5d5LcoHLG3Hh53SIEMH9lwNXHCFpgjPYZh
fkKkUKrV7CSnGhV5Nli8oHIf5zBj6NIgMn1GbhPSX3GXTgTiGxrP8bWOFw+/q/h6
Vmd/XIdW1bpXFyoWvCpk1uWWVgWRz+i68OYFUKyjeMx4NeRH0v3zay7jJAOtTWRq
WJ1/BR1MhLivUOG1wN4b3cj98k8xu3jFVEOnMjcjL6iLzU5GQU1lLil9zV33JzGm
hrtK5Cl18UUl2paMV5ohFVoyZc21f/a/eBruJj4ZwHNg5qLkyeuAVW4DptN51NdP
C+WDWt4CwC4+wFcI8DYy5VUVluKrTMOfKuF65DxnM1u10YACIGYY/k6QY5F9yu4M
glXnwkBOZLT1JiKRQehQOV4rIhyvgEuwzNZ0DnCw0sCQxoqdRrlJsGVRcY1e1P4O
WVdRaVQ2ShfzDKWLC6ZwOoDMjcXH0QQhAeWFWKp2BE3DZVSkPCFjNuj2A3kBc50N
NAClc9b6avfWCzun45LUVvnyiWN6nhLNH6yv0fsQZzfFr+ACugMlfLCsAsxg3lsb
2d2ed0PbmNSEOmmVv3ktkT2EOc3IOkYXjtYxwzSS/fVPoOMz0lbE+NtuzIkoSUSr
p7lA9nXyndK8U1YdI7Tdvq8vY5nmu4X15jy1ztYU32dapwY8EEikqNrfLF493McD
3L5uaFajrXXtWZ9ANRkWu5AY9oPvaCioqraUFZ44AUvyYCCj7wxXd8BrhD8BpHV7
7fi4fzXoOgJXzg6DsmGdNaj+grL82SwuLE0UaMrKAaUAzMU7HIybWfdVn3EMEyPX
Y4huGZADqcqYhdCdQVT/iecy4PX/dmgBkU1O5TVZ4cChYP0BeYsWnFPVN1e5KpYO
Jd6yvp1fi6MlSuBwqi0j6u11/133te1u3jOWeWQppT4YsmOZE/EqN2i4wXlKmdJj
VtsfTFpn0lP+kcNFxvA7sLLoGfYS3wRPdGHMRO5dis4oX4vcBaLdkN0Ltz6akkZO
Rtl+Cf1yOHX+on5G/GetxZAzBtfRjDHlC5bLJXynygeDIYHICT54ujD+BDEuC9DF
DrvTS0DnvnZP+jyH56EQgZfKu48rUSHme2v/1aGFQNLcQDYzNBmsqMkCcE9EjJ+b
JtbpBKs9phGQnHRCnpZrwKS4gu7I8VaEMTz7ntgFi4P7F8PlYza54p051QEt6kRu
hH/LGeldwFHwLszxnfduXRZAh5hMheroELhscO+M9cOKauWt1E0i6XKirUuFRBuI
5mmngSNqaiBuj7x91BcWKxYM75DM1x7tcVOha4vsNqL+Qa+SPMV4WEFf0HYCSMU5
Gntd44OoIjZEfq3O0zGfe1Vr6sC8SIDQB7YzGSXm7a5o63qVKUjjquW14I00Gi/d
wAGKJADUe1jWT1EBiMSZNq+D5sRWr/9p6l27zLP+aLzPcsV5fZ9QIAqErz19Po0U
QABUI1N8zGYGeXZU4XKvCpP2evwdmM64MF8uGOcnxk73BaTjkQRmjW/O22w3tl6W
L76y4JfbFDHEjAjgqYhmTIMxYpoPnWej6al4fbvtKChHihTS5OX5GmTO1ysZ1Xn7
7/Cgzl7Gpy6fVTRYn3SWJhqarG20F4VbL9VqcUU53vqzQhSHMFsyPk3b7ys8plDH
ofrfNWE37+JJ4OLz77Kq4TD6ln0/mAdenvivM0VXeBsxoPeELJxGb1fYu16gmNeg
REuZV5iZSjkgWVZAko2DR23Y2ZrxtRCBIDuHJz+6qgKcilItslRu6Yg68ciyw1xm
U72HYQKyyE0nw7G777QJsFhR8ezE8LkVVTnvxqKIvqWQr+oL1XjY95yJqJh/1BL/
a8YxAtE4HjmMve62uBUa2JiL92y9yXJZhRC2HmYRULrEur1wUGXYaU/6/ys9ICO+
NvLxFGD1kEeB2XK8K3wpoHLpTn7cxk2ROe5Tg6SePj/5wIPWxeKv0IhVcf/IR1Lz
sMpRePHLAJXrDQrdfhsPMk0cDo0pW4nXHU3s+jK7nST7xh+gLSUJP32ua/1DrjWF
lywe0gXX1XALaKKcbtgtP1PzVWvRQO1nw/7/F51jM7nRKLQvDRanr6PqSycLCHFP
bY8XaXyqKMBL1HFhhctCr3aQike4xb9JBTsUoRMYerh8GnRHztCn5vdNkJOutr98
Jw8ArQ7SAjrZjQTZg6QayxISbRhT61951VX7StHOcWaRQJwwFdLDfmR+vAnXFQd8
SOvn5+HDfeji6TPedD0APELz3xPuyt5AG7IIAFD15leuENhS7Z/mcnH93Mvlkq53
ZUFZGexp0Qnp64XhCfMq+2NYvY55VwIV4Qe07rOrT+/egqEUoJwO7WKlLd8E7/MG
uF4h3dNZYbjMhCSF1jsSW81+Rcy0c1BTGDPgcHjCwaB99yaHeqjTffINk8eLl/xB
2StDdIDgwv85vdQEf7DGE1t8De6TPmwm6X1H82rcLUDILISlI7h/fVqTyOSRsM3U
WXmUUCnXjySGKoJ8zi1O0t0kcXgyQQnhJ8Pf4jxntq/gKU7weSRGlKqwxpZXzD0P
Yo2a8WME9e4UZ9+KJpdvC+ed+4tFu90ZdUkLBk/XRwViQhxQ8JZ6GGb4+CfvooVW
BBl3GuFOck1LrLqK9MbmCuMQUFHudAjNXE5uPXSg4pYs9P+LVg53st6IxAWIHVwG
cy2HnOZ3LpLpImR4k7EQegCL9HeE9jkNHelcOKaBWgovbQ5N+CD5zYHvZDxUnbtX
fKHffo1CdWb/AHprLCcz8oFZh+0pGsaB3uOkkD8f6RHTEzu4IePFdZ1Cxbk5/GXG
X8Ir0TFe8GDJjwKsL3ZRps0D4n2A8dmEBLtZNtzuVL4zMIWvHY6aant036A9OmXF
zbPNz856MfyjBXjfPSbKYBqkOIsbscCorDJ+KOY78Vkh++L6yB3e2/ONvmgFd+FN
PFuZFQARStk7Vw7cwTj3ZjTUH0jZKYmJMNTzjAIrbibIPYUwMqjasN815emFd2Dt
Q+a1ZqVQu6yt/Gg+GgJaoKpfieXXGtFrY3NeVFAMDLt13LPQwRvg65Uleh9b9Gn5
pApgH8kNpb2vK2KU7kz1gF7t/xo/aZBPSMys7mmZo7IcZqArd5xPb5GV4bTPF2FB
yanvR1RP3UjgsgSL65yOmOnLRXQFBOOnX73eGyRacv7VVW2yBfxFNCSkIpTEvXyQ
6mJfN1dblQZleH47UJminzxlcq1uMs8sqKWLlhip22xN4wma5xKHzeXKLI436h56
8a3wb9zg/YdpcYh0ZQD0L2pZG4qOoA+hRvCGkXCMPf5YeqjHwI1prsjqPJn3Hqyo
jFD8yHECBPug4sDelGUJZURs8/FiQnc/aMrS+kuo/3bDBk7TU6ovXY5zJ9o4QhmK
Vnxz02H73vWM+RyUH8QIOUb9mw3kYLEkVB2rnM+EGVrRxPys1lFoonG6qfydi04j
Z9lBp2duUgCeQRhcVTK2g1HC71iea1Hu2aRx8t/Z4J7P7Wc1axBMt0C0OkeoJ/6N
221k9bpZdxrr+tLicBN7n43EEzUOs1nJkq8ywcmPRPwa3jz20g/HfMlfo1fsDobf
lpNaPbaqnVK9GcR7sFtaiHlZjTeGYyiKJQNnymXszdDP8SDPFAojkbrYkS6kv7+X
RIPw80Uu9IXh/DcaOIRwDdtjTwOvN0dFQrnrpeFZWQF204krwpzN54OSZebdQa+f
DkbEfEq7H040BLNTWlZneZir5xsgYrhWTPAzdT/xdWMt57cwluSnPKrl+yaMhClU
fyeZNfCzsO9hbDJyiAHjY0EA41lUObIG3aBr+UZ6moI4+v1Bnx/SCgTrFfllhFJz
9TfHr6nTRckP5f8CSa19HJ9qVwrTry/9gyN/PjLSWNLy2ixaAc8Yi12+CRSVWdT5
6lJVuH9GrS8fDFyTUPtXCfTt3vh8F6/t04HkPGFsYM6+9lzIdeCywCDV9IL/qWSk
iZKruL7goFE2ecIzvY5xSmXmv/AJPuxzSgRNm+O8ABIdIDOvduPIFF0gDTjKVC9v
84seRFXiF7AUShOFk5bLZKAvsdKiGKwAIolbup7UcrO5lTmP8OtFezNqGMdwyjqe
8LTPNRw3EjpU2ofwgbtNknTSh3b9feufEJCqZnueQYlAV1/3U4OHm4B7yUj7F8ct
1E1wxKJKW5kKehJF4rcXAPaJigkfIez3w+zESGAxNHhR2cIWZAng88Bu59dIqrPd
0rboC+KknNhe/oX7MrzYuBS48c3NOloI126rS/NsNgXbofMg8Wa9SNqt1TKDw927
Bj+rDAbtW6mMWARS2oqi9xJ/dV3ZHst1AZzADnrInkC2KPpkiPF7ELCqmnA5MdRm
oP9A10/Rt5wBq8rEX12m6HqdgMqFOVs3PK9z2XH1W0335Tw2jCZqXk0aR+vNu8De
1TZSXPNPKUuklTXekEqOIaaec9eqT2TtspMS+a9aBPOeo0cbJfJg8Hr9FzOoOttU
Let6NNIdWyLQvB/qitFI5Es0lOfnEN1YqyvkhiEVN+fuiwhvPuOlD1Bb5XvPC5ZQ
C1iDzIOQZuaJF9nVhQMoG6o/mlZkRSyVh/lWNb04GayNm8msDUQHbA/AxCOAG661
Xywh+OHxJlVt008dqfOtb+j49iP1dlTwcjoU8IZeAlUBg4QBP2Gz+csmOTejCuEy
wE9mIcr52VqjId6Vf5DlxDORDtoX/kpZFdhYOlfmJbYcycFO5DH61+rDRuTXnWiL
RzBHC269BM2R0nfUcj6U0xZtcfD6LcduFnPDvA0U/tVB2pcJXfe8foGDZu0hzWWq
YCIjGUmGzUqNjPoVFF/BDAb7DpYKoX2veFhNCqgnUdwDE94JXLPbHgOz1qV4Uuly
8cywfwG5B5/aBMxT0vcD7U8VtqH88W59TRljl+PDql6SyNZwx2HJSZajc7uaid7a
Q88TdtfVG5xv89PMJT9hwW2arR1iVBVzLlkRKA/Ep427wgnpT7bOnrWbRsE89NRa
8pQbF80ZNFCkJ73AN55GxXQU7BtFxBHc/kQZiRe26fF7fRWBhTk54szHgrvXp56e
WLB20EH1qd2ziATg97TmYK5uYnc+DMi7MgGgfeGXSD3XPfXIMywpMHHWDd1G3UWI
Rb1Rnm1iirvNRD4OVbolUtjoxvIc/aZUh60siTlPzGpRzuOfY0BuXCT2W2k8qk2a
qY3UswRcnFTKUTHRBtqSrDEBSPuzJNGe+ewdp6lZLFsyHfH+pzaaCDjGwAFRpWdC
7qorlwSI3UDr/OrvteMEh6zxEYdsBvEUFoZ/gyTtACP/CUjZ2cxYza9q+OJu1A7h
+ytv7QQK082n9CsPnpBP4DJrpLZLGY4J2I8A67vAOFihsZl3MPSf2Dlg+WjApFvJ
6Zkq6Q2XdwdTD+wwVH2RSG9Emburg/BB8HJRO9JIDtZg6mSFrAY6fGT3dv2khiJS
J+b0zlhMIJdRoQ2n3tkpYB7jmO+1zYdGV+CGhZ4GUhaIYf8Nu7jAQLrlOWp+Ox9Y
0sy4X/mUEvzoxDaYkUu75FQhlwNXPh6Pfqtw/wxSDjrCj4mdZZHmntHcoNNOEr+V
MFE166UCHG7Oq+O7tyaPE+k4BfFSP5xHpbZEZVGGUoDtxLOeQX8DGS9QkEgEr8yz
7HxMLqRbcWsKz12iJRDtOJb2n7KcLSeB5sU7l/U5yZFCsSL3E3ndz4DuWEmaz30V
BGk9Q0FlV7Ovn0FijY/GIhVrTry57rHMqlkBZPoa23CrjE3wDThdTL7KA2VrSoAn
cA4KCBSGrCrINlPdvrIVJCTuI8Wm5nK+MXb1d6gugwdu3Hl3NZMVUI+Z6RwJ1Y1Y
QhzhRFAUMgYNoeStpIL2fTDSCK1Ew3wVNVM/y/nyWzZEzzwQ4g8mJe+H7aV782/N
IogH7i+DjyIn+iHgZbCAMLmvNe4nKm70pZU7TeJSdI0rN2nTP+zu8Ikpc/xKmI87
Ve3IUyQM2Be6356gzw6zTbbLUFhewkoSnS0tEURnLMzVQ2G/yETwkFQn88farMB6
3aIxQ4PE1+BoFlljf+GB8HJuJbgyXjvffmuEbaE1GwITAXqa5xEEtS/8nI1upiHu
jh/fdmZzKjkdPuNVV6WmiV/lW1dhlZKEFpsNFsg1B59dpSGjzU0aiD+NFmpW46mf
zebvVVd8cblTSbG2CW576CfDq8MmVK9+GdLwtOdET6WLmiWQPDMon/9ILaxzgq0Z
QaG2mVfU5neiayhI4sh/3D5+/MO6CtRY+SlVjK3vHt/C1BODYBEQ8jd/8HyI0lKY
MbtiWJPe4x3XG0WVcyGrWO6DkuY6Gm+xRFMYrzYjA3XKaEGUqaaNIhuyRQi2G2sA
YhQYmOcN92SGZsFY1TuvyEOLGIHLhQ9SzOeX8HYbB9V/lyc7bMfsR5iefH8XIE+7
6w5IcIsENw5zXUcF8cw47LelxPx/S7u8qAuT6NpVGl03nJITE+gWeIz35pg1H/09
8TS/wf2iKZ0n0PCVUzhiKjqjT5Un0ZYyMC29REWFPvhUIGSgB6EwF/Nl6fTRw5ua
hjLdKwtcreAT2H1HcE+IwZg30CBJcSdx3oCq7PwAtNdYOrz7h39sQSqZh69ugUIv
c9sVz51XjDhGgv4i6hFMpzagxOaiXE3tT9aE8+TX+DtGRrIwtBbpvKQEA7glBH+T
q55EtKoeTq334Zs1HfqwNmvq5ErnNKLpGAp900TOoqIud6u1qleKixdfS8I/+Pya
nxoI6432qM3OeQQ1oHy/q75M41POd4Vbk4jMwTCLsdnZeW2F+Nr2/4858gMZlY3i
eoePaVBo/cg3Re7Tx1jSK38ABrnLGl6BBvtUbsrjFVtfOtsiAIsExxohOfNs+drB
2IjEZprJeanCO96xsKJi2w6+SPgMeY7Yu+xMM7sENoRptidv9/19nHogDfdWNWYJ
Nw5hWWsVMDqpp0Uzxs6wB4JQXcund7zRxKGFVE0wJeh866t0QhW7yG0balZfmbNi
bfIvdu4IqCPacdQgRpCD94lMoNUVSeCoMSnjcbXpLrQ7XA15HxKH6Smr5VNfemu9
gVddwSBacWR4gP4zA+EujGxJmc8MAyZijFQH3h+mKj7uFotvQJyBZV2W0otL11nF
6XAquDFxCMqxI5YumifWMasPxbgAobjEvnehhW0fcGtZCs+O3bFU+emNBvUVq6kE
1JyO/9XfKQFYwNMsDHqCWnMWwAk66Cr+bsOFpH9XBFm7VXEEDkPHc5aF0MAeGbiL
M0yw/a31nQEMdo91ntziOX4eZ3iD3eLuVX1SEM5SRsSB8c06OZV39zK3sMXZFvM7
kbmZ1LJXtWQ+KBg3OoxeRekkZTf3/rDNb5XJkssie7JiY+Ny4hvSUtPMDA3K0FhO
mwGEgqSaAcWaV1sLc8bhOozJugzNQQXoL9O3ZQBLhIhSmoVtlngYgmmQUe/DxF3m
QXL/LLqHZzbhTy5E72ZD74q7jx0F/jNlLBp26mbpcLomvexp6j6G8Sr9K0CXJ6Gq
dcF/63BjZCCL2zi8Uqli1LcHKCmnnk2H4cL5u2MLFFAMaIhrVd0wGf/WP/i9aX7+
r8PQkfqic+YCXuNRybFTL89SmfLpVy9Xa04FG2fH4ItVpNtAI0STYR7XCFWYlzST
3fnYBmNMPCX8YNp8+/mG0QngB9HcgoYaZhbGAnQ4r8YgiNRiib+0qF03u4ziBILr
ac/TXDwgtoVuki1RyJz3ivCF+NWyR4tfvFVuLkl1zBm2uNBJNpY5uUXs1XQZ9WgJ
O1hPbWsFuN/dyIxwCwMHPFWtiVxE79rKSsG0E+9gbMu2u01JKyO6fdO/yHvgVmrq
9BGeOfYe9NAKjeKBoLGbx2NSWFlCOKKxvYx4kXSgpE6yw70sWjD+T2hRpJ/rPtRv
SCLu+BGVeO56af2KlrVY26tF6PFKToPUj71iwbAy41JoKYQGjrm+9ImKh2Qmg+LJ
w0iRQElD6Fwtg+Bmen9X9xyAFU58YZBtqrNNl8cHrUxQWDosg+rdBlRoIs08t8yu
mCg8XcpQSLKEoq4LIgSwmU9HqZpl9eUhFFTzxywFmeP+IpalN0uZlyTMvUrUFJvL
CTZN99meRo+ixkPDwthSF3yWFVoyQ5qi1+7Hww2HO9uuTKGgfC2JQWyZhjuRkn01
RtdPeKPfxPUnujU6coUiRejkpULQFeFk1jelBMmvcG75pVBSF1ceqD+mT+6cqJvV
81I1zYAUiM3MJ1gsuN5HUhaHLhf+10zj2OLgwO7Gcs4RCoMBg1u7nica1tjL4JQN
6qseObEpMD2r6lFVc77XchduNfjuMxH9UJ4goTI1gjhlm7RfeYlUPHZ2N1kWfjwp
FyZq2nE6UNEw+Pw388ePBkopTJPFCtMbSf+tlrz9Dsqu1F6nZ6nmpg3fHqqO8CGg
TVhsmexpALuvN3Zt6Eoc0zTfgNMnUCulrZFVQU+rVNIAX/hA/5qS96USuunWhfrE
oBcEOiCt/LZwWKqe8iRDpwEtxp1gpUYsYGhr1t8+x500nKytSYk69nfgTj4MAodT
hCQS4XZUElD8p9OXBcOtOzhHHemsQRjSf0QSQ894T5+EL4kWpz6zXo1BOAS4DI9R
kKVWh0e8lgJBxvKRWGd0FD9HV9tl3ZWMQ1T3RVgjhZj8gBuWRLHoprthCR9+qD41
oxUkqW/CeSkH8+5HSIxJcGv1wyc+xEbVa9soS19uxWDocv/Pt9JhMJ1nf5T8nv3b
I4YhA1ElhDvvpS92oHGymMfJZMTouK7jXqUqWvWgOubMb3h8LfqVjYS98qh/WAwL
ITCuShurmqt0SqaZcfgH5ILT4BCB09va+2iv4Btm6ZPuTOX1ohEA3dC9qZYRuvHu
BnKtyNcEb8HPQPlvmULD2s51B2EhsWQqcctyMlxUeWAWFnP6COrusiQZEn/fhhf5
yM14YozOXa1WoRmLI4YSwsjNWH7c5rQ2/tDzyIIqDQP11lnCXmGxMbwvrtNf1jsC
8Pf9ZXexhdaAPp7B6pdZavuEmuRuSYebEBWqP1X3N58RNSmhM+tFChrKSoXBdceA
53wnwtmrZg5oO80FQ2AhG/b5LbDSu58eCY6wschp1LWh9IOULekwCeuurv/HvjID
aYwd3cSGzqgD5jUdzdJQLMd71eoiAPhyae57jtu41dJDcddZw6GzovprCrdoI75n
wHdGscsd8Gc5/OOddITp8lMeW4E7UFEgomU10uq3E1t3/0wy/1M+/SBU3ORfbEkE
TYcE2nonKXzWkI4rffu2xgX7pNA3F2OzXCgcFb8EGjpV/IMHi0FdKT0O4+1sderD
LKhcxJ/rY+l+dYgD6pV9rSWl5jltkW9Hsb3/eEz5TcxtKNWEkBzBHaxx/JQPFTwX
pmrNM4z1tL8HTSKfCaLMObVmy8ESJAbN8hw45Gw53/FH65601B1R4QMczNbdLZBu
nciAZzADWkk4uCzuh/8huKs8EmiVyylUsAYKLCA10pBbDwUZjO+Hq84fXF8tbQBV
ND5emXWWtu+edbYYcMJ7fTRlgsAGsT+APw3rVcFLWmqbjsjcGb6MnyhXGxYwPLZy
h3iH5AjTL8xftZuq8KLhWUn2TpqEVs7EJ0Ktta3tDpMjTbO5sAL5OlONP9bZgRMp
IoFCJfPITkSSBQ7iltUN0xRoVk3/SnG6BVUsGqylU9EV6T4DitEjBCLdp5u36QWt
f+C729qgAoVr0w8bFKrVDQ7ZPdutaoOoFHXGlRArwl9HquMtIGU2+URPQkAbxURN
sLGYmjITz2uHH49a/2PeVa7i6y5bP6G6PYdM2cRRmkmomL/qTBsxkFY6QzEeTbW9
q/G3jc1yPQ9uSnUdQ5XbWEg94TIJvnYjnc/7ZK28otRcQAaqAMVaCgmv96+mlGb9
6GV55NrNuyUoOo+RNMtiMC5bpd0Y9xockdNi0Tp3JgQpViKMRVldd4PMIZbTpGoS
eozRfywWUX5g9Uodj9rwlTXYTzK+f8Oz97xVm90HmWNEbMlHQBV6egKy28D2/oTi
EgTYR8VtmRnMVvXYV5xCni/rZ4rovOGuHx26VLRjKvW/Ch5QQmFxJIlFMuNreSWn
ri/nWhCSa8U6wKEtL5y31av4uHzRe9u3NPkkO+p/EFIMm8n4pmxoz/swCOL0vh+W
BonfhoJPDnY70FYhVB72tdOi0C7NP4aBloAPAbfXfGIwSDhTId8I9uXHOOXn0OFC
rfuLnLmZe0ZQceSsHciAegR1moEOvhTDBj7VjnNUvnIJYM3lAGXfmg2riZZO85uQ
PAvkrJGDdgs40lAs/CocTvIMngil0LXc0l0vfWDm7YHh8YeLBIqVMKVUuyXZ9cR5
mihL1hqxhdEE0keZVTcv0x33bz9biHU2R7hN6qDYeDIvMSil9XFHizIURr+t9PEJ
xmdQ0edXLKSGyTsawCgb2+qXrRZTU0ipOcT1/z1XNyr3mjvJrIjD4J+5ucQZE4PE
i8JkN2U+W2B0khLuTuyDOA++eHRsQYO2A4+6cSo14b+u2U88XgdLrAKRWsN9e6HJ
znkGGQS6FfFOhZxouY4kcchB1/0XRQG9SKA+4OgENXOigYT4h5FwevZUOnByNXS3
B2DBwQ/qTZbQJV1/B2dVOyzPPrcYFOFYc6C2CETGqcijj5gyBYtlHrLd6Jv+Ze7Y
EnhmfJtGlIhJA/WINct8dSR0phyVWVBOoJIXVXHsIQrrW7tt7OE/Q/lZk5hacyGz
P+ECBlEWOm8qaV3Lsa/BZmRq+Eb6F7bC8pJe2FBdZ8zYXcJIiRqT0bKJLD07e3Ul
sV7Owt7nBmIFWckhWlhfghubpyAYw5UroNTD4NyTmenurc9MPxR1TzcLZyqILRJN
1XwepihC6W90SbrHhy0voPVGA++wUKW985ohCoA5OVLuYdsD2D2iV3v9WG39RmGa
JhrHu5iaHmwpvWQqQXV//fNkU1rTEviepjLlr8tKj343RLgXEHEiaFIjVrJwC+d+
AgtZGU1vz4uHrONy+pwy+QHWRsG5033uu9af6raqjwyxyLpURo8cX6qElPGZMsAi
WWwLTu2Ug+9ZbJMvUR/5uLw8/F34+csMloIW3Xeu7v8CeVk9d1lm5lLKeQpYPByZ
C8SXRIuwBNjQWFCNvZzzuvu1eNemBDp/VYO5HmGEIaNwEWSnLKRxVQltqsnaO9K0
fnWnNqi37WO7Dzi9Mq8TlWVVk/O3G0D0e87W4Fg13lTHXFne5LuI6tdo6m/xTLuY
BfQFQepn77FxI6ScCMQU2Oxt283CRPbjlqHer9x+DwApuuvaTBZ6nOm5VPNlan4u
ykdEhZ96bkcCn7BbncFIsy0IRgfXiY8dGUo7XSGMXgiKhHTrnfNws6oRV1prQqhh
shH/UhT3DIaKWHrE8SsqCboCXyLwVKoh3ZzhqM7WG3R+rv+rH/LzQeSA4HeLvZft
qDLS5a9iJWmTIE5wg/m5bs5AkNsYNkQhgeIrG7wV/uCMaUuRHMCdsu37kvkOBiNr
YwRBtmvRl3qfxQpz27lepDQH+NQA1q0Q5D31yC5VZI1jsun2OxQxYVVyxq0sm9Cx
T1DOHOXmYTRQWfG+e9D0pCgzi9Tz1Ob/Vk7iU53GSqaS8DcGU3id9NxNa8QdnQIt
rGQRZLNztHHYB6XgpCZj8Uo3vnnDkY4e8sf7yHS1+HFJGChOp+TNDAXDTW5Oryhr
VQAd+IUj3a/zmH0CRObFhKEowf+E+DuIDLRlCJb3gq9aEVhEUcFqxN3nQQrAjkTi
RxjJAvowlkw/F4yqvB2wnHJIhTtgdpYwLtpP03bE7WHJqo03nUKp4Sh1bbOhDRRq
3yEIXaGZ6EYMOtaTfqIu/ZAefZH+TIkuvXViT0Fmgz8y83Mu7pdwrh2QKeqkhwj2
qE59+lZ/ROo/fOl8236IqfIHN7i+GbpYy5WP7kLdnEz7kSIL3CE5rnjNNt10Xc+i
JFopR4d+toFRvXC1TZmYov/Z23muPA1VOorlAVZkO2sQpyNkY3x85Dje7Cu8R65Y
Oil77JvzO3bjuSRwuvSrfZpC/n1230tgxyRnnlIBgcab+M4uiTeCiuFSixtbfqby
0PGC73cwjG5ML6HwS/cMKEnSgVSQwHdFjPdr0mkwDvlDVMKP7H3m3NrUryScYh5x
oB6qF8KMV0QrXdJzhvZ892MqXsbTh2jjL7fBmrZqbJM7h9f2ROcFRmBnQhvOylbP
ourIZTTPTk2YWwNMNeO3mkSypnKmdwns46Reu3zN0LW2nvq2V07QqZ7Q7k/1Hv95
GtFj3ewi7BJnn3UMCklpm7U55PJ0oqzziYrIrTpZ9I/UicXT26AshWBc0yAt69Ks
e295ucjDMOF21xKa9H5gcUC2yAOaeSjFhI3X4fDHgufx9aZfh+AV8yP+qhQe/iQE
M1xbPgpj0WkZCJYJLnFVSB2KBeGOhU3jaQ0Q5kg61EaU/HPQkgF71vvGzBomC7f/
B7HTk+cXbqNnhNkcabFBMVwD/3SvBFBSRsqI7zyRdY/M4LhwGfkEb7Q39n8x10zw
Xx09tExo3qYz80DwBhRltotJTeY74KgqN1CT4Z5+x97N/UHKXQTb60ir1pODC2zv
PGYabYxZdtow0BzqWeqMNvp36NPwAGd14wR2/8sBruTht2FTmdLK5Vvlyxz6/oUn
KVEz108edin2RhX1AJvGtekjj5YE1ssWG2tjwsZnQDO/s9g2B29obb8PlTX9NE+2
uI0LMBuftc7Lx0idjnSnj4qX3U4GxJme8JeBlPHSyJeTcKcW2O8mrWBiEHeWsxPa
54+yRAFY7JvMLiKR2wo9rbFMsk9lkwziHJBXuZ/gb/y1QdXqGF45Y8itFrrPj8xu
1jEomJGHHDpuTaGKNC06lJSldFMHM+TXC0gwO6d+r43T7EY78ruaUyxjeUzZ1nYG
OH4OkJ3crPnaIOrSiTLw7Meh1haWx/VSygTgRmYQalZRIZcYgOVfVcB2yJXDertm
rCYTty6b1xSx7d39zM+DhJ+KUvaL8nN5E/B3mlx4y8i0qZmAO+AfhvJ3F+mkQFdE
keckCikssftFhkeZm+/Qw/xI26KZVKxcX3IBFTmwcItDs0Uxn6vvcH3bVRFREftQ
kItWUmMjBqzAPrYPTi/WdgrAV2CY5I2O3CXDKv6ZkE/+uTYNmmVNUXy1XMhKIJda
GqzfKedbpUcqpB33szq1UD4vHvQDEk4h672wy/mlHTc5O7q71UPfWzjEjsk6Io3f
oIhaKwyGmwgLDV/Iz6H75CrxNVfJY0TQ+Prw4u8XA07Rpkp1FYfV15gGfWDmt9am
TshscIywrqEaG3gYVstwPl2qcpUDNSGkFkhPDviMCfJv/yaNVHDYk4lKF3xpspeo
qtlinbTJ/nN3/lFRTL0bDBtn62VtcpnMLm78F3Npljgm4wKuw7/tX4Retss+N3rY
FB0rKfzKCobDlV5XE2kZDg7gko/QLzSDlhG/oicmYzy6UPHiKwAj4l/RecsFwOBB
8IwuSRaXMwrftTzO0hm4CYe7pYtCBjn8QWIBMCbToZJZcGMa4rdqQGZsucBQ09sZ
sOSqG6qK648Yq1WBqT0pDQbotyu+YFMlGRR6Z86a2TVI6ScD4M4Hicn+UHvnPIJJ
LKQJ+vOyHvc5XP9F8EKEOj+MGWMYaoLAkHfEdSKdYCItTjzXf9SEjzjXME8GSl9T
bOIw9POIzzZpLV0BxnbhPm7yfZeD42KFLhm/hkZvahvrgfqtGL+oVpkbgXVuSuPC
zmLnvr9aCeXfDLseDkFnga0/cpn/5BnCKisTycXgmWoNAlT72plpE37jWHF/oKo/
nym9F2bS+0wDHXWMi4koeVih3i7+d5rZrEIQ+OajgqOtuZ3UURQoxyvkG6kmmWl5
2DnmdmZxRA0M35Od4dMUSzFVFqUuvvpMOQfun5VeEWF4rd4ZIueX/2J5Dbn8WktN
Lt8dR5nxp4zqqoTK22blePXVdfrFNiAExqKSwshwx9PASENfdU0kPIJgw79l03u2
9y2SlmTw9U//bTMTY2Z+gp72fruFFhMQ7UMVGY61RYExw1rT+Ye6hAiF7SUJDvag
ymoaWDK8EUy81CPApC93BqPJeOEIuwzcdbqn+9GEbsqqiy0yeeoM7T3+aQvDHd3Q
WqNIpEoaRqZfqqHeFzVLOSVUOpuWR0hp60NDndz7C7U8g11lh7EQZ4VJrPIg0NRF
CsF8gSl5oIlCRsPbTfPbxm4bC6RbcY7v0P2YYknAAA8dyTzJEIdDQt09LF8fnG/G
ilF5ogoDlAfAFd5zjVN9Ef2pYoGK6qs7eDyGpGSC8yKyvOVPs3gQ7rrznnwIM3mY
M3s5DebeKqq1mZKj66QRZgYaYTONQri2iMl/FCYJ2Qk4JuPFzbN03nj418mN4HIb
P0uyCqsMVstJwXMMMiwPMT/VI+xKKnT8q1Ey1e11GRYL5A5XCXamuX+AlAuh7K6T
HYNvWSHeH4qxjRsIb2wtKRhnEsPoeQnjHwu3VTbywTwdKtrpa+W9gYpxx1N5cxr7
s/og7B5q7YIgN7v1eGIEaVDH/GPmmMgwKcBf9TJUXNVZbBFgmraGquqtku4Ijde4
tBog/jwIGZgb1q0l7/tGc9YJDxMIHADl0+lfXtzQO88jvdFRSUC+fFSYLpIzVLFu
fWEy8ZZ+qgBS218QodR96JGu7CFmMqgQplVASzB2G5MjplOpbH087dWw38Y4DYud
C3i5/DovAZgV9NVRsEE9m0GV+FHHoH+S79Ivljl5K66uzw7iBpWABJU3/PpkcJBc
FtiBlWHW5Gp+pEvlNdUURQi9t1NWNMKia7h2Hf3geyJy56eqwUHQn+1CcHjanNYv
UHvm5W2yyiytDyyGwxZyRSxL56qyrUrfuDSO//G+v6iDyaHn+RK2PdD+i39vzyAp
ioy5mmPuc7nH0HHEjYVdXM9ijRMu70brTVON+DbW5vjMU/W3hSoz5yMuJPTpZxWM
FfLSco3fwvawr+xzXjAnBSLZddRLPG7nxIjd11kELgx7+aO0/1OYjygilZzx4eRr
deiniIjeeu9omPuvyjTe7r2xmDX1jR1CGUiRvwC0iPgCARhzxbWTiqiDDTn6sVFo
+6g2AuOthJppCK6RH2CcJUEYwCYgaQvUpwJiXRcxh+UNon43uS5OKMdYz8CA1gWR
EuwmZIDEkXe8aZEAx6tIZjYaOAtIXJYtUt2SmtZpxMJkKOiXpfh7Gw8aGhIS+MfW
7g7UP36otE/cTL3WPmnmqqoR8BOtKDrjHjco9FApUvzVjrQVoe5l3s4MOAE8wDM8
mM6kJBQy0nXzwevvG3WzESOZrPXY1D7PyiL04TLZyPzpc47njzejPbRNNtwzudzP
EIEmNE//ymBaLgf65jJXY7LKwi97E495PIwkmEvfXiB3HQjpA1fYD0JxC2+I5pCJ
JlAf2BFghxf8X0eIgQigV4oXG7daNizG15fBX3DtI4cxk5dfUF3oUDXHDJRg9TpZ
vfUXkd6T23doX9gspvyiZosviLY6F6e9QtSCqoxsCHY11f6sj3ijq3poqTkaprAj
BtbVfianDadvb625pUav8ZWRo2YDPQxu6wY/rxTkRWUpx/00WGnod96uAjoZRCLP
4hjDlQth80tl07jRwiMlJAEgDibX9DKEyj1dAi4FdWi0zuJYl+SexEtiVqAMNS/F
m3Gaec1rylEkpgni/KOcNJH84rNhnVBZgWUIen35BXD7XYhE9GiRPVNtBSGmQeWx
TCdYDgr80SNYmvUO3gdqLqOv6fbv3BNJJ+4ONOhUnKjulVJtRjVMfP8bMbY9eABb
yKuFUx8dCLL/XFVSubgDOtCOicvXPvMYumGDGmm/1yKT3Bms7fyrfX8vMTE7dqna
EvU0P0U0BJJLPGgF7RntGbT3DQ/0c0MMTAiwNnhe4VCKy2o7JDQqbhbqhAtsCnb9
nZrodY+52CnccXVP581pb+Z7TKGDLQIlmVrkeyf0g9NcvsVj6Ayti0hsIFIKdE3e
T94GV+PKdKMVzqXNqny2CNxY/eiBUPeGe5wwPGkKcCJezpJh8fIm5jUPhodmxpch
ZMoS/vzsZpuaAOr7uX859UlskQ1DZXqHNDSYgOz2hpTsRdWWVGmYJsMVzpoRBI4R
HaKQOWmIbtMPrIwzvibEaucdf/6inQ0YXnYRtQBQYL7vHQCiQqfD9hTo+Wt/Zcqs
I6kHSjRl9wJaz495+dshuI5g7QVj75eq2GnZIM6weAFl2Mwhn6vgFsWX6VUkkb2J
8RykU+0mQm0xOFr04EyYwFT8RgsikSw/QWopGrdkRiwKYbgc8SAo0Ym/HYwZKBxR
JJamaiZGp+dkzQOugoVva4HHzkywel8X+lFlSEuDdI5n3JhsXmPRvzBBrGQrtKhK
zRwoG4g+ce+n1NAz0smxBlM/GdNaKL4ZUl7iE4Yh4ERayOZbSNWn/TdLWwzyWgK2
iEYoXzQJKGhqJn9BmmyeSILGTChhLM6moHNuxS9Jshmox99a0nce1ASD9qxyXOdh
2OkkpkYNEc2s4FJUKmi2X9GBeeJXw0ZICzM0KGTWnBd5w/7v4Ucz1tCzIaUS90c8
usbhzxrfdbmVs8HNbpo+ifWSpRrp1Dj/ImwYSb6V+7dAB5dSMRNO2LuBwuf/zTtq
QBSmLBbEz04h670SdjiL1q+B9e1aS9CXY2IguALRW2i0HEb4jcDOhIQNOtu5jqXb
ZW1CZNilF2U/Bd90VCwzs0n34+CvMK1jfVsJyibk0/utaIVY3khB/l6wccjIz3ge
LbfQfXNm5VZE0Qx6PeWZG4SAt6uYsvOMGGbIo4qAwYXP1/0zt5ys06ePEMLH9ySr
2u/NBS0xFSS/Li/RWPlOs6KVgTDxSFj+UTNaAeAg624Ku04JJQAPjlHpNzClJDuD
4zwzGmcIYF+Fg48lViLXRIguw+S27I/XaHHILfTiD3YZfdU3MQAqmjmc81lBpvjx
etrOCCoYSiPJ/Emx9dwGv08gLmx9mlJPKYQDs92SWgU6y+bUxzcX+DavCDe/z8mY
qEQRgoLmUrNleGNgyY9wKSMuMC5YjJJjnudOBGPz2tunnFDCUDRC4PfmWIh/ek4Z
/iKwtIAT5C9FjHmO4UtVkK9sYakjNIp8QXsMUyPGadrAgO58rA+wfgoOcscfisPd
AqEuZHITaSkWMg9WBfQINrJLVdfIGD2/UsZtELTNQpPs7YEtUTEScHjexZSkODWR
9alOsL5+EgCDtUCMszygW/Qzf/wPlxCMQgPsfe1XyJmIY0ieCNMLNRN5c3SqDTeM
YvpOFj+IpZr4JAH5JTzfgyOwD3IwgHgCCnAOnjTYxnP7fNCN+YZENB589dyuN+Re
7X1+aZpw/7TH9r5AggH+RrETT2cGwqbrCmHWTpJmLQepE7fxj70Fm0/m87w0dEL0
vbSeMhRqTDrFkAzfdhdumoJOUtEOmQxFkssYx8OOMhDTvF3ILOgRDZ9KpgrToeTW
yV3w6ww2m2VCYL/Lp1UrPhub8QtxYHG1dOI5ZIMhRYGg0yzHghr8DyHS4qiu7LFV
NEzUtmRcHqrTbVa/C2N75wDteYF+1PwPCzHlWFSfN0ICBeb8st3aEUXi0a4YN6iK
IBi792ESVdoJ6aAJUlstYSGmYCFIKvz91SYhzQ26iqSQ4c8Bpqx8aBe+e8WxDAmX
TYWCVts3hOUJEEspzsLHgZ0qri54dcdu5O0beud6YCBIMYlFzWhEsJasmtLmIf2U
46LpXsLTXbUJ8/Z9NikDA7pcK9yiqa5Kw9i5T2FWhcNR2B1CLd/vQYZIZFo8JpNp
DPo1q01jXVs5VzBHMbxZKD01ST9kTZuSIOXgBcFWxfEcNqlVLDca6IewTkjm7P/G
kqs/ffsL1KzYrYc5xlAbpvLZxhwsc9+/TBw0k7dAbsSc+oFO/AYXac9MTM9ichXX
V21iUWxNx2I/BNa9YV5tTewTn6WtLfJY2Rw1CXEen2DjhB0RGQWR5sxqnzPPXY03
mY7eGWBtZtqWBBXuFMWVHUHC0TTTl8SopSEmfoyUtMigX3nj4iuZuA+/WXkCJCD/
sNR8EypTUl7BFYF7xAMyFOuiC7doS+xArYxOmYfCFDjEC8xuvrOb9R03JOLw0fRp
qrf8Dz3j1rgPuv01SDOs4/4NSwSfWVGouKy48Xd1ML0WxFC+Sd2/+8VOJts/o8b9
p2OM7JkTh7dUp/UUIwIyxvUHyHRquncdIJz7+2K2J5Gxan+t7Zd+i7+j8D3f8qSI
PjNNshramkwCTXmjPrb2vr7ur7o6A/A8SYuEI2jxIXgCdO+aLEjSC9X841mwiGYU
kk0YgGYPP/QiD6sl1IQDmVutu9NaMUqmhdYRQra6cwo3K842j5vtpDqTqFlzcFNy
K6zazLvwKwlh5+NSNhC3E3yeXWMlXTnO60HvoH1ZvEMT04AeRJ+yF4mEUcY+lMnh
r7eXU/shBmJNCMxAGubva/XsTHprvVr7A2dq706RvC2+/hBQocOPdSM8sMLXNrXD
zFdUSCsyAleZVlWTaMpwX9fZV9RTvHxbT/5EDeoxFnsUzThDwji8+mbXdhx3ku0R
ZUlDzDA1OaM458uCth0rXrf66qMVhGBnGSJtMxFryiu8NoBK5pPi2HFfmfExEqK8
UZ4zI8cQ7AP+kPQ+u5VVTmgKwbbAj9QM5mYrnFuAez6kuxiRjDZeENW0Y5ic2ODZ
je67wZjryUT9g7+RwEJBRya2UnUsQdw2wdXxz+X4cer2I+WoJzvpfqnz+66WNowT
vUcGcuzfYbbG3g9o4ObQ0C+JhYv+UdQ1aZhaGiB+skHHKPwHe0ZNQGCnrxcqDOKp
ZQyEcsRQ6hUZxBIhPlVz+jyGWjUn44IrK9NzMGj4wu1JNlyUPF59gRf2iXdRi/x4
Tl75Aqn6xF8EfSPRrNyrizHKgQTbzHjp6bksyHXpwgsJR9omHGBWKRWNDt9WOubn
6TzxL8K3P5xqSF7EdPTwzSWdZBp+GRJsU7ZHxTw/hxcD8vpZWoxbpMvZ6ClRSNSw
UNEhMXLdnObyt8wjqNtrsMbysK+Yy5BjGeiKu7GKAV9uTp8pglrDCB3n/wpuz9mD
ZjifVDBwTAAQ+ST/C8soUyhOuXe4y2tfX909A4/F4EUANeX4voM9GP1wjvCkQwyE
Oh9xfr/Ut9SgIE39/+xsuv/1e38ZXAE2cdt6w3iyaoY46H4Z/KujgEAQCtx8Mbyj
Uv1jSjbCBIJeM2OtDhYLUqgFaxoIYWKhl62qgJPo/AgTNPOT6fTQIkUnISEn9naH
YfSBqMV8TbXSFg/bDt0No3rbiC6EM2nDKdK9GaFclnNB99R369zrsytzSKG3Xmgq
l7xZr+kLLrDYOQguxnK1tvrrYYALIjI98hHY0zBI3FseNMMXufxqyDqLvCyV7AGo
jzDT7D0RD4YD89gtRy8ATFCrDVwZk7iKQTusXAZ8LJKe+wy2K5JkbKpY0c06F2Cj
AFDkeiX2JDLmaoFbanJ4s6Uwiaq3OqmWkKbkSejn3kToA/LqyFZZQ44Ss9t/K41h
OA78XYHGeqUoulEvzbStvRsJ3Sbw0nCXtbNGd9jX4KpLCSvOX9IT33433uU+PA+J
3B6AFj/cOsdJ0E9eFDTGeOKH4hg+LK517b04VvjgBAdtmsSimyDzoPdTOPTS8Qba
ahpx7UfQrMASpiBuHyw2ZnGSlR+VKbemlEmdNNTCPSo6rTBDDZvQ2+c1/lf5ppZ0
mG4IFVgofoJ2/vNJ8sPmQJXQKAagFCSYGBGUJFn3L+s0JobB8rhElbw/xXK9Q5PA
ZIkuLEG1dDJ5fMBut7ViO7GedkPpcGvCY0fOaoaLCJph5nfeXPKvY1JDExibE6rv
HZMDq/ptjVcDeFUFmgOviJc/4vvK+wI6KKC0xT16QmegaOYKO9mxocwtCaiCkzuW
RzKyYtSw0kHRSfczz+yh5eWMZa/dLdN8jAEE0Flz6DC18Oc5hmATVpFtWZ2QIrts
7viDMYEMI0IMF9RBU0um2jjWqzJYrZoy0V9D7VVf4ADajD4s2gUlP1VMfVn7ginE
VfcAbYVQMaxhlIPK15+tvPZ/YDYXrrPKSp//TUWfUR0754oo39KR7L4ldsFCeKsI
B8NJyWOmeU/oAaY7Px/BMNZqeKHxVwSaA1ZrqTnwlVoN4EuxNnLhbFTj460LcHJ+
ylSvJoywmBouxbnb6pSOsMlHoPo1/QfUzILtgEJ0wsbI9DjaLIzmSeRGpc1RiF5A
dR49d2UmV+0/eEqIvkAqa63AOWGtp8uPHh9RLxUrN/JrJ0h6PJvfvPujJGzDCt7c
NbsnXv0Ak9FQ4OjMKVhu4BiafE+o/ORDsQFeR3Dpu5BZFgE7AJ4LVHHnsiQtzfax
ujn3hogJ6TlNfOxQHi94/oC45G3QGXlFo7Ij9RwTd7nRejmChttrqxgq3W9Cpjse
Ridwp1iEsv6x+6xEBX3WgJ7Ql02B7nHKRYNiHIY4bqnCqmlDkenPiWM3zuVi9M6l
5UzNsI8KDYPpmFN16MmlOVbz2I6/HDueMla9/DnnH+QyhU43JESTSlCg4KsrbxDI
s5ymnUY3XzrX1d2tRPVok0woQoS1AtVPHAgEkVzDkaVuCUKdQUUuUH39JqFw+RjL
Xq9JdOuvXjQWGtOXIvMvwC9PGgICyiKaSUs7A9uEjaQ8UpomsnlQDuApQFJIF2hM
Lv86Q4wybz+es8Gmww92tYuv2Nf0lL+fEkII+hW3WhGxduEzvom43kjBZGFPb2b5
hkmdeTRl5G5FaTNDJeGYtJ5bpA5stnJXQHdCwU4xywluD0FH44UA+KNHvhExCXcu
2ftKUWv0ZXi5zeEb+gQhQW6+KZWpoTJiVqOL3v7W3mBxLtoLHUP/FykKmAeU+s2I
Ri7cxKxDoa+EjicgJxMBBD5ohUm1BL7VRwq9rhJBZoXwFEeZbLUk+KuVBbSsi4XH
kiOygqO5Y6tVh+tF2mLK/3jDIjr5gwnlUBEpkFDwj/0kQ7LZ1/TkL4znURZaClaf
+BinoO3t2Wu49r4OBbXOYeR9zYZwXVhtUyHNNw/dESe0ARg+Xdz1aB7w7pt5LC3X
WU3zQGKE5GsBFfcRccL9BikMtipkjO17fQ4dAdDQAgbGJBITstrmYx7rnXC00hMn
yXONxBmps5BwY+o0CIInSTmLt1jK7oXtfrbD46qQas8IyvcI1SokDLeDveq6OJcB
BKVzkgiyQTrHnMIi7u/sy46LzTnV0bFCUvyGYpHVel49DmNmihmhFeCABgdVHB3d
Zpf7hOfdhh5C1bipX4vId+MBwhHl+9iIjXg2+1WOI4T5/ckIkGLFG0b0lTJjQAOW
89n/MXbM+C4buMD2vHmrc0si4ZJHGYorda4e6pdTuS8PLWaGIF/NUxQxGTOyl7ji
kqztPMb1RGPncbJrEekitrSa2uUsqua0HS4QEbNAvRZs2tzYSY60h5JXx6q3e30h
xeSExBeseRr3a7R7obI3VdFUzok5X1N1vYaYiCR9zwSLfQDqkitsafQ9qT4dYk75
VUptd4h1oG/QCmRhUM38qJT41dSiEUvJbU7HtVd67MFuNulghYbos84IMf+qvJXX
4QFOub/xnAUVVkiDGPeK99iSu6a+sIvYpbnFCeDzNwnXJNITPdqHUEiZ/MlzKbeW
ZoXGTeH3Y3j8cyeXxRkOSegZVKYrahW5sZGiwP7EO54S9gdC/5cOBCHGVs266TSZ
ZxfCCp0I6BZNfeGh4xZkR4FumFJWqCMks6EWcMclOQfyEp9XpZYUjRoVtk7NMOuH
fYWxpkM4blYsnwl/ulcsTHf96CY0L2llIcBSU3DYYW8DsGMnZLbeVB1WIl8pifIj
6lK8ltaiSXSDewAAIbA59dnHoB8npoTzwKz/54YtEpUp++N5/bwdJRgg8OrcGtXI
vQfp2WEkm5Q/7BIRsw30QBkmNRTtNYeG3YWFmc+XnXgqw8fWgR+MfNzLJWiMuevr
HECrSTi7wr6UNHQVMZByvklQ2M702pZYGGIkt1f9Jhxnj7g69EfKjMmbpKEDN0E6
+YaRc1Mw1yyXlEpgf6RJPusTwAE/bno/khUBtTEwWZDdA3YyfYpJ9rndCpfOsxNJ
1rWj+qmbvXj/wxwOJY+i1YNZJiDrY1TjLW8eu0b6xBy1hoOENotC20MbE8lZOraH
tUoirwht5EBz1uFRMG1h5mQ0Rrt87967+F92QdWI1L1MWQV6Ujn+AQSK+ee41maX
LO5mI27LM0Fzf9inqZgRSCSgM/CxW9IsMKxsZW5zeazZVP3SQCUArf00FjzzhcbN
8Dq83VhwY2mMR7jVUd785unM3JpH2yrFsI+FZTAI7dfjjCUs/f9pX7aOyk3O2rOv
/H/IMbcbJKPkAaobVoWRiuTvwSgPlYU5FhYnx2x/08yZ1jT4tMvXk7ILjtNmtdYb
Vfo+qc3aHr5mhJDETlUyD8yh4kCXv8zLF7PkUPrqQDXQsuPZPnScgHRv5Fq2J2e+
L+4nJttvvZmvnHB9JZFCHcCpIfM6bFXl3CPBqqFuJTY4o4/Cfz50zx024QB4iSaR
YHQSt4fLpKjs9Rs3rja46kNNghaUCcrDLeeUmzsgtMtr5RuvYuXmelUtUo6X8aQO
BCwiXhCsTxA3MhcPC8ZGA4xl9ZjG0ZQaobzkY/pyTl/8LA/mbxL/fFScK0UV4xOE
3b+XJw7Mj8NUC3ynH1R55U3dLnVFE4TdcsRvg4dTryFbQ3GhhYTqTpFQdBspq6cL
fs5ecnBgl9h/8W4l6hrrL4s6CtQZhb9I70mnkzFhwzBxUMz47Yx4Tw1NFgHqsqMi
ZwrYVZlF23UWftDlXnCnjARmZxKcajl+rA6uCFA7kRAD1siICGxhkq6jlUCqBTGK
Qld62/pYyaYE6kr9cijmEV8ttIuBLl66yweA1xkY+/p2GHAf2QlzuxbvnY8N6Ll9
BZeKVjIwYXwReUlTcRmDLGamsTc9SVq/ELBxBAHaYdIH0Nw+Sm1VZxVzIKPZv8UN
Gz1NvPbJt1CPQPFqojszkQsJVG0SgeAmLKu110TYB+66EUzc0lWQttO7dcWLis0j
ksbHdNcAISvlsh14v3t+0FhcI83vBBhEORGTKha3BZauOiqTSQpE6wsuZ5+b072q
kFRD7LBqcc2LNLtoFHD1E+eH5J1SPRkAFRJXmSavLNiiA059t82S6BqnSV3qw5kb
n//SmkWUnEi/ku7fhLmrb5WAKzP8Rd8l1k93jY1RSgrggp72SV1ZOEpTcy18Ilgx
rLqCU4pm/vSMD87wP7b9mk8HKA77yBtnd+hQ25zoTENAdyL3HO7ENf+10LNQvCZE
hAUZOBw3CKE4fIAS0UUttftff2Uf67yvneZz0H99pNRkgDZrNnGGhaiTCDC3WzWY
vUL+x64cwJ4UiaaySKrRhRl20aBkOQpOUwLa9vKZTiIk3qOljboefxjSsO8te6LY
Vz0xbMv191pnSi5TUV34yNKFVvhs+XK1bgzUnvaN1Pzu/8NW8nm83Tb+NyTVgDiW
1suNUxSKiLL2cNwqOlARRrHaubwtj3lmYMdqxMpg2AxBUF3TxPB0zAJYE2UgaiNl
scgFJOR/zBTysBsgPYuRfkD01aD7aXitTeQsDim+LFzoKGzIRdrQmBuFAOQVz7pZ
gDEmpMPNlBigzcY0ZCAWhIXSNjCrib+o/LyQJm/EQG3uI4HyPg9/HnALExjkRJKK
9ZIAczV+Fs1zZUPf2bl5Ftnv0QOCj1W6GNAod6XxYHxuVV7LN4iENPJlL7ajDvvb
/eI5BcWX8yFHwwx2H09lTRcf7nE75WORWhYO6QERGI2JDUydo5SSEyut+O8PYAt1
5OWz4cD0OfrWsJvfbSDSklZMqxsXD1VJZ5hUFCjWKnXNCGF6+MCCUUjSRxzKqeeA
SLkvbzgXBT7Ry5eKjeI3RZYsQ4fHCp62m6kd+1+tssrOcY88F7WxGeRnF4FwpkAI
nwkHipGJ14H4mY7Rp/tbxhXzuWhht02m4CUi2fCaEoeE5KggMaEJw8kaB0NSV1j5
E7pLsvXz8/KTFmdPToUr+Py+gyJmwz0wRghSQfiQ87hU9x+oL214mQIsCQt4z88m
0ldhCuRVBo31aOdO4sgK/Dy4s87RHa3XTA8cNKuYCXfE+k5fD98qnRRYNvZx46LH
og9HQrJkZ8L/sixeGgLYblzjvIn/5dUBkwJWJmclGvuI28e76FXCxpd+5gp1lkSm
fNpPqe8OBezZ/1GDSTYJQBibB85QZEhvA4ST86403DOqNr15v9sY64rlOV9jMqRa
dY/Th6ZzWIpKST6zmx9MhAJLTTuVtAJdOER9+tQi3Rq92sEbKcvyHjntlEHfIAyG
xTgEUGtlitKJeTmYH9IqBpyj0bbkmihjXkvKaQ48YEOLlCOGtAJ0Q+xHI7B/KRv1
R1PLFu1bpL5Upvbs+eJjdz9y7xRdGItpiqWahx77ZvL3TUZuYzfZzdedlTd0EUDh
CBUWMVF147Fa9QsvV0hxwYNEPk5EqS8hZCwzdLN6ugM9NDwU26/QTN6yocMUKlGH
YVD5SyYVaI6neCDrSTE0FY3l8VQZ6H/Y+vojbSTFeGA5SoTrpS2nwrP7TXFl9faD
iMAuzD102ncu5pzIpKNIkpOHBbYQ+PwU5ZBBK8mqNwaRBvqt/w8lhs7dY4wFKzjE
5KNnArNK0PRFO/q2Uv5UrI29bT7GrBrk8hFK1Jfrp7nmbmOhs2xijZy2iJyxPLRc
5gGQkncecM0HdGN7jqiCl+ui5crQsULMn3dz/YX0/HPJ53IqEmcmuu+LiXMtSgdP
sjH8LmQS5AYfbIOpc6fs07cquI6OFccVGFREnx6wlXeJ9OI0pXE0p/go43hfjHQ1
9t3R1lFLs+OTYlBnDXmxA2YE0danHYw71PchFoQvDf/u50Uc9K6NgJupEKrPyI49
t2AJSZUBV2qIryOtt0DpZMmnpziLa5KkfdmBUnJYifcZfmG9oLQxm9qOTDCBfhzu
opLotrwmsjFuKCx6oQq69O6ACwR2a+irMBHLkHw4Z4+MDGcRSa0k1XETVqkreI2O
+ga5Di9xj0aiSkYlmq1DToRtlMHbBC1zT0mmCNhoS7qN8qJdfRRssd/LYfVg6yA0
MGnbkS/C7O0w18znArnInDO84PnmG0vtZ0crZ0KuRSuOF/sTnARHsqrx+tz8SKyJ
eV2T/vSDx4lZpb04ZbF2o6Cza8UPPvcrp6B+aln/vIh+FU/kfGLx5FcHOus+KgzW
rGdBJ6G1Ljewh+/npIwmmU6JK46LkI85Dv/7Xf8DGzHEk1z5vcHxIjUD0KYvhkwx
oyjI1in46dVKP85Jb6M7In8REWW1PPbFz6dafs3Q4uaiAcsDNu+EqFPp7wX9N1HB
GJchUDmgrsmXUDMybUEuoANB+4p6IYo7D9cPEwOW0WtzFBNqZWM8WQRl6c8cA65m
cwcZQismvhf+3IX9ajZ91+HMo487AT65fW803dN4Wii4FSVknpyOQmzwndKbiDWc
Ymu3IFkvn2giRp9uHqnI42DAi4psBUPzwCbq4eGLrhUjs4ri9mDrkmunIkI1y++y
0UHSc2onyyYsuub8w/l2CJavjaaMZjRC/s95epKGBPsNfy8G5Uqrue32d4ovbtkA
UscI9+8E5Y4y3KYybXifF7s4iK7Pbw6HIfrZoC1hxDnoMw9OfgbxwJGGVtcuw7Gb
I091ba+psklSrlaUY1e0oQYbsjQXbgGe7VYro7QRA5zpmfEvbGpUPJ1iOqF1hlbL
rpieNtzBgjvKs9fjgZl6Tk0h86xGZTHl/zhFxrk0kTSuZVBOpt0SNN+OidePMb/i
jfK17JM+IGJmeyHR0aPzdU89t+SawB/j5TSeV94GWVxZaxf1WBqXctWCsglxzU7L
NhISr5j9eAMK4L0Nrm0N2Jsiw3cqv4cNkit9KAzEsUJIfuwzqiY6+gJXlqk27hYn
YbCBrMuYSlJl4M4geZKASugx9qJG2ET30tfxcAR8J7CXlo3DpnyoQnJdnc1Z3jLw
ofGJcw6GhERqywUrdU32ZMti28uxk4/2Z3L+KI7eTMVdyioEOtnyxBNup5Wv/EuS
SpwQln/tI9kSIS/QoTYiROB00SEyz9deeKKm/IeXAb7X4bjd4GoP+cnQ3Vk32wu2
yYFGZxoM9h4rK+G5SrQFbv4W6kup5GF2ewRxNMHH1Y1aG/nv1ovKYv9UNHyNJ3Bf
ZMFQ5hHhQYp/rr/a9R9tlQao8mTc9R9Y8BBUioyaKRrl8bEVI9IQjX8ssm7JTrd9
pGqyDLlEEKFvcmP5f2xSMQWVSXs5qLbBx9Qc4AAMH0VD+SYO9JXQhyp2rtNEJVyK
CTYYmxzDH2RyPfwC0V/w7YtuZNl5bfdaA5WsfMxUPivUuSB9ctE3cGjkn5G+wQ8Z
5N09eI/lgQSpKmff9DitAvJva0vRRm9iecJX2q/1uMPuDMPoTZuXsC2O2hFr2fky
toxMYDkEbnh6nO67B3uAXeuCxvTNL2yvQSdIXtvtG27uJ7LC7LRgJdwYPRyyJBZ4
cw60TzevhBRzoVra1oHxcj00GPcP1kbkG98z/a5fqdN6MM929qhsL+24HjawNLnu
uLRV3sszyRVuHQLnV6bhTJzIwNKJallSg1qFkiOPCWg3BGJe8BXdcu/yowMLmQiG
Ir0Wx1IHpTp49YQkV93XcBoQR5SbnHk/3Pv2GwY5tsmAPraI18q1R5FMAAYNpKT0
sUhCmaSwaMLD/DfpK9HseynAJIFZhqDCk3Tn9Hy1ijp+UzPkBK/oVEQcioaJA3EJ
du7Azi/dwkMxdJpe92szQiXl2PPEwudZ6rz/O3RjLh9JhQuFOJVBBQ9VgPlreaWx
q12gWdPknuMbqvglg9vnsBKjKSF/UQ4bpyDZnqCAnWTiUYFDyv5RMBk8QAHGbc0v
QbhVs/Wh4FJFapo5LdXwp5a476iPeOQv236Xo8arKbrrrbAxnR+zzCBaDeU9tWtJ
1oitH6jOTAZfFUYKUnAwG1JKQ9EYHNVXThkMpN0zZnrpC49TuHDSHwtnzEETuuRW
UW1dj59NBEWJ3ee36GEQx67t9cKnAwYsuIX8yrxioyWu3MglVKygRell+td5754X
i25WduPflq3Oa9VcIFCkDinDO9YX5fPXC7lC20Vs03tT/e4t3WxqEjp/qEzMBqRZ
IZIjECr+EahLNMPtS4kqZB2s5Yt6xyZnzU7gNqi96OQdgOjl17hPf5GTLclkXLIF
9A5Mc6xHS5n+RKOFMNaegKjee0L+sUMPnZMc5oZ0LXqrZhy3rOzdqHzRFzwdyMo6
5NIRXIbuTDKU2vZ5c8F66bIrLNGWppT/QPTCOlxtNR4klpRazSIcibvG8EO2p1nU
7S+bbIBPN9YCKl6HDirr1JyqMrDvtrwseBGh1+xVgUfHXX3y+bB/ksmpNT8CSEKA
cJSNnpIlo6MrC+DcWFi/2HQEXCkXim1ew11Ul8cP/UuUBFMcc5WaD2aJY4Hyqel2
G3B8+5rl6TStuCcea5BXU6QjgW0gqlu4q7ORuqX2MWu2QvxQCr+2kgugLMKhuT5L
RphdkIShANGqmFOrJrmT5191qd2tLqOuAvIL7+nj+g5uK5nrXFZ0Eo3bbZRkiiiT
0FdVkGwu9lvdekOIEWOSwwCBU9Zv6A0JHJ9ta5I7Kmy7aDcMLQrlK83yC4tn8/VF
s7a2dxXG2w2rLPnEvTCd12lfioSG/xUCKfyBvht5UUZsim9gb/VjBN6ZSjZtloVe
K84VP6nDhNHjfgaTPDFI+uHwMdJn4wQ+YqkW5EypBeSXPwtn6eiCeWpuI7G+csAU
8pw3jUstwBWmhpVlvOI+6i0T8mA7A+r2txpvYLC8zLWT+O5R5xDEYgqfJ3FxsV7M
QN9/VALJwX7B0ryWyZN/wvE6xDZwrE2dI74aM/4Zp5xSvdadi4wSOG4UMzTxBTS9
RCR7r9mC7P4hKnyHOetSb2n5Id7Tjm8FwCLFpjZTxylcCz/DPRuA9R2OjlMBqmlk
6nobtjo95XS117xeA7hHp0gT8IxzWZI1561IXUAyzpgGG2fQ+cf+gUp0ramlxnVJ
I5bZZ6EBymI7RQN8VKke8vHChYg2GJrzu56B3dXNF0fNwTGBrWFYmb+pf0WMtxYo
zB9/VI+itxozJi6gSs6KbSq0r3BOSSipYDOVSJ33v7O/XXJO639aAdKzICMyBPA+
XuvzWxySdqAAuEnmyvXokf99e990zWkIUi+99fCFbND/NMMRsVUocAkpQb5rEr0G
DT8uavTGZPDwqlm0vrzHjibWkFQWq90CGkVC4kH3VDeBVLoXFnEzEu/TBmDoE81O
2AMXSIz3eBKpSPYEJr2loM/qjTDjMR7GbmDQkmgeb1WcCgxVkWXDBJDKWxuw36Q9
uwJXJU01uVGX1oc1VeJDPSrtDRETEt48A4VHBnHaPxqy9X6KhB8ycjTcUAfSNNk/
Vv11MSTCS13/LHk9b+iczdm1jga28QJD8qTszdqUwL/gkTeFLwabO7elYLve/IAQ
FPd44sUE+DrP2HpTOVb3A/RyZMGCz6ogg3B35dlhvVbwUcUCODZn6g/wA/sWhslq
ZRHv9mSZEcpB4aG7xQ/eOMI1gyMXwlC5T8rrsPNQsUOxE1TXKx0YauCxmx73Cc2i
16atxvNXiT2Llxn/mKtwVECTsAasc5HuWj8L10rTIo35inTEMsI088xU0E+uyfiU
4mN0xUjCE7p6i4eKIHa29ulB88szmNcgnUxQvcuKf7HiOFH7hqHXCAHqQJv6OVXb
k+42uCVD2f1YPs0x0FjGbF9tnODn8sU1r5+QPS6VmwUQj4F+T2PUo8F5JTIKZ4Vl
Qck+xOkvMTS42tvfMRPBjd5X9/+aI3wZ+SDRHn3jA7tpVTJr6Mb/aqIhvbNzHrBN
mrXe35DN6MBLaICfTZsbjaAlNOIME0w/fZphBkLKRE1LzorCtkRdOXFPGeAU7j3k
vbV69evLhbSRcmk1U1hDfVayBgJqeKiCsjCIcILAr3slIDfUIwoDMVqU1kiuejvQ
e/b1uB/Dm6oYvx20leBc76JsLBCfJeTgyW7W/fHFvWVoVN4p1+iRNvboq4EMw3Pz
AX6lvIE2D+ZdjEd8AaVEz8BgrMzSyQ1jBj7MegfcZ6uMAHbPz2dKweWQFixd2I5b
lgmhW2gwwTCX8aTFS3PQZN2EgGNBg+mtXKVuMp2VQRB6VMfjwx3tD4ApBUo/kEZL
Zle4UbHU409IHKELXjb+jHNfhOnw7jrpREuRehww7UcsZJhdltMSMtxD607/imUU
golw7i7bPUHWIk8wXsP2TuPKIT3Ai9xcTNXn7t4YuPugs4eldunXOciPWoef3WJe
RlK4IOrVUGMD6h2P2+cwTkK3YNL7ACSBsFlWi/DSkLg+srBxLrG40pFVdjylvJSx
Dq0QP7olGFjT7mq+gU7VM+e2eMn3D0qafZI9JVLeBCac9fDuQ5cwlY4EahKW08xP
pfam6zHLj74ivR8dK3eAkikivIVt7Uam1Iz7tTyHt32DNXtY6CiGiTIQbrqtRqOH
qra9Brf7POEOMa9GbSF4kfpgty8hmvuP1sxaeKCE3wokc+Xv3FeiEWVEiQVkF7lb
tjYxHxwtYrKlzrL29n3pyBxgyQZ8MEVMyqiS8c4RPFUYftIBL+6KbXSlguirJcDy
ca1x4SolD7mOBXD3UjdVfmdApcgKnRyIVQNr0sbe8nd5Y2HU1ytU2jE5impSNHWY
bj2759JUlpIgDSKmdkRVe5cNSc+gvshv2ee3WeOrPSwGzCajgDPnI8NWtheKfUsW
nyrfGaedxsqus45gN8otMo3E6VwiLPFeT5NYUGHaorKr4tZM/TObEbfk5tCbJRSX
A0Q+QM2WmQnULmgE45v3GPRKEVapiCqBYjPhuu+bljfbTayjIL4tZoSm8sHi6Cwa
RRtLBaiqRmmxKDbC1PV42OaHuud++/Jvi0iWlusGYaENiZA7ms49i5esBWhXX2d8
+Ky94YvB/yaJE4ASQUEIy3JM2FlbyoxbIdarNGYnsMm4ph/z2noWcwEjI6tvv1if
RbDbg9bbPrNO+XgZplJK7NMglFkVd9xOj55zmiHjo+29gX1iAktqdPFFZeU299ov
KD2/JfH5ebPbuvIdQlktW53MKi+6tUy0tU4p6RlaqxjOJgiqu19utTizz7PKFBDI
erA3+CP8LeW5PYuS6GwMKrs9dybPyCkh/S9cWL9Dwb0uUlBH+b0lHqPTNRyJAGAb
/yLARlWHZIy/TmiNSgoJecHpJ0mNBygEZI+e85ATGXoARNi5KRWhime/2mHBy1c8
kJF08CuBAZKVjkAmIZ/+PHECfSABMJyOm/z25HVT3gkj9i//BgKyxJHIEEoIZk55
/hhOevoJsExpOnwg3liu2Vrl/QHE/IEeCM1frdg5SAIihnECt0cQV41sSF14mHDL
1adRrTDfikqqwoTQcoySoqgard93aRDnZhNhq2eNHZgfju2K2G+1/0jepwtMZfnM
t1dL3WUKJ/rTVPa9Wf6DftGm8WA8Nme/ZpnQYMCDQa1HmwiTARdkLUyiTSW/onqb
0WRUPneB2UhUiUePf8OIXVXmZSyNt3NbFuIZph40MbJjj8aDVunJHCv9hqHKQ+pX
OiFQo1R7ue4KIjEf7gZK4i6Ysyjm6z1ORV477vxTUoqc4tMkG1jvHTI9pLFY9Klo
ncbOzxIESSbBg8H7NXaksk4VJKQlFasnAjifcXWcKIlE22IY41SCAKyrC9vaTF9i
2TuJvwPAh16Bgc4I/NlTTv8unl9kOqf5bXblpJrz9AD9FnCRsHR+dV1itt3Y5JO7
NW73Wzq/E8OKZtBohj+ukXCmjdMgcFUUTBG6PdiUCGNZMqqIRXeY0PdI5l3tSUXJ
JZSKC3g0g45IhRDMR874kP8k+EO9PXYBDlHGDFh2K9iOOtTnp9uM1/pgflPIpYp8
tVB4XSF1XSp2oiHOo4ERwYDhZCkr61BtoaWzwYtG8Yw25N6O8NB3div8tCLuCwIB
MuxpdWXJscL+cn4p/nsctJLXxbuKoWmQW5K2mwA3RFE6rjT98l8C8NE6odIaSGVP
U53GIczWN9eYLiLAFcR4HWj+Nv4tWZpTVqDlfq6IOpYIXgkADOC708oVoPazjrLa
1dSslShtAJEUuSKCQfRBOdz0XPvt4+/zTirJTxRUW2K3XkW73+/A9K2bFcZecA7l
XZmOISUTVq2/+Gp7kipfWrJDxzUK8tTUHeM7TsZ6GjKNXJrs6bMKZpA2fCRUmkY5
rDLqSFp9q26/b8mJtqvsDy6gTNJPw3D55MrPMVueGsCj6rVlfnIsPI3pXRUqGsnf
EINGWhCnLLs2mtOZsmLe4VtXOKlTjHueu8+9+S1biE8NO/7nfBDgo69bM6vyXzut
t/7X2K15o4B1VllCoLnufGwyWU1yTi48cjihc5VAV2DsZJz7ijYsRuUIlseBxl4h
alNXGtjJz15BMGXj1/QoG2fNvfMUzRCoTZNaquJ2Ipm7vRBWEb//dv1UZclFdg6k
2EEzIfHRei1g7OwIB/fSTUtK0L9LzCABofOMLdDxJ5B7zClCLOvITI6YtD191Ygu
REX+CL7EQAUIZfylKnEgdP+oni3WAiO2/FwEiXwTZAkxFkV7Hq4q+h1QBPfHf4SC
sqQjVEywePevWwQbtjayzRUbJEoBVCsYWTIc/YbHFuIKmrjWpL1R4Ld4+AwlDHkP
66/TAtsXwxbZNTfWSP1j0GPR4u1ySoUODhQNq3qEdLNJ5fA0aYtTjA9Uu6FGiqBq
OQ4FVm4OtKyYZQiRXBWk+E8cHu8tT0sO1D0vnAnrlYRzrZCFV+bHPs90FM3/b0oN
iRtgNs9rov3785hbw/pOHgvu8XtrsNDxJpv1xRnv61pkoPIyO7nnLvn7GMKUcaMe
wkhMc9o87iKgnthCd323PThHc39Ml7x5s/OdRxs1x50jc2VD+a4czLxbMDiNPzHW
ynFjmsr5rx8YMX3RICXeJrR5tNplKMnlrPtoD6cfhrBHRSD5R5Wy/iLP469Tcnzj
gR30HOJltivlsjDcoOdNLzmrwnfo5VrcVMj194srULmVyR03gtksKN5rW21CPEbc
JAX7mwrBQ51qnXjgmtvqr7L8RTkZrR1BzAGZQ0uO2M0tTMe8fmW7x7YuwUIuvOeP
LGnGs5uqUkfxFj3klCI287Brf/CalcdGRC1RAloHZKVORe4jOUsjTC3lI5mSE3Hv
D7tgjt4ttrDBSVTE0BwgWby6gltlyESSbObkH+jZcw6hCod1lk5lcc3cA3qZwlUT
IkuRuStocnot7NR4eJ62knlM5F/mZY5YGh9nYke2Siu28W36bdNnuC7pYa6Rl7Go
cAL2dCHkHeHQa+Kt4vrtKaNO2TNfxu9W90jKkLl9xVJvakHIGEUV1xWhyhufQzSB
58RC13aj3Zki4Tri3LmrRN0AKGyWGrUQXScrRkU8BUahdIHgg7mQ1hFbjOp3s6Df
WXXLED8O/8ZezPRK/AfW7/eTXfZEnZJZQ7u+Xav9wEcoTq/j1VFicpCvLEi4Q6vm
o+f8lpMphmk1/pTBXg7yJ4l7dZ2gCgH+2Yja9Qz9w30JS3OBfRDHNHViUmauLggT
4wiHUiiJ9tS2It3Rp/Uhf7UiK0+tZPO0PDoEQXReMsEXvnqQ3S+b7iSStivPNZHN
XE8FHs4bQeLEeiuxx6vvAgvuJLQa+3iQ1ehAtYA8DaOu/e2EflRXmms9DCv3tR8c
um6kTzqLh7gacyXNlYwtobDzEHc/Pe080H/wiZXr0Ce8gqVPrcSUoij1u3v+FZC0
Ghw4WVkjb1nUk6Ye12GqQHNY/sBY/L2YDn820xzyB9yPa1r0eBH/WZdNaETxV2w8
tCbLeJEAFQFq31mtQ+vnjZ8IgIaHh5AcKmZ89YDZQZ8cEQWjXatWu+TGOhmuvbme
cYlavaiUoH2dOhudnbo4YOLja4aL2nBk854mYWXBl7IsdBjVlckrSk7XGk09Q6Ao
gcrYevqtYNjdmJI/kqCApLUoc6h3fb5HmD8dUuXrPJBYgmy7y0ETzshdVR4Bo97l
yBXoS4QCKbmUQNfdhlApD8lDVHwqACn7jgwSvBJ5nPQ7TRqmeD++vwJS+U9BJ7xb
rmrHBMBPynhW457pNlzJhezRl4xzowR+PFQbi2fQtY4dHVI1MF78cz/gYm+KywEz
FF1VNQBydDmSyG3W2VzlXJ0CYBLPq+2vhk8NIOv6uDkmo/Rcb2vl5k/e4yo6HP/9
pJjvzoQIQ+P/7prkHzbUxXyGGt9M2qoO241f2MbobOwi2xkwkwO2JODjrqfUtxwA
tqe6fwC27oFmeB42lZTJziZTPuWCm7Jf/Jxu+A6up798u688jW8XefcFfpnMt7J0
dE4otFnzYSgImoxn1ioUlcbkR2r0V9giPqoQ5dyL0bMtC09AtQjoOsueDy580Gqp
kwjPbcbAwOzc6WE1gggN39g5oA1d9w5+gRXZuOMKLG4gHoW1Nx3TUcCMpZN45s3d
o1+1WYB9YhhufQgAIYSU7wdkby3jtALL0Spxr9hf+0O6yAWu4d8TsgvgJnhYvLAu
/4yAK7z9BaPVDKrfK3mRIPjR3kZbgzHYqWgE8I5HY6CtUeN30pop5evjxRSAuiaT
dilrCGHtN79ETBSJfQ80YOyPVRfEBcTvY5ytFM6I74uPWPCujhSBYqeP8STKDNcM
PViDqPkxrLsaHEXv0E4sL7xcHfPaQOCCkqtb7KhWVXgRHTZxLMPlfGEd3lm29PqZ
QngwKcqolwta+Mp7hLGfEftCOabAzHFW4nGsEz/lbSHyBiXmckeuLmq3PmpmNpmC
0G8J1Ir+x5CKywQt6qQsPO6aKfHIeKTTr2nNmkB318Y4aCLK7H+tg6H4Slv618AQ
L/souO68pYT2afXQ6Kx3fXhyM62G+3EQOfWvtKtk7dh+nXMEyN8zM+AYwr7eVXck
W8GhIDLU+KKK0S8HlVgwhU7gv5uMhElO0kWh6X+AKTMLi50HQDAn5g2Jwg9gKF79
+fS7Ggk75Q4f5FUiqSc66p5YuG2mIlLL/68t0JSV8U/eOYC4dUqkq/0MPHwmGfnE
/8GdCjxPegCt/BIY+JbbeEX7a8l3bY76xqfs6CSMZiOgdMeI0t1zmpO+fISfR9JI
Mn+VNXizKUgXQ/O+GRJE3nh92jQ4/WYldfvzO5hFTYjbWgeAaovdRi1Clh+eIwYz
IU4cUkIHvuKFJslMwcBZCmqJDx2PnVUOXSSc1vGpt3RHYJ7lrZdT/sOcW/6fkha2
guCEicVCWT9J8RzXPT5QZmxYHc27L1ud4e3sI7Wuaxug9lJDj5PPTRNoqwYH4oet
gj1paIOw2z1lJRpzavaaSXICJfmTZnXXrHy0wjAPI5RyKNPFqWx3DUgh4t2PnbIy
MLh+J70LL6fmObIWmfP+fl5LJ7gkMc/Bp/86YhW8OPeltMkxWKDFpB/O1aO2MZpI
KdUktiYAhT3qV8+aX1AVedIbR1zUrbghR37ax5hytGbKXrTNvtAKCULKps6PDmMd
zcbUPG6ybx0uewMuXTX2Pn3sWVfux+1drbD7vDCRin9XcOg3vbuHUQ0LDZg5gmSb
jvmDnVciNjDZxNl8pxNaOKal2RL0URD03awAQjXyPr+BKmndEo+/W1GJsthCfAk2
75Me8cBoAD1OChEWuFyWmUVgh5E/ckiwHVRWmfwGGfE2+hw5W5SMj7/UQfObaWAW
y8PRq+VT1NgfhNBd2aiTe9JuzOhdHLf8tHUyDM8prISSYuoNVqZb8E5rYBoXLThZ
T4UfmtoXSojsPHWGnqE4ur/Hk/vjYVNJ9+GRtbe/BITVrPjkmvF+q7aqH1mDAV5r
a65LYa6ZBLGXPtp39uvKdLCcEHCFV/ijbAzWb/8t78lHSXW/GwvLQEdsZd1NjQMw
/1DmxEj8b4Rq0szXeZ+r0rdld86t633PbvC5V0dJLQIR8911gmlq0pwdZ4ToIjmR
dWOu0Qb1xexymv9TJ1UdewtF9iu4IIN4Y8CPsCtTMLVEHS7Nd2KxzNBgS0BxklHk
lNuqonsokR39NMrNji70vcjQUlWvFA83w6sxB5HFd+h4y7USxJxJAxBWYjs2Fafp
O9ds3z17bub7Je8xdjB1m2doSJlauCJYYTvct4T/eDuh8++FYW+3ZMlOp7hma/Ev
cge7sYtiJJ4wlNakGNtfnHuH752CpVBDHQi/BQh1ZC0Z+JAVIvrt0fp3kGr0SpLH
KQXBgADoT6ohJt7hgDNUN3e7TDSFAhsK2572j+gu9OrMlAp9uPJjpechSI+HdW+Y
MU2QbTkZn0pEV4s5Gw1HPIV2LMb8EL1xa8Wh1lTvC2v1CD6TgOF5Pegi1jSOmg4y
0C+r2MJruJCROLz8xDtJ9nZg+EAgyldYl/3je1TN2t/prEyzEG7kNvRtiP3SoCCh
JtUMxeI8ZGBC6BPy2US6BE3SgSyRqPyYd3J8Z3F+9N6RoNsbrrbtPHgbdFSR9IfT
wh3cbg+OwCKE9cwc3nHwluCX9ps4jXzQR8enkzjsR9L5lqC+3x4gHf3UEG9H0KFd
+xazC1wBPcuXhcW+hJhlD7PdH988FSCJwIyHka3T7ttFJA+ZjET1i82kO4iisKKV
deJ+Lg9Wll57foGaUKXxfQ6x5Zl0vz6l8E1n9YIPxFmO5wc6dg5inBeQlqUo4Eun
2iZb1Up8BDCvUFvDe4DqWs3YFdxiVn9Ab2eMWtctvMiKz5OuJVhvo/PmBABjBRFy
PcJEs8u0jgPypkDzlxE7PuqzxrTwdiEWpRDslW26eT1Ww2vikm25Np+7w6sZ4v++
5YtlTbnIKail7dZC6N/JgZDsLcUA9oAWcqYBXT/sWsSjAeNBRvLkJ6lMGqgvvJaA
1hzaayv03WcgBQErc0jkstH+zV5JGLZ2qMzyAHtVlLw6xMjvPkAfEzTkxQEZrWGt
7n4xRGXirH/Be8bDorhjk4KP8Z316TMFS2V1Iv5Z+26zOOKWHhLxQIU8GaQWfgil
XzoNs7/DybA4+Q3Go9oArYlvyzvjv9EeZIYq4d2NvXzP4FmP1+QUC2Ep7+7QrDPL
5nShXMoFfbz5IpjMgbvs7dMhNQDgznn+IYIMefriRYQZ2uujenTL5SvKbLGY3U+p
HOjITKA4r1wTYTVhpGtMrBW2cDXPTVGBINJukVKMRvDc3lsM8mgAPybh+hvTw+2g
GVMKJ3h8ZKSbTlJi/NukELOFhSqH1SUP8eBkbEbcVC8Jao72mJrw/LqwsthJsfg5
bbQQ2QNu+sCn7RsvZiepBN4R83Fu5Py0mKZWpUMEgwtt5dofL7E6aPRUhnq1/Fev
U5Ge2VJD++fwJ/NvOLiBC/bC1A+Y/nv4NFJBOzGzU6ysCiSHLM4qE2reNg0rRnYo
HmtiEjs/I8LS9nyMHFvugUkvVuxy23LNhdkFe43TrlZVVuFn0ir6NKErCoQsfS/T
kX0a05uw1hsbhUNvsOs24qJWY/aRa3DxIOkSlXaSJ7hynBZt6q7NGvkt8QUiPlWe
xQv1HqAj/EuiHVo4JSqEC0kWba0ximd9Ny6o31AwaYDMkiQYdSEQd8tCxiEVu5b3
BcsC4Jh+5Su98xoBPZt9alBy5iMgm7qPkEsG0MH3OaOIGlMWpj9SHswYg0sTQaEY
NYsjaaH0ScjQ8fhKWrbkhBI5xq8aYvsbOq6pw4SCmNCSaxx2yygvbtqpE7rRQQTO
Zs5bNcJcOU13bN7iGDhJsN03wkUA4tbbrpNek8dEbr/2VyEMG+8x3CAtk3nrZ1lJ
pqy5rkP3167Bvusz1T7HmawEX2E1vN6Ibp9iR+J+ucGm9sglo5lROd2xdrV1rumz
aOAzyrznVsL5fSAFjxhRqP7oT1UVQNNEosvKhNcKlt6P536VrAPdJn1m0skfwDyD
dyJHD01djZ2DPjT6GOIpvZhBCi6Y8ezdlshgoHGWKHqS8vnNCbwGMo5QolDLzqpe
Mc88Ql55kEwAAe/WrhJH8mGJbdl3FXq3QpVU7Rhp9qt6OYxhE22gi1QH6t8ZZkcN
YYCHLkJl/7GOuZ4ja2k/405cCaSadT9jM66BuHMg+ACcXkBWZ/Fp+8dRfeMhY1dG
SCi8erhmFpEGOi5x761Y74+xDi1WzMMBWZDzVx1CN0yg2gDfJcwKKygV2NRPM0DE
ixBO7aB+lmKjsXU+3Pzu347blbFV5sUY7oDC64BKRnAmnkwfeMtORAn+vdYVdc7h
ffVjeFHYno9nX5thBytdepOjenjh4HvfaFqmJ+6Wjip3aChRoqRDfqgzIcIPXTte
U2q8X2RrUzz0XBCzar0aGMyNZJ15PWAcFL42wVGrXv8OfIvvJDVYWVjtpfwhRt48
KVUAuSX57ZngE76SA+Cnz/Z8NbD0WWq1zgDTdJSQukmhKKZhEaOKaP1IZr+hXsNy
GqT5xsibrkkVzLlzlqXOMS5yCSxGiUcLR4AIGQ9mhlKtUZJlzRr3vUgaW/At8Syi
S5E2Fud1Zm+F4t1JUf4vyJseAJAIe4zb6wsNTcd1rXsBTunm7HxLkaXBrAgtiIqB
I+PA5ZH9lbZn7JfMTgyrqd6b8pJfLYt/jIN9CA6PQMOkPbw1p9v3KEpOgQwcJ+yE
yQTZOSuuMHGgVj1oPQ2eJlOe6fYDW6Q4yrnBv+P55e3N0FdR6COiGuG0iUOtrwwg
xR06Laqe6TNhchstgPqCjAZTFR7OKSfMvUQP32tq6fkGGeZVFjeDE0jZFMPCVe5k
bMB+ZIW8k5AYdks6UiwfWYL+lYF3N8F297q9fX8aTo/Dbk3t5iRADDOIoI/4ZHuN
RuMAlAlSWMGLs8i0SpidpMjD8gOEeSzPhT++Qj0NhRu6IhdG5YC+F+/xn6ypSVZd
nKemSGegQlPJGNPkLf7pnGDB8J20HTAygZOc3OgqAGlQSRk/rSnOgfpWonlpigrt
VauCK2Zn5+HRPMxYmpFBzYbpJ1CpwlA3PaFl0A4l541IxTxeJPdY46UCcchU0KzJ
sSYXR+S881pSLUAjWlZZ0vqWfOaIhIWvufTEyb8KWKAi6JQsNz4HTSnrw+4pReKc
oWnrAD8GbapdIRkSD45SlR66HZIcax8va3dqlmJo9GKWf/+MgIQugLXFj6wqYOI7
92LIMJ3h70wmj8/xlwJ1Uw/Y60CVplnt7q895zPDueB+mwoGur0/RByYclu5zqAN
V9CW9HeXFAB0ko1ZmyRe2fbODQ2W8Em/0wn3cc01tCii/kUhiUYzSVrDDsNZLScP
M+XCTuBw1AIr7M5Pl+kcNxhP0y5x2H22AWco5/KUN6VnezgeNrj8hjjVNFTh/zD4
p2jtKoZ3AIDelKbzsfiXW3og0fa7oels8Q6eBoo86trgSJrI0YjtgnHekJB42ruv
Y5Oj7JiRs2eFOINZgZsv7OWK0o4lY0oTNEm3Y42BYJG+jZo+jIPquCSZ9k/xSbYz
Bdfr9JRJ8dk0S5MhA/TUAZZDBQwT4eQVFkbgAZay7qY3+bW8+69FTVdJu9k/F8n6
eCWqm8w7lcniTe4HWWpOe/uXfj7QgBPV0+ogLSdmLH6d6cDG0Wuk2UmKogBXsjD4
ezpP5Q9uPTqyY0s4EPZCdpqwd4nRP745SePiiML8iwX9LEA8TMCuwuunZTlEbfUJ
ldn/S0vgFixPdb2zwgMEcHx0QyQeqmEq8grGTWcZTyMkWp4knit1Ekh4zxsvf9ly
TAJOTRWXLDkf+UdEYiadidlttm5nfmhYgCfoz4W+2Vy2su647IAarRsNLTXI/hir
xO/TyaD1+piC23G75+KGiVoz1Ci3Qs7BYbiY+78/IOruEwEOlrwItvpUxe2ilj69
D6e0VB6YcsqBbLYR6PawJ43BsqI0dl1RResqJ5T3lPvHbfEMIe4Se00mARR4bEgn
M2RAch4ooVJNyr/58L7yw0HtLU7OUGfgPI+OgblY7D7X3nGNwzjqfzxSCn2Aw9TD
amaULMwVYihU32VifC6f0MZkCp9XObIUT5CIYtQQe/QJ4GHNXJM82Z8Uc+tXRI1i
wQvDEwo+amge1owkD/sldTR7IT9ZCbvcAK7tD5OKjb+b6WRvGvIW6B6P4VcC1qj3
sApGm1pGFMTb06ny5IWhAADZFeE0sirnaEzgsJBwPwVf9z7wtpZkOMncCKHm2HVY
btZuQp5/8OkdzMv06bNZ+JudDtRfCRghbZzKRlNhQkV36vzIvSs0VAP56LySdpCw
HPj9y76p0BC21+j2U5mYwqKION5F6fZcduXvzzreu5xxHkzC3JERYQLRzQTM1aZ2
5gbd6+4hJtYx/39dVd0z88AEJ8E5onbGayfMWHWCPLqpJrcBtrOt8jwErfGyR2Wq
hAg8jliMWqpfvW91hCwz6kgrRIXtUWCuYEV1N20R/O2P1B7iGY+RzIEVwf0d4IVW
wsVATHeVQcDZnaF9Elsc5rs0X0OLQ+/AzP6/0Po+apIIk3Fdv4FeX/Y2H4gJidxm
k0GTBJ1V01ALvBRwdyWwBjNupjCDmxKfEjE41tPCZ+xka6n6DzBPN1Ja6tVimPJz
raDpokPzc+RocRflh/MzQGXEF/6COhyKXwNGMdUJ9m+eR/rTfDS0r/RC4AJ7hFsI
VMxPiVU64ipJkgGYnsZ8uX6/k/QTCjgGqtN8OOZKG/kV9mLPMU92o77rEAqBfjp2
6YockIjzjiao7IxbRZIZB2/nHnTWx6e2C0zqoUFMhkM2CHMveq2PSNV4fjQ+xdeB
metfodPUBfGktHqvKf80l9DMCjX13UJW1cUx38GzKJN/AxQfeNMQt/mq44RROSc1
OEiPkThew6SnShHvjEtliUlT3l0B2aB/AlLP2Zj0gnv/7lWnn9VF4h3okKnRLEVt
ta8b2/ZAKN7JJr4PNn1jwL39Et88zleXT77NY4L9APxWLhECi629uCPPXHEEeuEV
f6U8y5P3aePlodnIfxuIiIr0uUBF17DPTCQYwNy3PfqDHdq4hlK/Vbf1XqvyUwdu
zQkIHtgRA03SP7bQ5jGOn5bFvxzazwzJrw6Z++s0gTX1HYx6/zKUAsdtLnTNqS/+
/FkMrtiqGj15CtBZSU0RCB/gSM7PX0w+fBNz1c/VzagWKfFj8G1RTGG+eyoRcJEm
5Pb/GRMiGKKpY8wtuovpC4vjQ4j4d+ivEWbQ040WhPfP881I0fmdMnu8PpC3iVoG
5GLAa3xRMFKxChDQqZD1mVDquUVDQOuIAwVpYQ1pXhGFhzd/SN7SPTtMahdFgmDG
0fCoNr486fJot3DlsPYGJCXNgeFySBnlpaLtIo1YjoKx5O+p8MBXrKwFqq59Sy3H
kafRgDlL4tTufMuZXYZz76xcN+F9yHvtJ7B6ZWEpK7WNU9GNSv2Vflg5O+Gk52Vw
5fTrboNQB1N9ovrXnq+WOLfCHJmvcMdSCllQmUxFt4qTy0yLiyY3bdCkt6JOz3uB
1PFghKi7/QqV8KA0lMicrahYShbfxNklm4nYv7572rlzMq4F9k0/oAPUpv/NA+Yx
q0BpMIHl1NkJId2K1fNlopYNFn9dvjG3o6WJKyU6CdEozgfLa4n81KK8TYnesadk
3TP2lfNKX61EkWw+KAPpyK8cL/9wwXlqhgJiti+xzweKYF0yHMuo5ei/cyIsC9Gf
2FdvJ4ZRsG8CeJL/PMOCnXiprZ0GVrJBlTrB/JUfcAOfrdOfIqg1J8rakqcN5NmZ
SaQ41vsE0zt6rzBRCIiyUql0AsPNR3lMI+pCjxEFQmtmKUqVTWmzEzBWsLgMRLmU
EIyMzF/Ok6LRCBeSP97e0GnQ9w4ksd7FYSlAxeODALBelc1evvdN+A2CsxXLn5ks
WVSnZagTWrYXfqN/HoSzABQK9C9fD0B8FsZerG5QpucLufP8GedYZJYwUEy3DNxQ
OA3jPcYpWoaBIAh2RPoMVq4QSY1PG9FrwUeUP0yTldK0vMxbv/3CNi2e9w/dW/5i
4NzuSXALoVcvZ8UCQk57ujR4y21V5zzc0/p+TCEahQ4jQ2amKtyT4WNVJBdH/ncp
3otpO1YgzRXqckzf1quiD9kfy8bFR3TgkpfA/76fQuoJdr5i0GfAykOnu6TkvpgD
naw30mY5+X6g8qeNSgrVuEEcc3yfDnEJK8WvTaqqMO1xQAOEGsrgnV9fl+JJdAcs
jshMaL1vDm05YiKShiJp39KSLocYfYFB/tStBCdwErQfHitUXOtHUEK5BVa1AOhQ
GBzZuIbZi2LnklEhJ8FgGi4VpbEs+/Gm1ypWnmkYZf79KBDvuN8qImwm1nWIpmE5
tmIyGOISeeT0YcWWailfZD5sJ81wPxawayzwvNT3iGeIWRD2aXArkcRMO+wghbGM
AwnD7g9gkbQIoQ7zd7LbVazAalSVgfOqaPmvNHcWCSbi3BCgaSzlp38oFR1H5q15
W70MeNoERmv6RoebJiAlRx3+QjKgdAT9vOGc50t0cp5Lhltz0R5UOkt7OpecXkSc
JWMEu2C/p6LkuguPzwfUKes5Ik5evzvCSEpxeYRQfNyMcoBMAmHVA+52gJ8WGwiE
L+FOLImZzrdeJ5qRrAcglw7iTUbkeWF1E46D5PPbKJBhVTRdU5yGiMI4uSCq6JKu
i7n58WeBeoPsOKvgZyx/wDtszd9j6Md0+/AjiB5X4ftm69MRY2VuyD0CaAMMfjAG
XH7CvaVofaueCBC/iPWrRqVsA5nwt9k2I+86VD3rAXsCpngoIvVsyjI0/lK1+L35
sMxZWcHoUOvpwRE53kyZ6p2ie3rDVWRsIIPg1IDHjX6B9LY2VgfA7nJPwfnTzbmO
BoSt4ThSjVGLiNt8oH5CZdbWWbR+dOI/9NMnmFJw5FyutErDsQzhuU/5dhQaX9HE
nsmGYVyy/gmpvLn3LBgiUpmrhiu1aXEkxDA6hf0ASZvHsiq991HWEYT66ArNq9xn
b24o4/hOP0edCMOHlqe8iCxMQmyYGKpMPDXihcQv+Nnc+s+Um8f56UQGU3RTNzNj
uxIZAKOvyQp6Lq3ffGUS6ajfhEHMTE2WeMNI0Q22aqEr830fNvRmL2alDxY6LG8b
4j1Pfubu5qknmPrMN7nUV3rrHfPpSmKBVHBIAkYcOWiOhTfpgcyL2So66Vri6YBG
2Y0jFZbuAjSzCnOb/enUxNaE8jtP7hQZyVTAgZ2bIkX3OkdFwk+UmkTn+fuT7Ao2
uWzNASmCAJzbxGZwzbhSQzeD5SaxasZwxaFH3JpXOxDsyUb5jw0BBSt6/0ewgsxl
1VH+VQO/G3uZuf+eTAGkO5hvJCUwpwjc9Hsdbowy+yKxQB74UCvC/+cSdBDDT37O
5bcv63okLP92HIbpAB1wWtXjC1WvQSA3Myfw9kvDGVaewAM3QjW3zoS2Mc+d3OXk
b0jAsSBtV3RZuVH9QpX07eKSaMrIk60GKVK6uOUVeJrkNpxL79QWuGyxwyuXVbz4
22Q8Dt1BT4lD7ByqqS/MIwJeWT2V5o92g4GZDdhkAEnnsw5BSUm5klROSVXJ9OhJ
u2erhRFTB4pIiVpZgmOVPKsBeQJZZG7ymYFlxIO/ucaEXoimGcnq79qD70ij7gP1
gslyzWjFpuqKg+9dVn7LkYZ70843ZOnD0lgZqmYaAPChvxNloQ9aAcV5ATOITpz+
qba8/GeIee/JW2PFecGALi0CDdVu662lNtuAcA9pn7iixQkupUe6tnxiMJU62Bhh
HoGp23cYdfqNpXUZBKIi/NQEOBvH8Pswsp6KmM4JkLqPUpAF0wm7mECv6VVXYu7z
J+O02g34JZoZnnp0phi7U6Otxpy1bIJEG7t1kBuRs9v4hlARyXFUmDcSD/9cYqPt
j2ZwsrM4A5OwTHudupMT3WMThMOFGmD2a/hLZzEE3NPGO/T/OIuNT4KpCZ7Pocgo
zDMQ+XLdPlhhU2/GBMAu4OV1kh3nbehSlzQM7y1J2kzRXmbiwGLT41pfYmGNY6wJ
MquZAHCA7nw7d9owsg4YBdSPT7RRnWnbcqbOcvhu7FdBIGaBX0FYjjfzgQkAs4c2
qL0mA6G02dGSMo7WxbmkWXov8eyKQ8yvhFwgn40IEbFEL22HBEaeDRljJr2R7kfO
8WBBaVbDzaIrc2fVxVOYWutJ8tWmp+RsqOxXkBok5yDlvEvL+ALq9SNLtHhZ1R3D
qZj4qirmz1xRU1V2c6yKMmsbS/4NIKv2xDL9rrB86uOlUQmUc3WTfzzC7VSKzHUw
l8zbb+NE+IWsibezBCN4Z+cc3cYLfzu3HfjWKRgCKnTAQC/Hmy7hLZSjJ6ZvJVUD
WoP5pHnfrkmBpMm6duL4PqskIQMW4Y/ybcr+63q8UAwrBMNbmsoge33JWL4RKbfw
Cb/SCCzf37R3ya+Gz5xWICkLVooW3sTda+Q5h0Ppkj5ZKsh8W8gR9fTGWfITq7bO
35qq23zkWVUmW1FadyCgFRPwS06HcjvKkw2wi+JHjfw/tySd1GzZb2dQGED6OBK8
i2HRASxb7acqrxPZnr7DoiGIn3WMZ5lFz4umz2q7e3D2mYhWX7BHc6t//UW87udI
3speNJJAQdLEAwcDhZERm8sNXGRfOnoywBN5r4bMAi7s1zudEwEThOwcOeqKi/iu
LkiYp5PXKaM3xoHO3ojnWprQC01EQHc5Iz6sedfG/NFOkhusMb5ruDtm9KJIByg0
JEBby1VoaL0REDvtu+3sOz3BJHJr1IfMkuhWeVHiB/idBVXTnSdeWhAOgGaQwINW
fgjPm3e2ggJMgcqyofJn+OMNJkQYmbLdeJ8Jmw7p0xH6AFoc4gJJygM0r/tieg+a
ohFGxkPXovrvKrJZoj5hT0y7x7mMOeiWCsslQf+gifZPd3UuCd1HQ+4b8w24AYcd
G025nZjptopr/EnGkFo+wzSR0LsioFkfFSB64tDsIBpg/mOopWCwM8T7lW7KZuLx
MoTWZhWkG2q0tc47+229XEADLwK+NWFjMSWPoWYAi5HP1VHjV6cHf5DffJ2KacpE
GwsLtuJ5wmbSkeqs+zyPx/CuoK4NiJoFjfqMCT+SC0g2kWqar03UMuPdWlEM+aGF
ngHIT+qJQT6MkzBAU23z2KzG2oKUpP/beOWIqZ0duo4qacd534YBk/E163o3yRM4
oF0b3J7gdiQMwpzi++eOWqGm9nA2o5zc4DRfK0RNd6Qgu65oHLZBCuIIJrd8D8Cy
JTrSfZXfBXeRGws8ccnb9dUBNRdGmHZ5eXc3qcsFA6dHylARj8vpFMa/jiVletrt
AvLH7P921v9xdmBIrLUHUtcJ7nil6ukEX3NCf9VYrb+KAm+w2cEn1JHJClEBxm0y
SG90rnMp6CDhGq8eK29WjiIkqRb9Y4+ai7jQ4/kRsE8kAoAU5yUDzaM3j+EEhsfg
w7LAXG0jIrjDCkUA+0GmgH2O6lfhiR3pxxT3xODcoV0MQ5drocAMl8suTzB1bioV
+05mP0TZEK6/hppFHZ8AJ0mJS0CApWfUikDYZWoklVXY3PxVQh0OSIMVj7qNqP02
48MZypZ6llnmgV3UsqKkptmfjiinUjV3y/lc435cdL4Qfw0n0fnVAAvJStK7y+0h
OqA72b70V+Mu0XOkLcT1YtRxlKu+E28WLnHpbDEe6D4VmK0FFNfxRXcm4IGn8ZkS
y4UxjZcKnmoqMDGOPiMQJrWvZTpCGnAM72nbYCcCnbP1gCt5F6fMSNNa3cYLP37o
DsFutHNRKpTT8836myNRhouPSHvf1ngFvbypevWtnfEoqfAJi+8anv/4hs8BjCDa
Yq0ft1gOwrUZNjVQaUBDqz43qycAn76D0/iNtuXbK8dkVaUPEPPu2iJIDb3GPd/c
sWcyAJRyqQDcPzXuOu5uGOCtwxwfe7gGPdpqb9um5L5arii+NUk69Vl63ZsUV2Gm
93G38XcWVcx4OaeIDZ+4EOh1E18sl7AinsNRW4kfgCk3G91QPKM40EMNposOhrmc
UuD20JbXoDDaWQ8GCwNNAQ/7G1QLqPwimBf2FOpUJjtyMySTkY2ErnQFDSQWLYOf
ZHfFBvLVKH4hlJqEfH/1PU6xplWZdEowPA+v1w710twyJ6E5PmMQTXFh6YWEO2U3
kjep56kNYKWHzVltPrReclYE/Ny39WH3hxcmjNzigYifx89O6XMlMWl0dquSkxTE
hFndK1LyO2NtOQ+R833TBM3bnoan9nMZTbHeWqELCZUz+TAph0Zcj25vNsrY1ziZ
51XQR5z+cru2Ys0e7xYd+/1UOrxPY8XkYiaXpKOahe0saQ5XrQpxci57aaWUR+Ns
QxHhRwojKx81lHkZJ2KpkoLH02z6SvqrjlG12MbRu4TeJzhkaScbiOX8f66bhzdA
p0e+5bpfMKGkTtJf6c49pwtOaSnRjL2+OBuKb9y6fIi7lIjefzPpjWMakcjseaBz
pVfV4QgTzP8RVwWlPYYZyir08c17f0943MjCRwYrCZ7g5dsJxtgoGVfE1ttVzWym
l306rWjqwdsJLrat6ZVxUhZ++s4CSqM4PLMv4DkTxkmqY/hkq2997bCWq9TH/KRM
ovGQVVV9DM2J/GNkwpPyfnTeJgU+pK/4TiP6z6DQl2c8mg/TYbEtYzL6hf4Z+8Mp
h3RTB7eC9I07Ycc2Xyrxp6KAe9hsYGcELnjUBHI6WJDR2lPiLlzFpKusHi53vC2f
V2ByUeuoI0BsPOfSb0tisbzyFYakPaRcltCPJX+h+q0oW7njGJzK9HiRYWkHLrP7
3eNk92Hmi9Vzd06xFDj5YrYLQ7J3zwxmcqhP2M5LV0Qx+maN8N0QDyAufJrfsJ6H
voitIkxvjBYxVfic+71wx6yyfZZ4vUDyuzmwc6YCXS048nCA4mmBcR1Lqv5zWFbQ
ear7X1FjrqHsfisqJJXRIv3HmGxQeB5NFCoht6p3/4leowj7PD8SUw7Y0wjySz4v
8YC6WuKdrubAOTB75NP7Cv2dJvWPT1Yi9dpwUBfKhRxU43SbciEEwCP/mlTqsEf1
d+U8j6SeLWFlVVRDAkEYe2jCNnNHhPTSenFCP0KOz41Z4h3lYtaGP1JKEwd19GQK
ssYCfsrLJx4VAXeCAFa7ESqWkhWnTkoX732CZAq/rafICsGIHqYR8HcGQAbTqwo3
DGJtj3J7qylHTfW1vI6PD1okuD+tHHfaeROVbehNU8AGzQ26Uaj9mXpVSix/kzw3
IqdodH/gf/Z9wznTm7gNgdWoGjfC9teV0cAnQzRoKabkt5ufhvdPlmIq/fpUNKg8
3uj7MMCq3YACV3gQltv0ZARwsbq2kvJuthpyynCKNpaB8rmztVTOCGt5l3K+VUNA
pWfQ7Q+iKIcwiEXSI7u2HIu0mliKT1eqZLTks/Gwci9x8P6xe6X3whmard8DRi7n
dVSz9bHWe5E1pBkuFjdPnldMldJ6laxRqw/zOkTAKBe5yTRxdv1qi57nI38AuVrk
9L0l98QEVgMeyon9owzt9uT7b5xgEYd0IFlWgKfyDaiSBzGIFiw2VDf5LBf5+YFt
7Yh26CszfOvPUoTmLFo45+GB8o9uBYiRFYAIV+TR2w5kSa1z1gTzjf9lFow8Gns6
HnwNYo5iwhkYa5ZbAmNFnvAm0mO8RP7bRabO/j0wJRTeL5685MzjFUrLP0maQH4/
hanH+HVs0+zAmXymFed3QdT0nmP0MKSiqzQ8EIIYD6pFPQKDcrebw2v3AbuXL+DT
yw1FGHdvlFKmqttYlGOQkIUkCaETF9sMSQTwYgOTuFYkTgYGAGhb5+ZcqE+vpqX4
rvNJ4B1CeGcDd2rBvDwJFE8YTFXvxz/cmTg+aAxuau9DvmWeopdXFSAm7pJA+XhL
52TjUq9zlOtsEnry9kW7gJW5uVP1zwExpeE5h8aIyZ9itF29bQXbFeiWlsuyAIeV
TeLaM4aB28OS46NKNU7o7qbge2DXt/3UE36N+FMPFp/LDKkV3aSzafY0i4+uzkfe
Y8VU2bZ8tU99aUBwDx8X5YVSRcChBxqN5MRsmUH+kgQ6nDQaYATMKfBzUmVzR6DP
wW7+L29FTCrX+E8hYzdldwCdn4NP4E09Tav5X385cHjki+kEFQDgB/kGrws83OhC
9o+xOYrnakh7fAs2aYQeP0K9Xz2DOpaVDCqVGCJwIpHRJgOsi09oUN4lUexNDDAm
4XVHLik7vHADuKh4RA1zvcmaZ35qLIHeaoCZH6JiGNCK2pRz44KSobjlyXdlXXo8
CaX208/8eCxFP2DOGL3YQIdvOq12Yvh0jffg43RazWMlU1/3OJ7upooPokew+LEA
xa99OGzGtx66ud71Jj3NCSaLHgLIIdV9j8C1WDYyI/lkLYXoIVqupw7XODJtJI4O
6XZzVhI94LU2U3STN58Hnr9kTLjQHDacIGilRSb4UYgFibzqeStVZ6vUIz4kydMZ
N0R29Pr5UOMxkWrYFfnim1bHA6LImTP7LbEWgFp3ZLb/K7tTRiEww+7qSlwrzcAf
3v5EJ0dKanbOrtkErKQyqDLkLFpWh3wGVXanl2SFR7yPRG4NuOLMUzQfZW1evgTu
Vv5RVygExhAEtsijMtOxqU312Gf1baZT+xZhBUUt8BIrw0HT/HabXo72D8OsS7+i
wd8zgd+9TlJUBLd/MO+PgChXfUr7rPdxh7CqCnJ4S0lfxAyBj9cZnw6W+ZnnNHqA
RxRBw1m4oOajwdALysi5Pcxdvh1p58RqgSuN3IyO8gMRFkVLJENlYitjpEW33OO7
l3CcmvscOB/8GZwv2O+7lvWRqiHEre4UUSjXsOhZt0ziE1PUzx52aKpkuZA2cW9v
b2in9ecsFZ1jHfyB2K8e+XyT8CU7y+/Gk+tGtYNC9cuo1w/kFjAhVJxEsnq7y9FZ
ZhNMKyslzIaIQubSQ5ffk2ocZVFkcuLJjoY7wmXp/6XLXw9N6LAeaTw87Ls0Zboe
7MccAIVbLVLhXl4ctu8An8SQQYiQib/2WfO00n7gafHfhFujC79K/ytAcSQrvtDh
dz3mVeBeRYb0ZdRw6B24hy11lifjrcxQ26fTUSZcSmwMhGAHatIIMan8G26rKqTe
8CaWODdltNb+x1b9FM5ZXYXakx8JmvkLHQRIpW4JYHF87ipn278HLxPYXyIXObDM
wAOezSezwhsQZ727K4NGYjYpk5jEUMg39kSn2vZ25fGvBI19gZP7tNRS0mE+Cuv1
0g8pdtD+4KZsG/fabFaoRZF0ioGimFTcSL2/sCcUGDTrvZcMaXlRtvooZQ5rm9WY
Y44s/URuWLcPAVDh47F2ER/AVSEqXLeIwEY8Wg4CqNiHgTVtCt12xAvtEWnXLeYZ
4ES0BvIfjk/YAwPpLn/rEwNCkI2ammKOeCY1B/5b/TdPN3eNR0M7uBYrBGU37AMV
odmnFSMj49/ZTJLvAZ4GrOj5AgHyeVo8Ye9WpF5DOB8Ab4TAKTLxkxXzSRCZyAdW
ZTxnizqSGVw9l6MbfslAzoXAZFx7qYPafhrXDanmuIUJ6FUNrRLtNjeUwRmWkQ+K
uEQ91Baf28WTgX9Zhtao9sAwyOfHQ/IshmuMrEvShdevBxfUTBS1j20Y2zKJKecL
2EdCOjVz80d2pVEwQMvbISdjEyRDt2bQ/AKtz2bV0lUh23rVfdXkmoELqcx/MPAM
CA3Tr7Wkk6krtt4i7c0ORAERYHyszeL5qn17QSS0/wSC7pdAwzkdlBPqd4aNlYsN
57VD0RD9GqpzMBWCPLw5fqp4+bspIaKjPXzOG3qlUtJ/TCZC4CJ2oWSaDlrE/Mls
ZXgXsORCoRmTsF51zjNT4oZ8v2iO4F43B9j2D8Z5R5cyeyje9Me9edktUJhp9rwF
gRXTfGcJ20a7y/+N6kiWRyPF2UMxTjRbgnebsGbUULIpFtjIDsgwOfiZacTWU5VJ
2aKThKUyl/zwaC15hiGz92GhxqzLJvICmYxMIko1/U/M89mhGvaGiU2ZOLfADtzY
trQG1YYaUH7Xc87QhM2di9ABd4x/TmC2l0Sv3OvH51nDF1bgnWUGnxYpshOJRUWc
SzTRMaF7l4vUt26SRL488j8shRTTTI21Mh9xFUo7zoVSyq+wXDVkjJ9FOs4BFh2Q
AaEuCD/yD6O5OUOiQgY2rBB5KVVqSUYbPdzy4MtG6HM0thcNo/Trp6NH3jQZ/Txe
omf5+x5BS+/sNa3oNvZHxwRWqBgUwcz2/PMOBRUWxqMRNpGZe61TAAtg0XShZX/9
1g1WJDJn9BdrqLWrgfEBoIQp+udguPiUD7ZkH5iYprdm8JD2K+rpmt89q3eNbpv7
ZLKdeeUgmJolXy8D8xpaTNF+aOpq+XJ7+WwQptKYw2ckgijDByDA3lAx251oKVgj
JfNfZqEO+TrOu5NqOPflYYcZwz10FuWFUeu9VI+6yIrTU2dE3+mdtF4UYVFH/M3J
ql5SKoxcgbSVGenXLLPk5YMUvvRMItUY1ig7ouQI1jXlQL52RfEclJ9vQv/vE8Kd
KiIa9TKFagdq7+fklNN4LhoPe2zKqa/MfDyZnyL1BqTb9qvNxMZEdivoY+tYegYW
asDamDqawUhrg3mpOFV14ljSfAnRFg/gXaVwjSd/Kbj4t1NleO3UHOIcGPHWZOzS
6UpHYwi3Y8o3kdF77WRmG8IKhPKOh8xe6NDTvBS5dAeqxxo69FwcklKd4tCUluGw
j7vgp5+h8o8GbFgqaK6WKPqFfIMYCEckO4KMXDaKLGhl+9QfWuY71bA5wWPOyaeg
hv0XAVJHl136dXJhupTNEzpzOpDNQnMsZatndaZwPuTLYU4WbkuCTsaRPPK+GXk/
/+LRD/Xe1nO3CT48vag8jBAPSC4Mtul1CCA+mlI/37e/HMZnTzfNNEO0zx0EiY1A
FIKzJInjpLeUmV8XFIuMe0v5Hkea73xfA1PKF7+DqYhqETAAr5SaZTB67ZpJ8QvV
h21UHPvB+AnwsIOLgCisGY87R78D6apxrjw0tNLPzowz6qQuT1uO/roRxIPgebJn
aKkprEsnQS9WLSwIRDkWGWwlTty4kt/O3WvFOn5yQlaUjb5HWhM2ZIDMoWHNAbY0
AEjtjqbmLbBtqOXMk9PG/LH7GkzFqKSWoicz+MP1yGG7rvr/cBC0j8MdADlqqbW9
k6RAZ6sVmqoCMK++94AbQVKpGpNkxURWLCVBE1TVLhomrK5B+pBfab7SzZCJ9NJu
swUzeXvZTNSLPoX+5K4OVKBn0IfOw8GCAcPnVmG1CQ/tusQ4WFmuuD7FgiWHhxcm
5J/fI3BD3j/eTvYbgTeVGv5Gchm44+0eG8VekbpW/bky7t2Koldb+YFuPUnJzxm+
3l8Jw1c+dbRW2RuIQXzQZgnWrm7bUfNtY+5sfCxgJWbeaVl4TgvMDUKvYMBhGzsf
Sw1e7h0AxTvCggENRM/odIhtwpypykj4elt74Q8LIQQLYqzkHLeg00ZtMgqJbRM7
djMZ9Tq5VZt7ea7BxC6q8dC/jLQtcLiuw39Xghy2ylfYntnBMsKmrY8gObW4iGgu
exMzTryZtM7UILr3ki5oAo7zGWZ9LKSd9XeG1/3i/hgl+mnYi1DbSKENZHkRB017
5ZlVcgB+V6ZMyjUiE8GNrVuwXSIXcIgjn7FFlt4+PRWaTRVbLWUPQyzusEXz8+U+
memDdgqDwnuGr8Rn/7PE9pWjpY5gtNkVOBQ1rXapTr2fK+Z3c4Zyu1PZFJFb+7b/
PfhUKclPV2hGFbGW3zYDe7U2Jh2DpqqFQNF3SPg+M8Fs3MXKSa2VGFSn12roeZka
W5LE60tD6DzDnJ7OqGU19kBropSBG8MTBkGFN3XNQnICsBnaUjcH7Zxa6bkWIe23
yW9Ml6tm0tGZQEXyNsTqQVkU7u33lVO8t9vNAUsJq7oAufeVK4+jneQIap46H3ia
HQIujoNytje7xxxfaSzAE2zVsjCgJjM9X9zN8B6vLB6B+Luz99gLlubQNpfD3KML
bvE90/aDscIrJcxB+5QAGzifabHeA/esz0W8pfIu4FAkxwzjtsdSxRAadHc+vq6I
1mdI2JA4t9nFNbWUtdwyAPa6It9N4tB4gyMXzh1/AwagqL1EtUVC8Zqj09SYVwZI
WdKu0qgnjTtv/Sp+nhY4kq4cBuUIXoZcAuifoUlsyvflEc+2ZnfUN5Hp/NumshGU
RVDyChX2AqTRF88pUM1K1NSNDDCzNw3BzAsodLMQDIfiIM0OOTn8qbPebmgoCU7H
zDqAQZ0z8OgBxpNSqkJDrO5HgDj648+Y2Mpqiv2L0R9eylEXmlvaoCPjA2/BkJ0i
2o9LWctjknBz59QlAuAfA83k2f1Q9s36iy0aQOfnJNrHSpGZzHI4cVDsVXItxZ5j
8CChImdXrmgXsA7Sd3EBWIxWncj6bLhKrZUQOfAF0Vzx5656EK6TDShTBSsfNH72
tfqEfsOOLtnuNG/ySzLcPcsmL9VIDBgFdeg7u7h347WrZFdYoAGhn0MxgZp+oG6C
J3xGM5eGj8GePuyCu8aHnBIhh/X25O25EQeg38sVFuYXurgpCHSMuw6NlpAnpKIU
tnsPeozrnSPB1pAWudYddMe8IzkaHjjNzsU2RqN3Lwbf3Uj+JrTN++Hl06S9AGHV
6gb1TkiMt8mJCYWAXCXGlhtHB9Ef755NdBY6mxfDSj4el2zagFJMmushi7qi4vUb
IvslrODYEnXhgXaIqozWF+dfJtxSmykrssvA3IlQ3q3Z7/HVXJFyYv4zS7rqkA4j
uwopuI2QG8fgcTJJzq0quvvW4OtW8ALDYg4ka2tEBBuGc73lbiM9d2TrUESmMUBS
pSsp/n1rJadZMNxbVhLOzgacM0z6133gqSCwcbYDWoT++kr/x2CScVdfOoi1PhzZ
u02xtRYO/31L11Mv677/+HVjl6rYtefMDr6RsuFfn/hPbGIAOoVL7hBKe966ewRW
emz/mFvmnHSLgcLJAp3e8rr/A6qyruvUWhnUt51g3uQCtw4J6NB6CB8YT50IMjx7
sp3255nSl2WzQZXxUQ7kXuMwDhFIiuAW6W2WVSH+5hPXnEs2xEtTuhUED8D+6BIj
ZBS/3At5YJUshhUjBcQNRb0ihWn7OuWay9zdhTx6T039QX9Rmg6jA46YvSQhPYOz
un4lCJkE4ePbg6dTN+qb7ZgKd61D93262nQeML+6JapLrFrxEJR8B50YQtiYVoHo
I9YzzxiQ8h2dH/1INM1JwwbF3b6Vx+RX+kTY11NVTvn8lc4UhMqdHYaTfbZkH5Rg
+GoD8hlWQdw+6KvbvsR+LYisxSOsgnywF1smUVhOu/YDE8Gew7VKqLm9JTlY9Q7v
aooD91uIIUCtIe4Jv+FH3jxjrOiGTJbtKfw3YnF/50495cfKm4f/TwD8/WlRb2TN
FjvZdD6nP9kkmOhzDVsWhq2KmhJB11J9we1w92MycTaX0pZcC7uLVE02TCprYTkf
nGK+T/hqCYdPIgNXJDbdA4KDBeNtKpEE//tjnU81yq756nujRqralYqxaoOrzhLU
tcDjzs8LalZ9mNg1UPccuzkTLT3GLQtxviGuDmM2g34JJFi1KLZeSuBgTFLl0Ko2
gBGbN88+tKhKaBgCMkJcLln0F3IlnMRfK7BUIvJ/A+MvAHQu8itEVq/TIqrkuOIn
rCSynsgluP3dFr7zPL0PrmWBRc0OGPu85carpZeGrGpp1A8g2km0n4AudZ3dl3Is
/oAeCdW0THvpszr2pnAmI6gH7Advm9C1lS4cE15x/NObRmmDB3Eb4n07HsSjOEfS
LuYSJvYs81Ef9pSrRQtt7CIMBqvEV2PTDRKJ9sfOHPM5gEE0Vr2WZ75vbIAAErnP
DwnqBzF+gVFuo2bZtI+/IM4E7Kykb4j8s5ei+9MN9uz/r39JHkLqntChZQUvR9qM
6tnlLTN8rIpCQqJ0pakNZuuf85f255OMGExGWLHhJJXnmiW6QPY+b9Lq84VB1ich
R917XX0/viTsfEuuXR1N0xH7t6U4+yjUrm1jrz4uZ0lS+T5GDLoQk2aUX5QZe//u
tHUpXHQit00fwMI9GDWHGYpFk10GnN+pz/pQkt906mA+xLDSvIHm8Y4B8rxFqBrn
L7UJuncPkWhiG6FaXMWwWqk0/GY3f1cSnxb7sElzs5vGH3FkZ7i42V3syJq0HWLA
o7oNSvU0rErjt1AEiXT8U+XsqcVelJ6TzbO2SDNAlXzXfFHXEDpuYxArwHdxJ54z
7kWtlUyaSw97qwGnX5cgICL+36yf4wopz9QjhJwGPWQc3goNu4wIvkyM+fRGJ+cF
EPT/jFHDEvgFHjzjE43mBjKVo5kL3GpMczbEaXH0Y4QtBhm9AyCUJKFT4CVVd4Fo
k5d1qshzZjDqWowRuBIrHePI7c3TY+KzfbD8CR5PAXKZtIcrH3U0k4QrlIHrnpP2
GSI+QDyTrYJupn7zAvMej46HS497bhl3NUnpBDStt8iWNmGeOWm4ElkdN6ASHY+x
A5xPhonhxC60/qp4K30J/krDmvJgCoePb5T7LO3Nhh/tssm3mtX5t4Vsz/PgZkZP
yuu8RKMwe8ouXgU6BjlBYdI44XMD0QF6Fpmzd3LMXYL6Ck5Yoje5sVMo/WDHZapp
cGbRE438t69qr0JwSMLtQV0Mv8aOB7DGnMlSsql1UeAgdgAqBF+RejTVV9T5E+9O
zJiHJAiwY/3EFvqha7W7aUUfbdnwQrhbuVFEe4UmfkjamkB8iQzaYswGwYT1Kj9F
fJDRM33BdOvQJjn0LbpJJhPOop381OYMJnK8g2q/ktGGoTbjuCA3WXs3k1MsWtuX
Xb1f03gO+s/3vkpqwKzVwcf3shx2aEFrJTNvNool8Zf4Ne2729r5OGSLe1vMq5U3
GauGEJ6OHOmnGPihbqflyN+E17smzUD6hGvM9nI0HdTNvyPq51ruOVu4wkO+DrN2
dUd+TzRgtuQg5ejTFAkiytjmdfevpaOS7Y0tk3ZntDpYIYvjndvY8Gti+o7jX78k
KyJJYNkj18UgK+yad9cQkIP3UWCGY40qOPaglnfiQZtvqGtx2B+B/fLPk3Y1/5o3
fWScMt9BcUWHwMIhw1cOVQUepRvHs4FB8Bt9oOVeOQSHseEqji2D74BjpavTdHfx
IG1LBQgO7IfKR/xS7BsNz50WRiIQhZBSKseBVDsYAY8hPAZ4vxpcl5qA/JM8cJRa
z4CxLfb/wEzEDDERZUcE5m/C0Df3SBJPxXdlZIIdWNe89eSzTneEpl0qTLN7tWSs
9+iM9XyrN9HzcAUpuv9mE7rFUDi1eEZyrddzlT5hl69OB6dS8Q9mcpYfc0JhMjlD
FLL6t9ntoPI1oUyfSvQDvu+TbJNs9RH/769g5NSitEv1BX/ViHnq/Qle2IpGaHCp
neCBYk8tF+aE3Gl7XuWsG8svfps9rq9htBWtH1izywm0MCCpjpcoeB+rrDyVDGRI
6Lj6+BSJ5Puji1dWL7FAValWgSWKesNJ1RPDpkGOIQ56bxjWXoutb0TZ82Fy6ik4
J/3Bjr0FQcJHd2M2TDgPX/Y57YbBdPMvQp51u+DGZ4U++GevKAdBzErJvnlTz/V7
k8WUTxMTyOUqQ/w1xZ2FOq9gYdZXbyekn5B+DhkQUVsyAkPdHMqVUoXT2SNMWUQy
gUZ5AxRrh2ndA+c7O9gDdkPNJfjBee21ybBt6xLHCzdIwN+uan2nYBJfPES+2GoG
JQ7Bwr7IKNaiCL6Qg4W9zbZztlsrpDAAF0HR9sr01DibS4v1yTJfz/wWrfb+WCKS
rfWqnqlrhCNLT/XmXsAuqej/3bZ4bfY98k7l8FnO2dID+mcUo98S8URCNDXEpYq2
dFCBbqHRWgk+yIJU9Bzx4AyILCAyFgpbt9oRHjER4BbevcSGGDsQnD/2iyXx+ukM
vUGo9yCJp/UQeSl89eWEaSaDLktQ9sr0A/6vACQE2HkQhLiCOjVivwMndJvwweZS
o4Y5A6Qng8U/UVAVvd7xxGp0ky4PbGOoulpdkx4k5WGuJLCtbOuc3prjIX7+2bBz
o+E+ujmEJ2RWg8MnlgvmUsEpsKG8mVChYPZW0Drw9na1Nucpp6fJDgOadrKJWOKP
uGa3LQOXzNLxeXBDkgj5YBIMWQzSZtG/ADgxNqB1Rwa6a/zp+LrQ4vgmNFwclRxc
xeSVbEwoxSXJ1x4YA65GpOJrNuM60eDIrE7nlj52WzsBeTkqpE6MNyRbhi85BZKj
3CBOBBDhwSHMIxPzmBHbkThS1AfHGO/qCHFXAsEr71VoP4fG0Xpz8OR2bNOK/9FX
meuJnGqggsACby1Ii58Pvzy/H0/98pCpfuofQ3fGElE00RiYv7Q529xR+dxCI/Js
6IqPDZPO1KItRq6ikra41VBElG8lFwe7ukBq3yidOasT9xoPw/uMEDA19QsKrGPu
SNiFBTcDsgNKJFS8BwgOfaONZwx9pTF31aNkgvRCxTPhZVtWHuqj/ayDN6jum45E
uqrrlygWoQzqrhxjsPE7lSex31eEfLa36hZsVIRwRakwqs+xeauTfXzbrk6lMYX1
35pFVr8rDKMeYbcBijWiiHLTK2g0N87EFmftUD9TAvELGrG9nbR+nIBgCAhy6uBU
Q+VYqi1Jz3E5U+wI0mG5vXuIP5HPOIfLhCXa/mH/ZcZfRAzfp9p98doijs2mpZxv
9NnKUqb8N3opqJHPtw4McI07PPOVTC1QunJ5eAJXnd2KGQKpU9VfYZIEB69xD75s
BtOXymGdp37lhg4DW4jFhm7r9GhxKzZDHZ/BRgTjqTO8w6qAVI5Xh+VPKrmx+mRp
pOaeLkvUElniGyIqX1dW1CPFOMBSe3ilfD83oiuIzIfvl/FinWdJ6/jT3+7ldLE2
LHMBVJ+pNkca1gtzD3eCLdnCkxoCdyJo+GZAlFjAf2Ko+LHEC1I+nZPqhazLeYf6
GCv3kbVlk1I3lDi7rQoOFhH4SD9hCbBOOF90g2d5CJPnaVdyePUZghzvhBLFph65
TeTNPlmJ3uV5dUXAOIYctV8l+TDjr7yq1DNGj/BzRpvldeO71xgcxc7rbAM8brqk
A5LtfMsMTBFl435VaXTq4BxExBOL4YfpsNfYrHcfGIsRsw4Eg5zkYbOKzDjrarOg
gqIvu04IrpK9mFpqF292ZL/6nzPfyoqQdWR9+4/+hHXSynwo6DdBJ18CtIHzjc93
HN56Zp3338iopYJ2xMMrGb9/utTkEW9DRXKMWzhp5pCVjzq0gHxKSOAW2TcwQyzt
xG1Ai1vXb3j/4Vjuuzy4zLRE/fJRbCA/etqcwwaPEMax6UR8N9aFMbS9ysNk3cpz
Gxi3EUNCjO4sYEZda7aV77GJoMl4X16oA2xW68j4gNZNqDIQ8UqIqbeRD/7JGQEz
J9FnImHGqvLBhvj3doWadAYr4j5Vd/ZWjpO+kD8qIL3KRDurYfDwsqRKuLXUP0v5
n1MWHz8fgBJBjeM1OcSVR4SnJKYUhqtARWGwZ6Qrk2jWV+ea+yLF/YmSGLH0yUmJ
rgPO+sq3I+eOEK32rLp/7mXs0PLbvgxl3I40IqIR4fDG+RNUB9isw69mj6QHc7Cy
1jXw6mn0WNthuyLgybFRLKoROtKqyBbQhHj/2OXm1IV6i6Dj6Y0xmGYPt6YRwmhj
Dyl2Ny59rJbn14e3V6Aillkh53CZs46mkanXoPdE4rLX0XYFz3rgG8J1jEMhscek
RdVFfw0VqK7ZjWmzAM1Uo1w9UeKUEezLio0RNtEQ2mpQln9uwKReAbF0mwfvpYfA
1ne+gDbtgJ60qCgvLOBz7HM/aaT7TguKW5FvxOR1bc4q22pYL6YV8O3VqZcYzmsP
NqwsigO5DewI1toAW1KOXDX86rwJOEY9S2ulRORZcUZqChHL/Bm6E0z/X2y8Dlk5
6o45puiQL27ae5EsuUO8KySfeP6Pl0wfNq29O+JgaLM6Vjp1IsHVgZLvvzWqHvUM
irqkZ90fqu1NS1nCiDy7aowMKno4S9QWaLiXTzf868SnscX4tTt97eztLwc53UvU
Q/RaJwCA1EBvLZ6DwnekAmHwr+LfZBmVtHDPHXo+SK2zP8pMo1TSefBSVybCiFKB
cqo5Bv56i5/KCTI/6R9ojROosqbLOJs7mBOrPDlINBlF/uYLm0FmV+fnYidVM2+p
Z+hy8tSbNMvlIL/uTctSn68v+NDmKBgbxe1RA+yTzL8KXF4XOhll2HDmiPKppPD7
M+NHakabbu6lvlz4deesXRwHzfD2EX+KpZCaH1on/b6SQRrCCEpOuN4qM5icQi8x
HZdAs6xOiNRl5Y3VbB2hWlumPWWjOJvHL3g787D5XyNy472jzcGwExb70/qjwFQ+
XQzsK3V9HcP0v1JHu/9kNDj39dc7DCaGHblj8aWG5YYBr0ZFjRiNO+iH0qV3kVGJ
A6kiJ+qqFMcj6f5bzK9prgvYcrqF1FbGkZC26pFUJmoHzetKStEz+i3C2SWz5X76
AeLYf3+oP0kzVdn2QffIcAuLo8lCKQJh7Fm3Nyyn2Bm+RAwLmdMR9CPpcz6QN4Fm
MD3FrSWMSggKOeFIBu6QSChgUmhLgJH7XOmF3tIyxi7Q4EEEjO9QaUlgpdIjBPor
F08ACsTNRh1I1dfljhnzu3BvIECwUMxYmkzpNTtjEV2EGAqaEiP9nWdRavkbEIa9
Itf48AjGmukUsTbMCTyAt8KN+py5prbmMZpc/76arexH03Rd99Gm2khcdQlBC9qh
M7r8+nDAKr1h4W/W2YGMF2QVTqiZB7VVhx0vYPYEJkDO3NKjzFbCraxB+wyKeFMQ
J+x149niKLJc0dB6VmZWpFbyh3z8ihy7LzVN/M+ydu/NZsp32kuf7qTGRfgYK2kd
jd6MYvBVU2NNxNWXpwai5wb9Ebt+zE7dUEhZGc+ukWGw0t8PYTNKY8GKhOPwHeB8
AGQZLiu+1W2IbzQhUT40OQwhxGmyaVpOyqKbFRTyRDGUjBYW1GfgzL9nUDzD5Mbb
IDK4rmd5vaDJJCCFoRh9wBxeJHz+t6XNc/His0O3lBDO0lQvF/WLOC0TYiq/0fNG
ZKAqm9gVhzSOG54d/UXND/MDSUP0uJy9rUDspo0kBZtaVr5GI/UrrQPBa33/pXz6
0fFksjDJrzGz0KSrIgCnXhe853FA6KS+hBXi/rxgb1GKQORxd/W+AJhUUbCAHTUw
tT5MsoKs9tgxiGR7rjPqS+ahUTNIdxUz+O467Gto4zX2DjdiNKf5enAU0iDiZ60w
E7RvAaeaVsN+GEVkVNUmvBzPrLYf/3RtD4g7QxLzqJPk6dCFYsOU8jfM5MSQnCR8
PjF2RzsWoq94HEbSUSlETWqc5meuq414KvzWtyrEHBeHNnZDa4aVM+d62qXrUEpa
mpLPluQSKvGuDE5YM/UPqR8inZ7BSfe5KX41bcikwpzyIR8prLGpmWXfxQ+zBpxs
RoshiE3N0vetD76Hit+caIskvtrWP6ZtzAlTtvRQHUDRQhXk7ivqTDXyWznqUs0R
MxIYSa8aOwDMLVMzMQ2UEwazQRVdZA0VjDec1QXDGUDOjugYTr/edpr6X74Bt6DH
R65ZRxJYIwmXQEAr1dTPth30cyDhQr/rAFz6Us2hBBeLdXWM4GKUmDHgLrbISpmc
OXk1Ck+J2l1DyYicmfVs9jglhoQcsKwcAaCwaoOZYhX+FEtUpy+4CucY6ustJhN/
Jhvl6FzJwZi6HOFGfSCKADelQ53c50ubPQoOlw4YSLrTLYJbeT0gl0poqQ1Oeat+
adMXJKBylZVcinehgo19+aYTAiXa77lBeFAWhbs+9U0OjEli9QjAt9ImSniCvrwR
KSx0kihS/oPUmJKJNAsUF/jEtQaELe1ZMAo/L3T+0DVrzUETUeFGCUhKkKKg/0W3
VZP6UEqfCZ+kNoafr9Nuts7Efhasfyfb43NtqzmHS0k2fvz0Kr7rZBYneW7XgyRp
lXe3BtFcjT4iMSUIxmFFPCCjGHnfsjTJlQxPJ7R+uqnBfGOoeE/8MjW81om/UeFt
f1J2hoOhiwagAatHivb4TJ0CcAye55daQOaxM+umTDIq41on06v6B6Zr+MVEAS7A
vA2WPTLNbENtEzAq2f+7IwLBo8oQo2LgGtcXUrYTf66JhsSSi0wDLjqeN6ISXiK0
0RnjQrJS49Vvj+PE/cAh1dHlQMdrUW0d3HhBenpIU11h6evP0rL4skPFiPwYwRCL
egiGFUuOelM10eAcaR+JQRUdJOXKE3SWR7NcpYX2zaX0uygzcAD9yQCCPQjSaZ4q
6CqUvIcU4hwKT9cmyo2vbKRnod4tvoijqkqevYuwAEPoVVXPztxsqOaC3Fx5ucBV
nxdYXlHwusmwf5Lg/HUpOR8AHcv7pYtxTV4xOQx7bcz8Mh2/sLHW3a9vTRETsTnX
bfa49cp09smS5kURvP6EyBLtV75+G1g9NXzqOOynlwY4S02sZDlGKS3DajXnjSye
5uQ4JURHMJ5Unjsz1wogE5f0nS/Ja4oFYHvnZKPYXtRcAzL23Gngq7eq/8ShFWhb
segwljJWyvyYsOFO6m8hMWDfXA7skxN4sWC41eQ3Lf/5nrMGoq7CQmZj3C7j93Yr
KLvesceYDbrllDZYxfdoxwEEbbe+Qxp15dSQrs74vbbcUmNN4CSNKoRLsx3gaOxJ
vMPLrdPVMWK7pVGWNTMJJtpEXAuNRo18Rd11tbwzdsfMF9slLN3YIplnTY0eryax
T2RI3/Ued+7/K1x3zjRrc7f5GBBWQexhV9bSj3zAlIi9YVLWulcujcHaP+S3Qjrx
dsH61c/ZzYg6z57PlQ9+0WifW+8GQ0yd8tPc47u4KudEzdthygfNNYTTkLHbXV99
tNKWpQKg0zq/X0vv/skvdZLAYdgD9/wUz2KiB8BvL2RjukY1KucAL74q5HsV4bj6
/8rzKjotzq9PBe3Wmmt/Ss7qcekHbM1pCiqr3QiPzbdHgGqbh19bzuLeUfS+VgEx
ZkURoLX0CZN32nhdV/25lvWnBRgu6bbtpOiNiNrxa7tLnIzbHREXNgWTHOtJmBbx
lOahIrOfINqqOAOHAc9Mu3Vnt34ZPXewtvSEUp5PWUz/9yw67VtxuiR5sTGOuaxA
GmdcGu56wikOdRNDImgheGL79mhfdmsYyctusYNvetCJSx2Rtzr2WTnZ2/9y7UGE
fuakEwhDKBZ5Yx2IX6g18PkNT4uMANZOZbW+GXP0lXU0Aq12gDUC37Gp9komue3I
5hFKFtaJOE1ZspqCJTr/pbNz2fCflmSLm+5USaXhr9cAPqWpS0wp6aRyggkjyQ85
Z1rXJrcGmvcmMjn/upA2oo2RP+UOfCyHT6eaJe5CX3Bj8xJhlbgslhhT9xBCDmTf
vrwpJYfe5p0ODtJz0VMb3dfuK1muV6+ZGE7nsHtbwugah3w/kB51EyfXWrUgh6bF
LKIOq1dnGZnb9YGH1kMhDHVrAq5D8/YsIj4JQ5jOtm7kR4MbDgXeETgUkssMwh3z
DJ+sWx02ezFF9X0wg8h0eb1N8wO8Vtb0oaCoF20gjI+LcAPGHS4rT6D5QDGb4ILE
7wpBr/nGZbc0XXCSJwGW6HOHwayhDsoOgUN3x2754znFNliz8ku5/cc/IP6SjA+6
KRfuy10UNy/Tz8zTXUpX14SXKMJmEgKxRWr8QoHVOc9vTeeCYcAGarlThwIjXR5A
CMjlUM9B4gVq0FNYfsGyHf8rkqqupN0SxR6auXncn7JLeao7EXwhC/22vrKY4Ef5
EW4zbLDt/tzgfenLbhRjAx4IXQYy1dKXdHV6WyojAK9l6jFNn4unbtg4q/Hl/G0Z
h2IEwAzpTJgjJUf+YFGI9KSNtH1AcQ0FY0t3GncTHqvB1S5xUcXzRaE7ltBTzxAq
2rSuaOUbIi+INaQ/k8JErXjq+gDtbcMk705zeIV/YXqA6oVEuiEbSaMphEBnLo1D
M6gSlledmeAOy0Jv+tkT0u81uFhvWoIXYZB195jtQhtN03ITq/Of77hxz3f12h8W
N+nWM/pZ/QVftL5HnP8cfNsBNgJXwJYwQGrT2xwkzP5gvpfztbn9pB0192f+uEw6
3nctICLz9rZlYNUwy08NZ40/pIbtd4WnyQa/5HaXnHkYy2pseh2u/23ieGEpuWuY
RY+3fQ40WHJgtAhLHcI7k8Re63A+a2ti6fTZS0hxqqQVIcUuS4dXF7qln+yMSNmp
0OwbU7ZQblZSt0b/rKYRCJAwfCw+Qvc2hvG9b1fHllB6wFO5wBHx+zapLggL/rrP
unBN3wtIyDEDsYrj+ficrF4hfEyBmojLYPwgmItUK4m0zBClhO3SJhFRQfq4bQ8l
nKvvpAR1ufVnqaoX7pmeGhTgcGaaPH3hyvmtahXwfnWt4QZWYYrUnGs8w8YF/vWm
Dyo9Aohhl0aFyx4GhXPRAl4fNL/4tHXPf1ULTTzHUmA5R5/DUsortrY6rb5O1F3L
hu/SUg8tSKWgFAFIcFh6SpLm+q7tZw5WDLwpUchCCeG4iw/b2yVq2cLfJfMue3Vg
RecvV45zi4u/juDaI4y4gH6IyDBuPvFXm6OyWePEK7PKlVkUtudf34p85SUAcqTA
GIB9H70k3jl9UWM54hWTKv9Pc75T7zYkrySZMhrYKapO4UiGYCCcegncWRH6LRBS
GcNSh4wI1RlQDC109Obmvo6FPP72AVw5PiNm6MYArtUbRC+beG+TzdNwgrPp+N1z
xcVGEIg+NiwG7ahpMq8k00DriKUci3WsYAWD//B7kLpXP9md95ZhModaOyl4dF8l
TlSagToy/JH5tmvyPAAA78+NZ0rEOzy7N5fmi2vKn6bhNh39XN9d1GZziU581HD9
Q64dZSGcKTqN4tqLkkZ+dHEPD+2DMTle/VVCs/JMAXdPy0SjqHvwnUOkAXyqSIPe
n7gQT2b6EZvfBL5tBumeud9vpRnARVb0hBfkG9m6iDtpu+Z2qkIHmyOBoTkEpTy0
y9ZEnf1uvp/hZ/MKNoRxNSDgqIR+F+R9jn5EYojJskY77SbbrBNW09D55yGCitJU
lD+x8tKrq7thbqiZ9KXeQ41KS6aocr+SrFPQs280b/e1T3X9i8kFlzvGZdFbBp80
yU9uOKQmzKvaYjKBBzrPnGHsNyHYmUJlPM9RSYv8VReW2bfweytzePcrovl7m3Ln
GSoN3dbXSQx1d+zKt9DWe6iAcIgxgSB85G1IL/oaDi1fHz3q1rdLX7Cwu5XiAgWw
LA/F/MJmDwXHeWmbC/yO4ZmT0yqqCZ1PdxwUJGn4PilD8LAM/5nleDxgqudciJlb
UMJdFAm9tKB4HZA0tx1MsnBkjcjRhzpUEaiCYZvOS7LQx4jlAVvjA0II0eEeHnsx
kKulhdBsQTHQaLa+1SX4aTcuxgnnENosFpaPYEBzWesjUgiqZnrDxf6U2HcOkgtP
xSZ8c/UuBPgmjcWK6b4rQgXA7E/kTG8x4KvlIhBlZGTN4+EJF6CTxzccETuIkEb6
8TvaeTo5/iKh/aPrMsCYavSJM2CkXTxb6m2PnaOPFzRdj5PO0ND5rU8YhfqIiCuh
nPj8losAePd9nWg/DtMDnwyCIz1lAUNxZ56uQ33Rf9mZ3aS/oQbpXseQUpN7jJQ4
65FhhiOa8zkSpaXkcgy383IxNgti3wPSCSZDFUeqJXKXzVzyB9sHhopFLItYXhg0
6kGuFEB6gLfkPvKKBBbwia9v/PRq8o7QCE5r637BpwLkWWB1SXmZS4/aSpM/BGOG
mv68xilxV8ckEgQCLt7cMGQd3BeDO5iHj0USiHfXTrW/SPRaKCUDltXhgTKZ2DVb
76YvRWpFOc37hjYzpZmqDrZrCVxTDQ4VOMki0iZF3Qj1JEcdtr/+nup5Wzp+Wif2
crLInGu7c3S3ltq4PRa9LpB8NAPp2iB7uKfaVkNOeg/4rkAWkC3Mmayev6o4Q6QL
zWFbeRnd+cVeyNhjoIAiyFTCNyi1xxghqT81phJ9aNFnInFUTdcz+UgQkRfBRipQ
eyomCjFG7wSFi1lTa3IL51bLjb0HR4vEQ2Naaw0CNGH5fC0LKKdLUzN6ZYerATmt
7+iokMqC4HXHECuUy0XbevPY8lxl3NycK6agwIOKiEC78ara82bkxWMftZPcCbfN
jMKLsIAjnmGD/kG/04cCV/zrof1pzXnAc1ywLFNPTq+c62SyqwCvLmXEofEpGV6Q
NlBNxoPAz4dPdPznZQAX2YzzVKPwrt8Z5o9J9/WYNYBSmGrKZLE+paUPBxRSjrB8
3x3hZMxI2sN9iOYmtoiCcNvZ/WXuAwBDR4ShjXTjpeHhFV/nmeEgWRSTtgoNf/AO
d9OApS2snp1urqDXVA/EMSNSFmJwPJO75QpoOTvhjSNf25HyKiVy8jJdnn+9xSb8
mpwoBDLxpVqgvkP7toGIexHMJDa6V/dzMadnlvUJcRtpcoRTUTfhgciLFvFOlkPS
Zh+nfmnv6hIlo5hmZu8NX7D6Ijz5k5bHtyMwdYF0j7i8XLO0fhOyqcLf5nWdu+Ra
ZcobEGtOk4mehe1cR/kFaENSjrFevV1rYCtrps/TDK1plrA7GxUO9ZuYOOWrVbSF
q54JTlZczrIVqUFhQD7lY0EtgLSK/7egiwjTg87Jps9MEyKZBC4uFhuxZ9tRtsBh
PQ1mgruWXLarlFUEFxsWKBdNGXu5u2L2qsYLGtB2DhMmmQi3ktvFpvOyGBeFUb26
QsIv4h/G90vePynZ/BP8xuEsMBHxa7q06abhSoeDzjhIxVYo2ftRaXX/whjz9e7c
WVC9i4H5jCCIvxLyoFUuKXdRaOUlcD2Zk9xU+x/4vHK+qXMJXAm0ms1Sbheszakm
gK/PJEkgrnVJN7NbjqngDDnJlHwVC1Lt81peXiVEjwxH1oiFtEW2AJkZnH3xuxpR
0fkdrhVYMOc0nmGBvwrLVv6U271bzaPAOC0bVnW9C+vCg4Lb0yacN1zMr5s+VBs/
fIuVT3DleNfH6EOaO/HoBKnoRfUYp8z/HQzM/hFJsBiX+BwvSNTpL6QANHdyKIFE
Sv2+K8ccZMXK2BvtB44nMRrWQbhGHxuUBrr7gqVNgkq9pgM0GnueVN3iX8tS/dl0
ioW1QMcrxbWpyXgxpO0zmxRypi8Nglj2EWUlKBXW86O0J15PX6tOdlQG3SbiSnKi
L6V1IEh9HAy3zbxJaDbmMrGmUxJBZZKCZlgqsDz/LPDR3+SdneuT48xkAct/BKfx
WkU7nyLsQzEw/Sb8KOUpl0M1NfgfGg4ZqSQUbCSq+nIT3Cvua7vHDPOMbV8zeINc
/rPGJ4GQb/gwA1E6kGY3zQVECViMR3tfDNQgIc0NKGJ35OmxIhKMh/tcdUTNj77o
sHXzsITvRfMjxj4Ptbha3g/0GWp+rm/5C+SVcCUdg56QmJY8B884dP1pctjjgy03
Va4hG1cgZSJne69gmr/M+p9P9XQ6yl40SsagbB4KjqGISoHVQUX10aHmCD0OypoX
cjuzLR0IKy2SG0oVgvtjTIGEwnReu13sNYs3btmO6UdTubb2x4Sv8tpwcMKMx4fg
DUki2HwpaeMYgRlTGfDEWhFRspJZzymPM8yUyWUh+UgKDy4wkusdfnD47IJYV745
hX3f3tkGOo+1mXg/SM78jzIoKroPff2sS/l9Qjlk3a7UYVaNnny9b3qLiMZqefsN
fwo67e6J7S6POHroFzA/0j6bj/qQHxcEyrabgpWjjtCKAJbDi7sBMBgEQVZF1J+W
Hd74Sh66IoxyP1lv3Y3PzFo7Epo3R0/HBUioe5li3o8+otpux598uKmneS6l+uI0
AOmK5PaOkcAEvhDWDjd6d9NYajVNpjAlWGPQBQXaIPPBfZFRk2d/qE3CeMtpQ2ow
nTQT+O1+y8CYJ2feJbuVEpZq/Rdbmy56y1TswPr0USntbJJhK9EWWQHLYfGCzHz2
aGvKUvQhOTmIiBI5U6XR8JGIHtDFN0fJ6nE198MNWViErBL9kubVGadsUYgS090v
mqbjdbmfSLCOtfJFbJI7u5fK19SAb2K1YSzPJO9Jj33a47vYiiMoeI280PJ8DYWU
r/d/BGl0xXiDmsCqyz6MzzI0zHRCSA/GPTgqJ8tRKQcBej1xYAhtVtWwsfPWJi35
KCMuBPnm1oVH924UsUIqeZmjMg8f7n3DWFA3lI7j9y2pbJV9YQMHWYKFQpAlLHJD
P0GUKKsgebgbxuYPYKIXda6dkG+C7wSZAjZ+satc3Hh7L/5UcXFfHHmCIXcUktsV
1jZwyDK7KUJ3afqb/AccdTX5d+KrEXxVqCCJa2opLTPNgVIJWoiAf+5PLZZ++3Gd
zz7uosUHGCNBzSNSJDTIZjIt9b8tjYnPtxEZ1H0biIoyGISwicjMs7C6n08mrbuM
zmp4KE9PGAYJnpzsl3Vu1BCdxKyj0ZsOVbIuV6Q0cW9pVUHVmRZH4RiCBY+P0Vdb
FrE53PJtvh5zJu+3ysKyq9vtdIKHjdCC8f0vdD3hFzfnVy0QsUeJjlXaR+X1juCF
lriKmVjt8mg7kj4dFNdf7iLPfjBo4OoDMxmXvX2zUjsZskOPlivZbdcuPbpIKpL/
/LzFJAI/xJ9rr6CTg1jXWwUVJrw3PoteucUC8zo9TVHS3gWYtDk1nu90BBepxrZY
ETrnCR7b2BTp6gbxxXru5IdlzuEMwbGpGLwSR3kNL1Yj3UEHSlMeNXIi2Tx6U+hW
Yf7BPjLMV9SDUj3mvr3EuY4nuT984BhmpcS8BRa5Ka4TwLbNDc9AINXsrzpiRe/7
LeLIr4f+Jd0o3G/cOpHQG3VI2Q7ZH9+eZpoHP40LiuaM2k/+p/VtDh76UEl1Za8V
ufMcXFs9QJNt+dubu9KuDwHc9JCIX/QZdVwpkpzpdZtFXza3YEQvoLegtsf6HlBM
H3wk2u9HkztF4UjWZIdx2cf9HrJvf67dDTyQcTr4/pnTXsxyLAHsDaL0B5oG25OB
RL4o9vo5W4HPYzK4lfk4F1SwOwryuXKCaiadfrfJPVNxnLC735O5T9FBNRJDmHzM
ZZUVfeKyDkuVE6N4Ywmfqp3ouj/dFnMWxb6uLT3z9fBmGEspVQYA2+zeL4Jhfda7
qzb2rSreUkMm3ZrPFYmM79a2BQUmlrKMB8MpwRL1K4qtYJelfjqpHgrEhSA3JxAB
o1DLJ9wvj9iXXm9Z2FALDQXp8osrsDiGzqJCMej1DEXtqeEoWqtX8zfD+qwYvP7v
4id7no+ltKsg08X+BQVT0j/aNjh6pMn5RwiaDSFU75BRktbxtXJpInfmc/JB3iAE
SIOkfKBDn9E+U4+lvKR6NXmtaNlzfi4qLeHcvamANX3Zej9r3p/RINMXnfQZz/DY
f3d9TTkug9aQSpN5Klic8tz7xOlWm5V8Eov/b9Q4LJWBU04QCyP6kzyrPgG0s+Zs
XE75AyKtrMLNtzXCJFaEwFzVvY+MCxQiaJXyp9l1GntCgy3OIpiBO2GNCg+10WLM
hWnbw12Knay7zfpTQkC4OnXYVtsQo6cDwti1umplAVOFxNy42L9J2oeN23JmIec8
RfRPln0TgVJ/fAIwYXOfjhii7DE4TF/7uK9e7sksFRFCZx65nibZmlWmvQvf8iKH
50HhOdqnh4EoOCg4f2/K4vhSZds+7EQqUyIOC1OI20I6PERueg0rod2oATaA6+Tj
No+n3aVm2JW9+SY4Jbf68Sx9pVlbBM0os21PdrwMxDLJQdYSzqqIJbfolLtdwdAZ
wtNX4TjP7Q4J1e0XFCm/6ng+saIiqlPAsKLPv7oiS/tDxARJCk34/8gikb+26bBO
jhkJZpOfQxeLgvvlvi3yQY4mQFFFOo8PG0vLeaMvoel4cPrXLSYobZtTOCI6baEJ
NG/+w215aOC34pmSuLG3N+z1ZKHn73cyqirPFQr9wvJM/zy4XeAdEEbG+J/I4FS+
pEvKZg1FvJiy+xH9PSKzqWh674ZU7WCAT5FGDcVMXmCnjYF0SHIhX7e6LjXEKd7e
AtmJnAqKrPeZUXh2nNafYoUgoJAuldv0+3pRAYYuQ1jxl2KMg/JHFURELxA/rkhW
g6YZ8L7GU7JCUM9Mv+kR5ybVXD0UVZArxU1WiD86TfiSm+HXkR4cjc0JBXhKpMvA
1aGLO8STV/TEAI+JUjpDv4+yxV5oNVpl7aNsvizyXQY3+l243EKmrrOuId1WGCFS
12yIlVxTm9l82xSatZJq69gI0COXIQgZMDn0NS2dB7KokjdZeQkEN/ag8W+T+y93
5wnTh6TgeT+9Ohmi3o9mHFvV7sc/KFx1IuPnWov8nzoKgm9vzi6tKI2g8F2azkGp
oJjIlaQ90pKwzJ7/PGNdMOqExwq+vO3B8GfPSNOyZac5qytgMEZ1XHkYSLx9Xtah
ZTfeB8jLm9R8fyTUnc0IOr/TDxoog5VWd4dDawWG8vQ2itmKMVeAHAGGZnwb7F0g
x38t6gXu9UfV3VR6VEi5r0HI0GQPV93JBOhopKisDFFdMX7iSB/WuEsXspFIhtZI
DL6jU83eaNt+vd5vyxmYCVBCQOaXD7jv8mw858FnTyyZRp242KbvudFaBA76K6pC
3yEoKIzK50XHCCtjKqIENIyUtmLV76m0F7Sj6lt6S9fejg35Zb+LK9fP6OLPHznE
92OfHrKiQY1x6fIe6zUey58IRv+bya9saFEcxie/34bO+lGrHRsep6K+RdP5CUyT
WziGI1tvw30Z6kjnpoXyPBEZxNIjHyPErQWodjBDzJhJp/9RQUSQsT84gAx089nC
vAwVr/fJ9usjVdIfmugFqaFYnpwo/UPlMUa9rVlxwqfGOhWvhfQPVHvJjHO9onFD
sfxHln+lPF0CTGP8xhSsFOtTa67Y+86f2KSOBhcb+kWBRB/x7BZyml+ZBpxgLtEX
LisbTi2ykWZgzZY9D6IR6WlCv/hf5EEl1ImcdmbdygK9HttDIFvjXez3hzsMUQ+5
W/Oh0eZNXIe22AYcVhThZIjxOpsI3+bp6JyDgVYGbd0FM3eBGlXk9UiPLloJhXNZ
yOWZZTO1X9SRQBVrRpzlPHMBgfWhIYgoy4h2xCaBzd4mflAxavjiJc+uaQgzN9TR
0phMh3802EID5JOYr33XZnelU8xqdjlSDUZ3XejL3971rS6dXGTud/y5eXvgpQuw
/r48Ol8k3cFg8cfoEDeL2P/D2LnbZOlMiZSTYA80xetQlpmrKJgQWQljiUYyHnCE
68u2EYy1aArq5o01K5vvZ8/4rDI3BU3T4YNlMCSK6VxHt+pcIyJ62R3hMJsxHBRW
Mz8uGqjyjP4jgiajaB9tZGFoRqgkRpPhIoxHhFP7nDDX/E3KLWSwgAe11mT7yIKe
roYNUDgWFFBfosLzj60N7lmWAbY0HNnD3fDvHy3oLL55/l925fo7Klau7beM/bsr
yhWbc3t3lvbuwa2u0Sv1NC3V2+kvBJfge+rwqA0wd/CU6yRK3b4Zjxd6KkT2LBDo
K8k7abJc5LkZYDRCRn7tgB+jFsOIfUWHAFIftNJ2e2OqbvIwQuUfFUjF8N8Oakbz
7/GQMavMyc9IC+OlSM1nwozs+7XOYT208ZVvtgVSlWDaPPTyVbnzPro6+3Cj34eR
1xY/m/v0gM/vLuD4alvX0F129gjUOsu16JNYeaRyxkbms6RDqvosY0Y6PlZfkraP
yJGEJ1PwYKiPl+oLxoXfaONxRyrQm2bG8lnrlk7rvy1aFsd4jrfty8LrGVa/PtDu
sCZWtK6qSroaHXXyMEdCuejatKQKde1rpvl6zGLLPBibfibfw7wxqvUHPEArFrfC
fSrngO6Swj0xtj0hFeax/6uLS8BhlqrhepdyxoQEl3YpMIypiaIx7F1m1YMwv1oX
SAmNAAmpGisJJcC4Z+be2r0mqbfn7zPCoYDvhNJMtdXG2KyJsOOKWz4m5p2Crpzb
/fJ4j+DOX82g+OG35LFg3SFixUzKYbOZEAfxVZAAOgCVawCKkyLOrI9Pa4Q8tFkm
HDw2x2WkVtU0cdM8nvbQ8S/ZfcJcT1ZnaM9IYq8NPzI7P47+RciseqM20QdCGdAE
4aTotfT8xCaL037yNKMZjmuUcP6d8y81sivdgyntTJ81fSFxRM8fE5Y5dHlbWZ3Q
LOpee3MfnFnikEDIIeeYLnjmFoZ9GbLRjifaCDNY+0Ve2WbW1diQBdZbOOp+KhmY
tQqLkJKWmrtsdaXxXHmgwPTWwvVvWbCarQXEn+V4JuDe49QSLd5J010SVmUWSXD+
hW6DWOodumn0TrCPCfaomNJZkLA3GA270zNiMNsyxBcj3GymPDqdAaHP5qx63FtJ
jaW/DhIfD2KC13IME6W2F9rcSCb5I6XkGyQIQNYVZxTt3I9DjDgAlGb0EaHEqIWX
HI/LrgkZu3sP2pBVaBQxWOk8gvLm3sK4gLg0KfHBtIPVeQAiOA1Udt0F2NiRsolC
vSoidIlh/f63W9mLQGYEHEYJ+j38hx1m4i3y4PPX/AWikmWFOB6+6U/rBIYaVynw
IijVHzwR7FgkQDnnOy8q2LFe5WT8YXs/+mtWkJVBswDfJKbIpBluizU0WZadlSIb
v7WfuwUdnbjjZm42yWNonBoJSgnErDZ+4YEJpxCQNrph+H2Fmgbv1HSCcUFob9SD
EDthp0jIKWm3g7VOHdiQ9dC6P1hm7H52koOo9Z76fclvYQzs0Wh7+Coa4e+nGHJQ
PlATl9tr1FKaTGRkKC7fagRG7SnuCtFgPp09xbEUBkSv+Jn5WYUqwiMVF4f6ge6i
1SUR1cWYhP0M52p75g7BWMhfwi3TiNTCBEXmdJXdiBdit21vQFV/mhdU/Wn/98EP
f/KVVn7yY9US1wOeuSWWam4lVeo7jpOfz0ycsQ2MpD3Ia9rB1vcq/l1PG2UAgg7n
ECJtQEUCbMpl46XEnjZ0Q99jUGODswCR7a+Zvngfi74KRooF8yvbUlfc3HnK7TE6
AFnvJjPVlfmfkuHN9zRNHbNmb8D8oTuVBJleR+JO9e+7+G6xo+SikSY2AFvnfvz5
ldmWntBuIpI7LiH0s5hsR6A8OW8wjSq/8TG+KEtlRLnUIxUN8J/MDkdzKeNiUpGe
XxI17PNfmfcHU/yqRq41aCsOQr5BVhxzlxAh4l2ck1uxrLarSq7tY9w8W3Repqp8
zlfMuX72oecyDA5BpfV/z33FlBDO6eVPCZUGq1rIb0r4A9xSEsy92MZf2mwW75/K
yy+il9QqmP0opmEOGFkT/6EK8WFianxG7WHkfUwKhlP5GdbexRuvTAUYZlDeAMe2
x5kplqDch414n4MbMNetq2x7M83xpNp40x5tx5in66LCdHT4VC+AqA/7uq9aJQA1
+aYfIUNZQJqirh1GnxtZjfLTlmaxQMfo0O/6CriekazNviFIhXzF0kXYYzgdK+pb
hqjaTuQLjOCkIwTowiUSs7S3U+MmcAvlm+AZMmJWctvZmtp9QvKzU4A4YrozZPsi
6h8Pc8p2o2SLRx/OPfHJ8YNELMKV8SotBnB8/frn7PIa7ubFI7ZqC9L3/pleyy2D
oWB+QFj7bZEg/QdERilIsdMwrYkXLX5lTXj2f8yvdl8ioUONzwPvfG2a23uONrAp
znFQ+jQg5kzQ8xx9a6H6NOhdpGIeqDvTN282J5Axka/IaMT6HOMdXEsoV52dhcVQ
9YbPekYIczyeusT/LkTtpK7ytn8ks/OzdykYegR0r8pP1xAOHTi5wEkGMirhMb4U
tAPviTNiE+enJ0rtiw9MS1OPU1vVzJnkuzR5K4a14kWqxa+l3QNIHDbFWXQPCUZV
fizvuPb2kdMh9Lcw3zh3FxTNyTN+NYuIUz7v/XsdzUA5TF9hF8CEv5anYwokxqVh
cyXxwFkYv8EazmskJ5lWziZql00G5x/Z8WL2dGz6KSSniOc+Gkd0KJ8VfxGMoYOK
ikF8YO06nI1qFkSb0uNB6okN3CkNMVO2BkxKW5+Jkr0RaMNkYHa+vV8Q+oG+fGWI
ttLlBlb1bxsFBPezReg1VmrsmZzGxmJZ3xpfV2GuNrL+/VeFL4cDvTzBjcp+2P9e
8JkfBJ4QWiZNDJC9Vs2vQzs+8GqgAqvxKdSpTqOrrw68MgOhxHTm87D77oom6E1h
oBQm/SQ/jeG2YQUjG3eYgBStzDZj0itdnYUQCg1y+QAyP43GlCLlh2+4Wbaq51xX
9PXi92X2UMKdWt7y/LjKBvbw1proveb6UhAbxGkT4BAgEKXpj8CJXazzsXM+iAOg
c6TxEK+u1er6bXy2hmyn0jQYpVcBT+gUemnLVgqGfJuh9p3TvPJVmU3qhuyZcP/h
HdNgy40CP/b59RIuc9TjM4jP0KfnmM8EP3DU15wzp5fhLTNYsizHs0ROs3s4CSBh
vADS+xpgaO5gkNM2BtX6MJ/TG/Y7SsrqycSdHSMgafdN4ybGZVR3VsmqM17JA2DS
2g2j2Bt+IYSrq1+vcpDyhl1l0LGq5U11P6mQB5mfT+Dpxf/fm4zuYEPn7nD4URLd
UDAPwtpG7St/dAhLwL1eF11xRs+WcJtcYYJx2knmTpT5xir5fEQCm58No8XvKBh5
5X80E6exDau8pOcU2u+znGoLrIRRgEWZ6KACECYchuV9MB0yboSadSqp+ro6nX9/
jKVcPa+4iPbEyL8NCD/0tW7A0PYnctYSvwzp1LXVvzKm+93zD1DPxauav8YxpnwP
bmOvzqTSmcO0gqDdo9D2x0G4K6YnO0khtGoAMgu7mLTVD2eM4lEJdH6bFVy2/LNp
KA/vmMoqLr4uhF3M2VHMdFfTorwiTBauTwXLh0OKMzhHHFZ8xYZaAzeidBwK8/8D
NoDWv8II/MzHokDCIGi2GhUTFauKKNzDhAdBYLR708TGZ03HTI5l26NCkLRcaJyb
h/xD6UpuH/z/SMLQJF/6RuRyGhmsytORPbya25Q9d3phKS71m9kG/viOvfVyMW22
rRA+M/qGXFBgRTDiqt79LDSQIPhhfqvzlPss+gD6PbHigz3uEKH2gd5mPLOUvHWu
V94dndF+adQBx5UZ57KGmBqpPkYo3488UpRfsRdHoFgRgA+TsYf+QPYizuo62J+o
xHmwA5ao384ObpXR8z0ZlVBQ9y7Vtfi3ZWcDrzUs2tHRWfEpnXsHuZHjbqCCzYcD
domCDyobcEg4+k/VRnvLprCelr0uxen+LaDg4iCuyR1C0PBl+xONZYuU6vsgDMZ0
jv1D+uc7hD74/Ma7SakNwAtV5k4EHpGcjs+DTbOvEiLOen27HTQIL+PDvD5hdCU1
n4EcQF0r/g2qKF3nntwfPSJzX18A1vhEJpQpRcJGk8AwB/ssPXfkWZkiYGQZYDi3
g1EO4XRpvAZtl41fgoeVYXJS7VEYl1oSaOgPylEZh3gCNEON5ghMjNu5xRfFet81
NxqgPj9nnx+ODjeYBW8BxUw2eQDs8vcYPq8gIei0HA9DUIje0Qdhdi9n1jseztdF
0UUcPx++UyPmaKmaLxULCGWjBZIWh4X2x/Q8xwwKH2Ndu9678jww4FIL8/yPXE5I
9ww3KBjcSKwUyOVzt/v2R58cRJCWMVADbG6BL7W6+8bwiMnjXa0PJVRXL+KV56kR
WII/LfGQR1lJrclrxiaOe6LCCsYEKBoClGgUouWukC4syNwkVG+GnTEpH35g1uOH
DvSvWbd+qyicqzXNNikUVkTHVjopxxH/UV5tVP3kNPP+U34dg7NzlV8W3U0sjT7E
D0rmXLvmPsaHOcVCqDexwDmI2f5+/HNR0Xz0ZNNg+hXY0tV36DDaQsY6ZAx0peCA
7Rx+4xHoQDz5FVV0MUm4JiLi1EWCeRR2KbLqQW2oa6Ifa79PzNstFrJKV/e0WwDv
9dJSICUKTzeBvCUcnMdzQZjqTmY8OELy+LdEm7dNmO2vPS9vSXa013uBtObUn9nk
MVuUHVA7K3GQpZLcMUEX7jkga+QqxWjf2NNd1dbZL7kAUDTsHtNnmP37pMtMMV0o
su+J5EBiScO/iaBaMCRSJkIjJK2GfuOSLhIdGV7wMIwq20b4f7ob11nOIaAW2QTj
bNjN/xk5xipMG5h7MOKYMQV151WswLgR2cPd9eVY7j+rV0+C2X2YozY34DxWXE8F
QCtV9S+Wt9mrtHXqD00yqBK1fSS2e+iOorJyrscgzREc6kZ5Bz6//hVv0jyzZGOe
9b7rXKCNKEdGi4F9++jpcC1lA9eSUAp5sazAH0B2aVv9RiuvXjk+eqlyAVXycQo7
TghKcAC7NWubGajIo18hzpfPCnCiiiutlBV5Pz6WM8kdPyaUntW8VUch0O887ZR6
fmmOiEvIoyN9kJ8NDPdfiJDvPD+337Rin/y/qTszBxM6EHJkXjZEtiI/THcF/piN
Sksqh5+Lppt2rkL1VBTsk28WuafXXz1egEt3VGQ23gs1UTZJw4uH5nlDJ25Z0vij
ExUTxBbcXZsCnr7Bo3nPpVA1RKZ+3gGRcS0OozcFuL3A7I+U1uVjC6dgV0CsiGle
LWNFfswbHS+JACZPfOzixy5fap3BkPn5xIA6vMAD2K0DlnrhSC2tEWWavGrUY4au
E8bJGG+IqgzBKAYnj/L/QmwBGO83PWcKwN/Omh+euteoktwSybrfsKyjLyrCqqQD
S47dPC2dlzJzICPzGsLz7p1P01hbJKHoA1z4HJhb/eSBMhGOZ/p/YeYDeCNq8U5h
IlI8zbLCRwUUx0pSq16qnN99XGRfAs5JKkubnq3mMySjmSiBO+APaGTehjKrNPvy
fur38bcjjDKTJhZD644ZJqCemjbygieHadE/1gUbTE8kLcK74yAULv0UJTRUSBau
uRZrWb1ZJPgia+b3QuqKrXx9c9yYGFAwrFYMDas7yT+mIRsHkoI73mxXk5kC0a13
8C++f4ALKBEeutt63HRyEaGY+qOkYP+X7jNOcqIHcPiJaYTBhvAxFcRgeo00dNhm
BqS2gJxBxNS+zS56YEdXD4Q8ZfNBYM8C5X5jzTMaUUsTaCW0aLzvDy3iFVzEQvjV
KvFIhcS4ZWrKBXIzhRzv9UpS24kb+wbOU1E0+0n+lG0K0Sb3xKznYUlwfBj/eCcH
eFQ/40vLlKDdb6p+F8dZYIyXZn2CprUfHcJE8A8F4Abioomu5foyK187X5woThMk
awFRCodhNpZ71N01rHBEJHg8y/KoGiVZnlZ0E6Io0UF/qAFd0WigdoP/pYejQBJK
k226Ytne8YQ9rUNc9ubtClAniHBZYViwP2qopnZcatB0gEBRSD3nnFdSe7tXUoVi
2RaTLBemMH+2S2Um9arVWQtJNK3TSFMAc13hCP1l5oVPsoUYvdpM5jgj9IKG4QPo
l2egTyHGOzO1wlc1JBpAJCIhvgGB+Yp7hAMWPFeIaNCCdP3g9fD6/DnVh2DdbICL
Rn/fAnqO5eBDRKwg+KtqQBTsDEYr+MBzjXKDM5ey2R/v/Y+1zU3XnRuRWWolutiH
OodAJml5UpNk0J0FteSv7GTiXJewxE5ajzAYcVngoHreDQVHgbzAVI1oSh+ig2A6
sNltH5x2RJo8kcApplMUtiEwirkvNNeuG9MhBrIZX43OPpodZpcpd9rGUUranvs7
wiwhOKQ4Nct8t9bu2+drtCBV6s814L6sL7HqOBZ74WvdH/TcPwdeDVzcDPrV62rP
AFpb9rESHNG655ewq8OC1niYC2DbbXAVmgbMiFZtCd/0bJZh3sXbTS0Uj2Rim+Nk
pAVhXibRVAfqJvbzPuz3qj0bbUsVjpbmZmFFsFaZeKRDC87y/5pV8MOLqu0S9H+D
o64XC/UXrpw07kfdvCqsVeykPoqMsiNBOGJfmjPH06pkEvUnKj4Ch8uDpiEnpDPp
rD1kg9cJwD3arL+9d6TxDDgbA+vtnyO0/LD6gyj79zfVh4vuolkZkGQ4OBFu3INg
GUABf9y0QXu+xbFz9VjSmVLH8H8c58DetTl1NAQz7lgR3yIVKk+j8YgKGTv5jTJl
TNufzh5ctlBm6tnbNHqDC9ZIy8IxYGGlAGrf2Dd1kScc4neT01aWDWuQaY8U+/Vy
1lDge7EWzTUVkm/h+QAu0BVcHOAT3SMYv/FTvmUrtPB9P8eqc7ayWD6/MKWrdCVB
6eTsg0ZlW/Hcwf8STd8XAQl0s2grzLDDfZnYJejPepnNRJMRlXSw+wnodHLwRErM
s9DFKhapKWcp15tPuecvDn9a9wHNEj+P7gFDuDVqzamsyWGI08FoM+Rd8fkGDShf
MS9xqltslKEqHA3Olw/yrvZc/KNx0Vq/07beupRqccw5GtEbVjave0dGZrGjTJzs
78FadoP4FmOzPYWOu7MJA1AA792e1pmkhFYMm9AM862In2FKbFZd7hX+GJbKrvTg
AcCxAiT2Z+3+RdHozlaa+FNhvi2L24fEkMn7wV4SVn3FtDGUB55cdAvvQajzeC7B
cXkS6Q5u5h1SpjE7TKkUuj0LxJTrRP90H6totUt0wrZkQ84QEj+LQ0+4eGmC5+lr
bSPLYzZ7Z/bVh7vmDHuTDOWvxZ83z3FkaYzcF2G6b+Gc7U0/6CqR9YeF8NIoZAPL
R6baHV4Pk8PtppeIHQCiNLSs7g8/s27cO3efnl6YOKVSwVFwh7LbEyxU4SwseZUw
4mSScyZg8kZKgoh5wloPndq8KqNw8+Dci339d3wkUGziBi2NjDslGFbn5B2Z9nIT
Yir31+dKRVCrj0wb5NH+BwamR5wuJYu6CzsmQgVHy3y2M8lioCk5KQ7hqIj3h+m2
9ynjGnWql42cOoIHZgaTXd4GYAZLffDQ8zQv8GMkHplnXc4jt4QFMteMmk5ktx7T
Ryr1ZTzJaZD2BUQuVEkMIrI9nEfFO8hDxsRILSmU/TGHuGIXdmSlRFAmge1RQHHt
pKGBR//bebU72AzdZYw/uGnkQvxWu2C/I0XN2s4JEjKcJg4aVP/U3WsyN2hi4iJT
fTJq+NChoZS5jEyIX6KHo3/VjfzzABAfBHaEJBP2cs+0jte549qT8/x9s8BfIzc3
PZtBe1Lsr8HvlCL1pyRVz4FvjJ+RuRdFEGbCJ+bNp+eq7O6Nhlp6TvnRqMj0SA/U
/su3Aea+pDSTNGye02VkpRUAiOSicRdS4d6B5e1FA/VI6+ij1cdIRNwON6YK7Th3
9P5MIhIkFg4qi/vT2vJQsZ2JI7JhupN/SYuJB33SeHwyx4z94NX88dbrekPQsPuB
U6tG2j/GCOhPzEPXOyiU1aXiPfx6w1E++Smjxqm3BDP3hF5xZA1C2wK60iBwBrDE
RMIODXY8v3VVlQaol5XEDnj2FQn2JHpoxkNglYUcOaYvsDG5hprHfBg9FZYEPYSi
UGDg81G/IV73tRZwFMdlwEwwAd1WYD+B+0I6zgd/HcqnOSzf46iEteSpqBbzO2Lu
2xx2aTcbxim7C4gWVQCPwntgl5ey4ACNJ13gmwAs/rRAOSLAjvdJFf/+4Ua4AxbE
fYsfnHTrROPXIxkJONRWwF4x01ak9KmBw6zD02rbBYXeICsUpTumBQAY4hiyeqMD
BB7lryURIXRICf7638161qeeL8oX4kyxcqEKJm96BK7Ryhx12hiywrVcXHEiKV4r
zGNezzpmMYfCp1uxCqATs/EZxEhRcMKsCJeGy+fSSV83M+45HDUM0Vqvj+OWt4v6
l8EjZZiW9EAH57CVo1WpYe9scS1+/YxR12Ii04Q7dnuE00oKDJ1MKvy5s4VTkky9
RDninGBuwoU9wrNnAKm64OV9iLU04g4ITWh45hyqnjQbKYDYtiYPKG5ECyzAvY2V
JSebJPRTNsZxDk8rwV4VE+mOHs4LIZ+DwFQubzesFp3JRQBkaUU5CHSyjh2j85y8
h7rFZOGCEtEQx8ovqQ8ut7HurowE3H4CF5VaTbhjvZ0pIwRxUSXaEDOJU1yuZIG5
71h9APG2vIbfYFCpMnS37TEVt31239HKK1c3+rCHa5UDLGGz4aJYyumnRFNl+/mL
EJI+wpisgvpkJbC7LKLPETt6tIsarCSbyNhUkfLvsXjG/hoc5YGBqqlyVOhfJ7t9
IQM/57VI6QKMP55fmRTx7SrC4nlAcyT1LxyU/xe5bDQtT3cBVDXk5XMKgRM5RI7C
gh8ariQS6zPAVO6BSNc4Stfww1QT90GsRiIS9fRuvBma6cKh2h9EI9ckTR6shWhY
+DSNgx4ugaxLaB977qou7PD3c9mvHS/mylFO1sjLCh+r1xl4SypnrIBw3mAreYsM
5kEjb6G5P7luW2FLfeR+PV7sHGhjY51Zvfn2Gqh761BBu72+ong74/Y89rtp1fg5
4qRwpXJ28b9M46VENHEvjP4bkGdma8CfhaK5IydwV7+fsgS/S6ZniCl1CNvOWlel
tSiSXTdaisoqMOPCm9GXsGzMAK5u1wVZDWWukT0g8yiBft0pMt8jeGo3Ee8QviLV
ajSMJ6AumDZW+wWf/ae2JgFNL4brhjP8+UQKFQjoiy4WHXgB1rKoUv8NKQVkaFhd
X6Ah8C5eoFhj8Ll9X0G0EjouQfum4psJU97bEvyR4eNcPR8pUT4cc3c+rpL5ltpq
nN2DYsiO0HuyXjm+tHNrvtmcwZprsrkWnqSjAPz9kktwn+xME5p3LkbThzq9d8cA
gDzCoBN5b3xTSTMBEPuwWbKmDI+3SdDOePO9ZV2fAVC84SJhEs2lnAmWGWbz9aPV
AtUEq3UEK2Sh03LdAKY6rwRpiZ3xuAWVaXqLg8kERNx3+aL+pKDvgBK/BWDafiXk
aVV8cWygV8gqvoj8Fy2wO0k1W6hLEDK+Df9TWld94tw9Mt85VG/6XE4AFft9OoOk
1SrBVV4QRs3yhpZY8iDCrijdaTymEogz10rc9kiyIp0TVnkYx1UYTo2fCwj9y26I
CesH7DpLS4SCyM6CjOS06mhHAXm3070R10rgwuQQusgfAhEg5agS9ON72jw/3m5y
eKnJ5osjgffRYyvkGaXJ3ZvgklS/zfQwHnbExbKnQK4VIvLyKp5e94K/T7yJFpy3
wP/Blc/VvS3x97KQTRgEHXjVM3rgNbr0ktCXNmxdAdIwRg1oac3dA/ghDtOJRtwX
8CPl0QRdboU/17ErpmX+s7d3CNM2TYEy/cfcfIamZNMO6BQiYHI0ZHxu5iqpUtSt
Ijlq72yCAJNM7LTmNLbmxV+zUa0sr0E/7cQZrTLyJhYQxjIR4TyYNYZa6Yr++tvY
Ynfct+n5qIV6Ki0Qku1r60hVfrU0eEMftW4TrrYHDMOJ/AFOdyIdzweiPRgTWlXx
6yJjGhVFWIpI4wj9PIcyeWGlfTJSznKdCnCYrl1aVCcR4IdwghbhJ8HgX5rp6v7R
XztsPqXR8nTFhcYFUXdPULnm+tbNh6PS/6vUmdxeJ8Zbdvb/e7jwpK6063oPNPsP
WmY8Gf5n22Lg9q86ToExwQuzmLIZHkZRM/KanPuuXScbVBJJCSiH4ELbaSFHCHdG
WFDiyIcjs0ta5bs7KwYNfekuBbEh2NvqQmLv0u5DqSSGQxFWg0S125y6m0Sn1RGA
0haar4U90wQPeiN4+Zp4Q1b4FbLrIiFpNvF47n9fqVOImpt09wn36fCg7nkBe8aW
I8EQHEcqz/xj+JQL9d9qtKFOk8MXXoLqAihZgvTV4p0B+IXlfJDjsN634tvokf4H
Zm3CCNLauvCQC0C51SGC6yEW5qNeTktBr2Sc8yAnK1RuELVo3wf+QNuZvXlS6VBQ
Uftt4x7nctGRx6DseHuJkMF0fi4JU4hcRZUL70kqg8Ww41NoUo/IBxSe+ygiILVe
NUjajpX/ggdHFEPbV+v3xoaXdfk/fP/wDD6SvI1Rwlm6oRGMl/1j/vunWH8cL2EV
CNmCeEoti9qvsrYBjQETJAKPeQNUiHNIOzkW+umIOhsYBTB9158hKxcUoe4w++Pv
y/mi+QPWMfuo7ziGaJUoB9FD4WDrxEgWnJz40IFeNq7Zfy/cONNRqA/6ittUP7l8
hpg5rI+LLd7VzNCin7ymQrG4MPhCUVXtrBtgHlHxxtpM84JN6zzTkh8qsbYJJY6N
UcFlypscIHRyYjjpLZfqRDHZqhwrfCPkEx/W/Srzw/ShhO/v8TjhWb3LQMPbq+i/
2VaOAd4/zSK3WHW6EPMbExrdSE5K1oOxN0dZMTjCiP5AOoyrCm/Hbk+PcgwopEhq
vXvznJ5C0prKNkiM7nFEzRUaRDVzfLtE2p23+ZQZ9AA1MIHQkTfULbSyR7f3Llsl
/GNbkh861m9ZxD7qyy9rmWwjcszIyqSphoCBfaR994OWdIMWW0rAHIUmIs5Jz8a8
Ijn26PXt4odhe89o2BhhByc/Mw32WYi77EDu5B0DN8+OcCb86qk57eE8sy89rBFb
HuC+5SHOdcbRq+yMW0Rlj8LFbPOox9NYHFXU25Rtl37CZh2vDndepIsjj9ckiRvj
rq57On9/PB1OxB7WL1enTX18XZdk3PDVU+C8cVeTZbYVt3XH/cMB4CAGdAqwuuMs
SBcNM+ITa2RjfYWrTO1QpL/rjYuowpe79r1/HOF71cBn/f5BAfFmA8Fl/UrIXFHv
Az3ZSD8dgE1v3ngNAngQ5fmg8UEu89y3zdroow86V0ZgLWG8myCJIZgJ463YWabV
ZgTWSZWEntniOTuXLOWyg3xRFJw7PSyVtaCw3ySKZsM/kvflGd0+2LCmifn8VL3a
+seb5HXNuOCxDgMdaMweHt/3FMFQUBQUceFmrgdf/+bd4IIYVO7OrlvCdONQmj+1
1TBLBTrTC2qzheJRE0GZUHTmj6UwdGht6XpseJChS9F+f4Qt2GAkEFFh/CUKhLkk
XCwZhNe08QNYWWIBFGUffayGcbMODMd9SNlPubh3W2sCsBXm1CN6EoOWqbEalPOY
RQsrtfu60KyuKU5lNZnFV14wHYnSo/pjbbuLbIt93O/zfJneX4H7H1qFzJV3HN3e
b1/zdJ+MBFfRjjHehxGLgjP6UEAJPPiQ06w+QDE59fDm3uZX91jPV8hNBx12tQ3a
wUeSHYJU5PqPAOe8gspnv0Vs6kFf+xsIE7pBm/6UAAoH1sVjtwN5/KeOiia55PJv
vB5pROeq9AbLlrHipwOOtciYdDQ4gJAypZe8hKtMv543YMIALH3soPV+6GLBv1rL
SpjYebZTeIIJWHscv6/En21Z/vbjM87NsXIASiTzinIcjcN9BwGKyETihWrBg9j3
swceFDvB3r95kPoR4SqOwZoLy1D5SOIoBTD1q7iA8MZiLrQUGbUPWkD+lTfTxvpE
lTxs6YEk83gXZ8iI9FBugbzimIZYDwrJWXmJxsePD22u++3GP/DIaL4O8Dthu2EQ
FgwXoFVqzGXoFcokiLQVVJ6Id2kFuWvCaZV5xE1dDqIGuPEtPTSpAIWwkzcPmRTY
u853hrAqdd1Dc2zVsJ9e7NIwRG0OnmrmsWHLP/8t0QVT6Cyu7LOyIoQVsxlZ9VuF
dLHUCFtuNPJvOlvVKRE0S/h1qcVUNWfwFxFu2G5/KVCSxmST9F2dREtPLWFwB9I6
ImNa3HyVxFu0/57KThRbPoLV8JymYoRSgaIwxox/WJlttDWT45BljfxKEJnMA6pJ
qhfy4KyKMToGTLQxt7LIxxZzG501751BjpPEpUjV6k8w1vqRmJZQFr7CybL3Cxmu
wXuUCOMrvfjGb8z1BmgEpicPIvR9zCmO062zbJQjGpKqxqHUvMZijTCl3rnI6RRB
YsQTXY8jwIXg9Qmn03pIlE0+QX4BwPnSZav8dqVBRdn2O3eYICRA/5yIEDO7HTPT
jTJbDMFhvwwexhm2rVUBh43fThP0CLIdBo3zv3wOBlDOzlwmbkV57LiZ1zrF6+7N
L2M4du2k2QixZIOXbrG+HWvNENUzCkBV9otDMSyoCEfhC4O6rLANN9uoYE8ASjtc
ayHFP2UvZ+646FYa9qsRgDO/GnneIyU4HhUaLh27L0ObruD2X1ssmjRp72Nmivo7
GOJaTUvV8SvYE6jc0alajypjhaQ7CEq0feyJ+Q/KvGuWRglMjJg4ZVd4qIc60/k3
ZsznktvXAoXrk9OKVcuz49zDQjP/nNs2XNwYqT2i1pZTWaNketJbJRGMzgIfHTCi
9ZRMFdS3o+fW864mWRgVzAVfLR+v72AJAe5tJ2q/f+n530BzBQrqa7rkb9NlzOTR
VI5A8jTzbvlDaYGgmgixifvgEw+kY+flYEPT9ol7eD2arEalPYOpude4KJ6fYQ7z
b2mt0FPkfvlTiLOA2f/URmRl86pp8WHanR6HmbsOEAHHURUdl5sfcgJdsyrxhGv3
Ie5OYOS59BEKbJETmYlaP9YFulLoOsH66Pn4ScfSdDIlIXEsQLd4ELl66LfWkYQH
1juo4F5LzyVtBYsvs4xT2ggKvjajvkRSbzomXJeF/7+WzU7lg/bF3l6nN32q8e0a
4dMSVlzQqER/slfNDOhh+46Q9CA4Z8frmxaKgVAYoKpXKjy0nySRE+0oFqiPZV4k
E5VXUJ3HGYYy6C8YD9fgooQibnAOfezMwEDk63teFnZ8HvWxFeomBqRa3vefGuFU
MiWsjOE91SPYWYAwixD1qgD66B50sk8rvjhUCaJ98LbIHcZS6F9yF48pa9Tk/2gF
bLg5a3vGcO2oB9+wXvufyBZixq1GDeg6Q0TXFD0zejTVUfDBQ0/ebgNRqj3OUwQm
MOHcXi/39qQ+HtbxuweJRuJ6tm4mc3mn4B1ftQRqpwvYqml/A2YqvpEQx4cXq1Ad
bRXP/noKl3iq0+Gmran423Scv+Q8j4NMZeOsk0tAsBf4ZEPJFZbT3iP/sN/oYDKW
f/dF3igJM8ls8GtIypks9WjWLDdK8dajyQ4312fL47Di7DKYL0Qw+uPSCJr0DcrI
y19FRSbgwGyxpOPYCov41XMSNzOHxUuRrYuTdmpkKxclkh0//39wOLrIvlpwb9eW
FwquuL0d96BO4cyRJxzFKXGC4HmZpfmwRO2DtkNWf1q9ViHkfxg6IULuhUkPDzHd
aL5aNuRBLr8gqsnBbX6hNBrCNXyKRuEbkJZZueJR9HD6UxACXFQ/YtAl8s6mB3yV
W8E4m7w2B+fDq5/AIU79V/qrLDTwygIBL42rS8I9v2Zr+ZIkBJQCwFRDNAodjJpt
mtf1LINO5Yv5KiC+1TzJUwdp+Sx17r19M49glsNygO67VxQ+bWYAHlsSwamf140r
q6chClRX3c8fWYOzmXNZPMa37bxxgz9C10RWETzKRAWG7iDJ+SAdIJzDjpZf/0U4
HTiU0aiReiJCzT+k2JikFL6OsuO8bqUKOS0XfGZati+VVaaxEL2TuJxvuvg2vTVF
5Xsc2//br1WRW6ujMBZYs9IBNQOg6Pcw/WxRPlS272K98WQEAZGVVUEXeO370QlM
kF/KxNy4chPPMRyhtfXGU6hMkTaickOcvvHWrF+W3e1Ka3eLYq7bvgEJVw0UpBtF
H79CwxDsrC5UK7tusunfiVUG+gpZQcRLcqlrC3Y+Upzx+cMT04bNXrFKGBl1ivUB
9p+cu82SVhdAZCOHjiTIjf1BOLLVAvH0s9rcT5FKb6FdUIda76pZf62HBzu4Hpn2
jeJDwg6GPUeicT4SLjkhLZOVJ80H2oD5hNwGnW6rYvq/l7TbgQ4XL9ys3lQoZuMq
WVj7YezL2NvoH6pDgipx4h1DcYspTS3qilYoPGTNVdDa6wailCT+7o7KiAf1GNq8
om5myQ2jRIgUNP5/XeHrsCqec8pdp949jWj4VyQhwxTiqjLiYaOA3Jb3Ckte4bD3
4wKgg0ukdke4Dun7kxMXa/kzQfrk/8eL3PchDkJ3oOCnrjscO6elDXXXHjurgQFU
NHuLV+gaPYHQH9JXF4PamP3Bwkayg9AdwHVYoBHn8PtQcf1xhmL6Ls6QqLqiQfdf
6/YFkSpxrnA+hEsiqTWihhvGtMfAmKSfkuXUpZ20L5SockTIXatnhNumBXM8p0eI
fMM4f2x3z5O84xAfWg0N3oMqOZaFs+FVZ54NxBA12u8/txnR3OY8YSIDy2AjNuVs
jXR204hkZM+oi6leAUWjTrk4CFwvb1pnZKODEWxfPSKWn/rb7RB6YJMZZnc8bMFx
Ay/62idc3dLcuFo2czVFaoVi8yyjhl+4LoaZzBW4eFEpKln7xujsU9yX+q2cxPDc
Wrm21GflJ2nKIlmQmewnfq0P8ICVU62FSgvICdKgqkO0dT59v2sNByPaiz9+lxMy
vOyGCXXkQv9+5/5PjIE4oG5Arm/GMH0+rSG2d2vykr+Fa8JrS+FvwMhJpDgkLU4X
mqZ50My465EUz51zpE62ALB7IMxQ02r2ei+Gqkv/ofg2bmQp9sEBp6cuz5yoFRd/
iJZ2dZF9KCVceQiGMtjD+okJXd8H0x683sV82s/MA2JfFoInwFsp0E9+KEnu5+O2
KzCWaiJ0SPw1PpLNvYjP5XRYReikGPOaWWb93GhJV2cdKRgNKdLvqLVDC2U93MR6
cWKB9Jqbp/zBGorEJP3lX2w3OFXg+c8hZwp1N0U/ugV6fdLMvX3Y2mhza6MtenkR
GC8f/Z/4n6D1/u74IrURmKtT7gi7PXkPBTzazFHxMkJaZ/B5j5KbAHkadlx+ioPQ
M594NBRCyPtCT2yAar7lNgsykkQtyzUCvDNSOTwE2zquSVDlRr6O99N8P66SCavq
3FoHG9S+62m/JRY4nD1Bu9PQ4+Le5XA/El9UOVFoEpFzthTWNIivukqGv8JfJsbH
V9w6/u2VYr88A5ntEwy3y5PjR7ZZXwf+gRlQGMGNzQfgahgSdtHrym6Sxnv0GkZa
7sn8t3TRjdYznAcXqg1kZh0o/CKR6XAj9Gvo5ZNESK0TqpmfAOeYP5Jc0yq63hjm
qQ9wohHAEVHRl4vX7EJ7ui9id28mhi9UzDisbwe/0jR9yUg0INE7xBvE7YfeKa+J
Ni+0jYc63xQ4tGdxmnUoviwqQIa/SzsiR+TJ49HzFcOtnZjph8hcVC668h14+w1K
YjV4WckWPxp6GUcGDTEvEJDCvcaEU0sa4y+n2JP8u4RLKlj3CsWkV+QgpnNXEapp
0iFhkRI5xBGMnW55f91bGUhaGi6JOBLdUWVdxnZWBtX50+uaB2uSOjptYQaCYFYx
nENTEPm9bUCJgvws2upE3mLWQEH22+evqZIjvgaUOgs+3E31VjP6P4r4nn8iY2z0
gX5BXE2FiQpP96XEBr0NMxmnLmYfULaJMmWwBVMIAnG3Y5i7IFY/adSEbc8+fjgQ
i32n2lP4VS12ymCAHEGX2Ah++Fib6eBr/ceLfTZFyOefSQ36xXt9X1ic0XBtJpM2
KcH8X36fHzy8Y9rBlLy6eABzzH6fz89ZvsLc3/SiGa02Qqh5fsQJzVZFNJTP0xHR
rzH1BaffRZ8qdLk/Q82piXSGKSX9DXFLBicSNt61TPRv10URAUR5Arb44GJq6FCz
J0DtqC1fCcSCiOTspMXuGmFmqPEVmuO1mh/ejsaclnndVn+24n+IeUldml8/OA2E
E/zuiGG2O2eM0L9T8o60phZuGQw16MOrhaRNXUBHGFc/b1WHdmKkUQ+vYqSEYTrF
52aSjPxUlXkEflz5Y9E+YH1q/Olt8+7qB6/TyzZC5nIs94nbok/BlwqscEfpACSl
db0Hf7w0IuVY3reQsq1wwmz8GpY43z77PoLqj57iH6nIrQqplptmWuzPTjlv8Jf0
NF5Qkt968BvVxtpUMzXQd2xVXpin2c2w8fKjB4WsZFXt2sNKnCtjKyKbFjy8Y9ui
1MeLU5Phwfa/3SdcweaUJmfhK0KvcGBH3GIRcoUtf/wW2xpTpImYgkarqVHlU9k8
Sk0A5lUEOIS6XV0+NCQXwHze4VcI9xJrQcNiLLjh4Gqg53BJ6hA2Rya9jYNtAZN3
cIVpHAE1psUbeLXEfoFUl0LU9KV4hY8m+veI0p9Uuhz9ZolPbi9QFONl8WRuIVLH
5LMmXyXEa7NIY6R+d5tVZTpR2lLvutflKtCVuaKausTjLRyPzXuZ2qH3Dki8zD+M
knmbKqDCkldPeaSBZhWUazulwOzEMDK7u++EdCztgNFuBYEWS6q9V1wlMR7P7SIk
w1kyjj8PwsuM5qpyoMub58GG0d9IaQLQV6ltvI1xmc7BbG56FYWmsmKWHcZV8Y1p
zdlUxveqQDuA8m7sCILKL48jWynENJW+sRsDl8quuyyCKgFBUEPWhN7WXE+PhSLw
R4YuTga5FQ5I/4614l+9l3Zi6hfAy2wdJnwjzAL6lOApy/i1tMb3e1iOrlwH4ssG
gVOPE0oZQd1LFFJZoZf1pvujW3R7KZx/8Ye8iWMFl4ZDC8EyqxTkTkPgygvSvzap
kyDTqFhQKPJdjni0289TT8PWsLUTozGlio7CY6t4WBAhGOq8VS7bPQnS+u5awpZc
8tv9pwqPL2ZLISjYrFtZiwMQoNtEhTHHTk5TtYgy0Cm8thd+Q8M8GSNEgXHfPrVq
+bXua7XctlN9HRw8OsAo5lsRwRjsuvo8t/vQbHkxeqi29wUF1xE1GTg+4KY+3Zlu
DUlAwmvfx+OScrB02TNaCiL8V3HZclFwdrMrY+TofYwnIjG8z/Yj3OqfTg8Ux65Q
jRJa2B6AfGoTU0MTb+JiGShbAMMeJ9VW/L+5ZGr1XHqejZeKVmnxLVDaBP/ijy3y
rA9Oj7d3CsJlPaAbHZZ8sKNNidrQhcgTGUo6OzV2bJ6cbIkCRR/LMLnL3xSJHAR7
jWhivWkNMQ7iZ5HaR/zy9m3mawY7cIvoAqNNTkEAIaippZSy/Dq3vWGZ9jA4ZTMg
opPav1vvIW7uZ+5qB/sE0LhUhndP5d3NZZRRU7DtU5MlcgDnRCXzTk7UUQXDP9KV
jf87dzAX8WWJOOj9cmE/62F2K5OrSxQkxVXA42qlDvtIfKgghsNWBBiZ1M8MGGgw
KVdjA3Hx6ab6SJ3T8d0eysU561dTxpXoQ3JzMfm16bsyX1GNqmwzGFwqECcVtjNK
SqIWCMH5Nr6Hw3s9Luw9BHOoLPcdpD47ibP7LjyyNrdmFZWWZRf8+e4H3UlCnQWZ
VY5QkQ/rgJN9whBhrKrKEZYdX25hY2IyLfNwVOp72xuta3bDN7PQap3f5pLUQ41m
UlCzbQp+bq8D2fVw8j5MISK9ZO9aPIcLEvmTrZxtjwl8H99R/G2ArDpgBIIf6HZ+
XPU++UioRTK1CnHBCQsE8q6IexKkTpZjh5eXnbNtrzDUI0XBHcJCyvGE4rl6ZCG8
yZ5w5PsMaceyJe+ktzwGqAdwryImojY+ndcSDN6t3F1uOXY2QaOUCeLbniH77eV0
C6yOxVJRlgtrFMgPPGEtGtoYMCoshpfUuzBDR9+iuser6CwhuYEmU/eIMsRCBjLO
ayJqLnctQsApMyWPd6rIsstOEHFOsZy0/DKWX8j8B58/WD6IjiUWZoHSns1PtyHl
JGRGIxMEiFJJ7HBPmFFRrWxlaldA7hpRgEo/9Njz8mr7I61weL5YPRYO3j2shXQN
bfJMpodg6lSCcrCjuEeN0zN2mA0C1CrXjPdC0OcVuoesosE97qKWrLkEWU0/85Kn
bOcjfufOEsUpHElN5L9642yHAj0509IM3dN84JAFtN0PXw4rZybwuYJ9GsmyENIx
dWd7YhHWIEsijEUb25FIaf/dxGx+bAzHPFh1PxmG0ZmukxIEkhBsX4B7ZQC6mcxI
1vMBCxEn/GsDwqUPxEAAXucJpdVSr6ZYWWJe8Fow7gMWKKuFESRKP+ITlyf8G4id
YXNorNdc7zsDXgbclDyk0DAs3SpGyCtQQtxo0B+TgKmB6kEDDmaDciym/G/PeJLj
YVAZMjlQGV1utM81mi/Df4YakqUFg77Rxz/otrWFIootgMoZSRYV7AnL20i/d38d
WoB5GCOMLsMghkgH9Royx41s97DgHBq1We8olKMgLbvXgCPD+24Iz0NI6bdy0DbH
Xn9dov1QtoaylFFFL8+oaf4bBwBR4w+8AujVAlOZ0PFjYqoDE1uTH+ps/r0dhSxa
aMEJsj35ItkGX0xhS9eHY/EB5DJmLJS4A53XMG09LyAOErRjz3TqP2Z6rrwQWzYk
RXYh6/dOAQ5uUSzTByotRuO1llQfI49pHWideb4zWPf6CnhcLy7Jk2UcrEo4T3xj
gaqaRvt6CSWGYJIWS01zZTkBWIz0tROaoR2w1rROF7/Lv11ZvvuKxnTy16vRo3vK
jmmJPs+zdDR30VxoYzkbRdA9OssbRNt+RRDFzOVTjaCS2MGJRqjnNAjbBO2+9mxf
EcqGSDTrEasYsTcDzdtlENHBhGJv9TLZp6P/Na9zDMg8b/BPX7CH8QXL3ynsRAqs
UJcWwGyfMjj7cSTzEXx+dlD6QoojVVqkQWyuz5lNnuMEypktQTrvje9YXRay4r9y
au0VW0FzmdBWmkOHNG9eySKTqMtocXAl2fmXK+DENw99NVo/kg5s+HMtVdTTKBj5
DxxfIN7mLdQBE0ogSzDpDYQ/LHeJmIsJ5DzoA5JR90kobDJStOCN2J0DtebvRygM
gnUT3JnOCH5x+CW9T9DjmV6JlNMQdQHz1bRubO10reav/bkq/gg2X8EYCyp0pL2k
5YtZYp8bYXDjpHvV2N5/7RGoojbfSzNtGoT8XzGQ/nx/takO8LJP6IGY32pQQibd
9kKxZY1suxIuiRC7Gj8xpuIbbWje2E0+g89ijA35z7GUl7uNyy5Z7f+k+N7/J3mt
vqKDX+8r91Qlo4OsoKhar0g926OZ1FVi+EdYxJlDWvz4BKQ188qcwt2/Kf2hJgmn
YMmdGKvnmoEAe63bn4d87FNsSB60KZYLWTjJbPmety0lfQskUus5h4HErtwYulus
nvXQT9tDqr2EGP322FWkAsfclNxIWvaMU3+Tz2VZVUE7zKZz2db86hVjhtCLuOoo
MLt811C6nxjaRyUvYxcOhXjTAbZu2UDTjupNRc27OWvXi9fqJBMJSDhlqMAieHU1
KA549QRyEf+s4oxzNLMiGNn9fotGzl35fqclWp1DNKz/LqIWig/3ImVaYZCZ/UQT
EGWuhUv+VWLTo00OwftRCQ5TRZo6so2cQOkAx2SMJ8PqowLeptdy/BXFTUwZGjWQ
/KORWk2RqIIDhpXQyo2QaFs4DlYOTXIj379fB69GoCpwaY/dM3dA7YfA3TNYdF0T
F/ocShA0DhII/nIPJBHymRYW2DvlNvhifrRRZ+rEO+KDN4eQhHYAoSzfByER/rGc
uBJeaARvePYBE1KSz3iY6eUEZhMxVumy+QX/khkFSQgyIETmJrNnpajKFxdJjeF1
IHll6jnZ64uewHfD3to/bJJ/BI5H5wt2U+RVOw6wOFuUO7338vGeLrlDlDKRilmU
27xuemOb1ttmkjvJ/4X23mSjWpLn50kD4ep78t762WDUzNBAtrlKzat03DPduchh
zfA43/rxn69tnjQKMEluqVZt2Oo4ze4VjFf2D2YvkOoKby0QIEdHcNRKL0fOIsUo
jNkLtMqMwNnjTowLBBWmztFguMYQt1DM+wko0rztKSipJFOqmFrueOCds+y8u9q5
GygnQE0CsQj+h1ru8dyPcH1sY2N6jnXlwIJQ++viWrmFJp3Kv7KGY96s78J6TdTd
BXOSgQfUN05xXlHpWL5XiDNDMPVGxNwaz3VtnM6kiPghzMUOeEEkdPOeTY5FhKp3
JTU5qc+U+dAfo+uCDePMJgB7T7sso3FzCCuFntRinitjHe+BNmMqAjDZFT69N+ui
Ya17MM0IpcDBtS3sIhqAe3JGw5Ym1D/TS14bcOsVTD2l7nDpi0fo+2tYsAT55Kd9
heoMHKB+xXKwPDCjxzZe0osJUWDyx9105BkRGx+e0UbGqUcp/O1e+ilSsriNGrge
nGUV4+XvrDev1ebpuBtz3iRvfvkKrmOB6yJP5kSII3msYrqVTk0nLnXABqbko8zD
FKAHEYLF7bbsLyxyKikzFZ+hYvRJUE1k6RxYupzHfG66xW3kYoSNU6HkOzlMULZj
ASUaXTCGCbBLzzGOEbX8DzX1VHDvEm2B22qE8hSKnzkd89PsIJI0JgONAjCpoNM2
Ca58FPg0EFxFtHzCYDLTTk3y9Ja03nW8iYMNvmAdhkcp5dGEtCfbZQTLrHOydbol
Zjoe+sXoW7P8ODxQRWfg2ZN6CQ7DeeoscFTW5ZRjyB1PVgQRzbpD7Vs9kA12uJg9
oEH0+VEq5e9yjl+NLPa762QcutefjwX6CIAXjTmo3eoYwYQ/AzOB/JqDPaKHlb4B
5MueP3ogS8sIhk1SLWSvJEnSR0dj1s1hUUQWXPgpCCku60duQdqCZwZr9Z8Z1IR4
/bxLVS0gFXgnRxeadflXl8dW6IpLIb0UNp93F8E/C+GmXZyxDpXV+nsMBWPCrFGH
mPAIL1l/uIuuIecXYG/KM2NGIuJS95D6W4sI8fl+3ecrVq3CPY8ucKTYFuWCIyTU
8TTImG1FfoLlkO1sS9c42e9OJPxLHoTNGEdDmdfgrlgIlYQ23eDen2CNz3kPtUMn
qnL5omtzogKb6cms7mysTB33AyDwZsH9LaZVk1ZIDJHPMO2oQ7T/PUGonvTW/VRJ
DrW4vlIadxJsuBMjP+7ITWZyH1EaKx0PoScvK29Q3cHIz2h3LCig5VUzXQ+/kcvO
MC41b5ZaTUxh5hdyXFlivViXhFSA6z+RN7Rgyv68fHy525+ZB8ghZJcP/8cZZZBn
85WG4VtBIrNaK/clCZoLF8P0hzlusmudtpybhl81NaWyF0RPAKJshLfVZxlWIdcC
nzu93ZYe+puvN6lsZp+12LH6K6LY0o6pPzFh1l/FBj+HnAv5YVDCJyEKYRvs6MZY
T646WeC8rR1Srwd+cJaA48PYrwigL9xRaMWxL46g1u9sY1RmheAzbffB0wPh8c1p
ltdaJrTMqj0DRnishTTKIPP3ScgE7B2sDvBLAzzPLDxwYQvXXfhyAmhqO2pJwFjq
aBQEdbCjfVLi/8qVk3RRU4w+4C/gBY07tF9G+Q0MXJol7d1yAbhpYJpCnHyB21aC
DM4pw46YiLTKXSf/luoCEYGHy1zkcQubGCFQk9FR7j4XhFgIaGYdqp3FgHh+91Iz
hybOnXYM9s6H8L+09gRvlnf2bM740DmkhTaqX0m8uxO5FD6pDhTeNq5iW2RduYhV
rwJEXWO8mq53PRAPndGZ/OLY++iQw3bBJmb8vGIViolYSFsCG0ALXijk6wiNVFe8
wRkEEMzMXJBFxbpfc1h3oIj0kRcDxMUcWzF99vNTKuDQGTPLmqW3VYWByN8BWbUp
eKVHB3ZGC0MvPX43hvJfgeMEdiRLD3WCTwRSIWyRH1Y4WIKqcaKgeaK6vFmT3vhL
/Z0owW1kEVjcGLkdnUlVAGltvgIV0LLF2C4Dp7Os4A27OimUse0dBLD/o5czmIuZ
ykqg8Wy3rDOjlvIYqZ0hPBuWlXS16p/XwOeaj8qbuOT1uvfMwJOA99745DGxjeeA
yiRyi9mu5KyP2g1wK4o1djkA0SaNiCQPVQgfn8e5A414aDayM3BwGFW/50hRTd3C
2kSWviyzK+ShXHMLZnLFVKkpgoW0z8fhlKCJvKD+Iya8DMCGat4fo1fkqNNaRAMJ
cczz0WYqXIP62QYObFeh6f5874K9A5SMch7GJuIq8NJ10qqD3/XBBmW81/wnlhDZ
wVS3J4/T5TcX4YQNiH4w6y27AhT2jBltJsaOFsJUhP4aZJWNZyK8q/4f4460esr0
eRWfoQqKLGyhYX/xWdokHRI4ZbRTUO2llzB8AXLfqa3QZNFcgiOAqTPntdZWyXiq
YwLgkpMeF8tvW/i00q6er7Z3iFkkQTf8ATOf7IP9HdqBCXjX6Dn+swXP9PPuky2c
N+v44QFZKFRJbtCoq8qur/fjbClo6iCpUFoeKTG7W2Fk4IutOFDrIIzJ8WhXg929
DDIIfRsqaWdfougz/LqP1Ftz+MrMN6vTOeR8sHCvdFA5l3qvXS/SZY2R568X7J9i
Ouz4ft3XBJ+4XLWloxCMVOs60PTbtEhrjp0ToQxLBmon8MNwF6/Qvk4uZN7Wdixp
3o7qzLhp9j08CdjNONeUKRTWJBDwv55KmUaXeUca4suvz83PYYKCMa2oFqjKPpcA
nL33POC9BG51xenN0+FFyJ7S/x/t2NiuefrfyzloUsEb4aixyiBUGAAAtY0cXIYA
r3xCLoOGioARhzXk/OEPKLIyxXmdjEJWH1UyqoUVdMTFufPvmjRkcwwERzeN7MQH
b2+8JsPQ3dYyCs0TjJ7N4tXIBAXo/EBwPqB9qGH/G/1kFi77N11qpscFMl9AbEYr
gwiw2K/XW2D5Mr3As9uS+RfSMegO+jUNTlB8FG7/tP1gf9LWOa8RyxInDBd4s8wg
a/ma3QmMHgn6dII2jxlCp1p+0T05cPYNkE98q/8Ilb8dM7a2rVEn+Vfa4RXTSr76
eXMg6KCuGyrIMfEsw05AAeboOR7hOYyWs/KYRV2rCWPitzYg1IePfIWU+t84xuXR
oLugtEB061ahtS9iny9phIGUtzj0ZsxOX2iXc4/gqNSrlaDKB0SupkSsrSSR7tKA
Bjh9cyznviqCo7BAz/qiichZ8T+Z+vMUgUJFofDqVX98tVk491fOsnSlPbzTxtZQ
LxQ8bDZ9xGD8dYbmarjlQIpFCFa0XUmLO5A85kdxEr0p7yK28b0piw1eOYGOQbUP
UlTTRTYgvHUPz/SopMsE/O4HibRexpvRw0C0rIjFG0JCud6PNYHy6xNAjL0aF/LE
edEudwVUKb07uYhVCqo2uR5JXxZFZF7gZ2yKu/81M9XM5nPUrgsIBqMJQadaLZvV
KOmAgzxcuM+Zsc9SEH5F1auXGKQ1XJNn2LeL5rydq/njBTDx6s3eUXpKi2fCXWv5
wd0Q+oT6tNslreOzUJ5Lad+0M9pNjTqse3CRsWfThyfjs8vkdZxHk4kuAAswpIWB
QqF0UhYu9Q2g++cftLrFSNPWqN1Ly7tmqc/7Zu9fkG0Zg095mnvsw2dQ/KH0LkSQ
gsxbNnwFhnNnlKu2uHfaB8SFDzLzB1NZKGbPQvCz7w2VuTrLazQVyAbu+2CEQaOs
w0Sum/9YwSabbevvUXtAMQ0vm9HtrYPAMnxRTvYvtrsqRXUNLKT0Smz0Z6u9AHwz
puYBobxQagw3ZEVuSt9SXR9eMy4y4ea20n7ry2D6cHkwZucAJmhdj+D55vJ6+qIQ
sPxwSDJFAYyM7wzShCIk+e2wDye1Ta/5zHvCey84AzHUp1aMpgXIOTEqTHEb5Wfs
OngJ7O80CxSBwU/JF5DhfvLD9Id6Z8i83l5irXlDQka0fAc9pJQ2rCt2g1jusYTE
Wf4IwwWJnpAYsByfWTXr/47hIHpEkTphmI/2bPcl+LCVhlPZjuID7yqS4ja6F9bL
bb5qThq8zCyrr+RAW3RFuj8j/Y/028/Jm8bDYItLxMIjrR3HwjogX9kEd/Lpg50r
Xe9+B3QqLgjqUiOpn5EdO3N7ZwmwzYAVW5RV/e+Jy5AjInFIspW6lHS7NM8zVfoA
eL18wxUrdkKEy50yeThfaJf/2IsmvAE/eImArSOnDrVp58G8STludpRyjgBoiykY
SRQGuUg9jfCc3dqfI+rFaDyAZqRoy5RJ6pWa3ENIW/xlYNKZztBgct9ygMb49T2e
kQseqmn5NIpzVj0mlFpl2/s+MibpODCAtC1ynpC2sWkWqSpkn6DtAuxbXFE7lWX0
6a43gvqd6ssQksNC0pMQEbdi3Cka1GcauE9ORuFfwqKmOW3H3cSlqqFRGDomGiEy
RoBbtfrxb/loQQFLUuN56XDNC5iYPLlO5guJSUtx69lCY8Wm5tLgiEHhQ0FDWMbm
d5cKKXtjloiwUn+WaBEaNLKY0EMDf809PXGMfj/77HZXDxiCNFqC0TBPISt/oKR0
3BDGT9TsDP0e9QdtTEw0eDL9aSTlw3tzL6ZEp2rPa87nIQ3MlA6fjT7Op5r8tATJ
4Y6jX2SGdqVYqGapisF70PnRfeZmAFoXWlZzHotEgHdpTL+oomi0uGwiobn90UL2
yKQp6/LOgj9y/ich/csww9lJroINEf8VXXKMa2eyx1gV/l2pjrTzAe6T0TEiv/jD
9UUjOM78vN49HKO0VADV8O64iwHpIK6ImwjrArpwQYLxAM8DiWGswse5qY2k4F7L
gvDWh76n2hovNdD+V3pjf8yHToTKEeNzyZZVPITIXcj6Z5wwL+AQTaA8rGVieyQB
L88L6oAdpT5L1dTWaTYUcX1GTZSBPJExp3dmePLfVtWkYp23FTFAAA7X4S4hajC7
tmwLw7NkFEVrXzvXMuTWgGVOs2lInB8P+Lv28sCQRBCmIQ+stiSHFK7MWNSxOEy+
Y3bFiNk4q5Ob96COzoj82ibk1X5V8U1cDXMyhrekVrEDWCjTMI+ELZrSQy8vDCyh
F98zBkQf0LX590z/3KiYSrak8yVpwTE6bfzne6BBD/rCwiJBA0fb0xamonWPxvjR
d/56kIZlsSroKX/plWBYIW5q6R9VGSC+kB0bsuABf9/Y5masGyUwBCf0WnexX0jd
ZlCMF8ZZXmuNldrU5GEnJUqbRcw3zTbSN5pNeaeSQFqjc+SeU407xM6qLCmjOepS
7D0yI1jipcJKLGD35qXuNA5sbImXV19S+q1+N7gzBBAl+GI+5Bczl5V6oV3DV9j1
V0vuVDTeWQMfOAJ46yAfkmyuf+9kxbuWwfA0Qnz3v7P3M9TdaLGgz4lxuvLoqTS2
ZRcQxVNJh3nlBWW97uhRvYycDtSOlLZYuOcQDNyiipZlKvm+r+gHwSgnKEvGZSV7
/RSZdGjk7j/Fvbc0WF5x2a5JaN0n4N5VtKjzi08UJV234WgZIGUx6svD737CPkZb
Kog6Om/0dBAw0VbXkJYBLbZjM+DQSUNCHG5xNHGSvvNr8SXx1d/k6/f/DAReeR25
rmrg2akjyfKjNe6uzV0Cb/cLiqrZKFaq7yUIwjwp5HV3HMV8P9eX5MMRc4JS+UqH
gASssQrT8ZI0jtW8CbzpQRDfG8waxoWt5mTVZ7ygAD6ZrkN8iWQniBt7KBqobs2X
dhjnmRLCiW7qLXi4BebrHf5O+hb9/iHcpc5KWMLUKnfyAwnpJiLiCJ2LKhBipUUU
N33PpVHYqJOKGy6GgN0Ib3uOgDVcoCB8l94ksU0oRtfD2wLjGKDc8YykbW74SLhh
LhlKK9lQzLZnbENkAVYvXT7kWZ8REf7jcef1svGsETIn3pAtHJBqhlQWtSqqoJn7
Eyo7QcHAjctRhQe2KDJBWIwfN1Mnd5ea/p/z8lZpCbGDJsKX2xobWJzPCIlsw6Lw
zG00SOwxwUITaBC3eup9natj3m4TVtQ1JsrOKQOHh/dNI5Cr8rrIBZLjQStaze18
SKt60zNGwD4HDm62zxWiHjj8Ta7uYSOwOYB7H0tQxf1mZKXxOGNa1LHlhrS1s0GC
I9zprhB+c4ZKcMjBzUof6DT8u4wf2hszAKDybZJv9I1znwlYxnCJBXo2lFdC5+Wq
5jALHgVKJ6YUp1WblkuElkI8cTq2iAog9HmOzVOLGy0mQ82NDCJN0umgh35B7w/L
cFIXrR3A81oBHLWqGIjMpP0xD6FY30odcYR/3H1MGDPBuyxSXNz+D7anq8dlBxRV
eFkxvmAtcWE0ABZN48I2X3H2amYcUcc6JUFwZ6iJC67C0caCWw3+qCbAtzqrDuSF
jYz1vWeplinrzb+BFXI8lfz2tYstgdTcO2uQ5OlqZdoCXNJ5feC2b42B77rrJemA
iqOGO4VzFr8kLUSBmPnyvqSNSqc3xBoVLRhZp0AWjFzYSguB/vAmnkfnaLoI22y5
dWlqUvLdREd4VthBlaxQSCyYnrn9tyXp9fNTJuUz8m/V/uC/3QjpkwHwdOq4P0RP
HEaHSXzalnJI7x4b3Y4z/sJG+ME53D5WTtBBIoNwD0VugN0MLd69ir/1rtLGYGuC
Wg9ZFf6J3dJdZRK46OPn4Yp1sYmtjxIIEb9QhQvJeTHqzHg6rN3jw6ZFpqq9+Mf1
1oHPNXVGziHUnk0Jhpumk1YWeKtx6fO4N3X6adUaWRGY7MNxdsztt3tmOzKJhWc9
ds5gAe76Kz72glY4mKPuaqCMPliVDSUAuHokM8bmEz1EB3PjWVBqY6iBT1OpBCae
mHlP72lbUGCOQAgh8J8GQ1k2FzjlEm8cG4q+AohPMturMdvUzeJ8yKjzDRRbnVwB
nTpNsnqDdX0EcMuFDT2oL4w1Zozd9/deSaPlKHlvamGPRSui5EiY4r+n2pAkZERi
UuA/eI3QJlrMwUklHbb6A0ghfbYlb+qUC/hf84rLq4dJ9fOPaZsAdOS6+FrnUOfa
QYJlH5+y/pYmXT0TJv45ZswuxI+/+wP+rOEdsnwr/4VlyiPMp2FkPL8cTbWRJIpQ
uAGGk9uhKJonGbnH/AJOQYksVDn5nz/2WKqCBk5FqQp7Emz4L6hiBXuXbTNyWsop
HBfHAX83ICE4AnZXs1Bm1K2uTAGo/G8kiKrwMhcVs+2l1jCDdJVRzsVPWhUADNiG
cwZXfnWcFHonxdT7KjfwwIX8Y41yFBz6wjecqoBuEbyqbRIVWVCsfs9yY7Mtpt2K
0Jje+DRitZw+fXQpTVf8lhgRIHIjf7bh0Mh3+haUF96K2X+TU8q+CZLc3cG9c9FL
iBhgY8tnNRIerye2MlGQ+64PBsDofHdEcZ7iNJVS9klZXTEqdU1N16JgbH81q8nG
dtn+Vt3p9y2MTBrqJPulC9eAjwHPbo+ImKSohnhInU3U70Pj5BuuTdn6saR51EHA
TatQ+KLHmI71h0XVcfKnYKqB+Y1RNVIf2AX/Q0ih2gjqmauNXiqfpsPYwYtjfFfa
S5CM5X7Z91L5qLmDup4SAB68feHDARu4Xjp6/QyxhfTaENuCtBrMElpxPh5yuoEf
N1wsasvPRXflz9KE2KZxAiRWYh9kFvoUsXRCFSnTbFIv7AGiaHymkpQP2yRjUESM
L0rmhXsVwoNdPBxrHXeBu9FvlsKTGTvkKQnog1xtNZFbPxtMGtA27+bKwzfKbjth
AcDBGOtRGeNThCsJyCAsLw7D5KJ+TbB56EpJGsv4AgLq9Wb3ApZXODqHy7XlaqiL
uUin/vl4piBDxmsEVT2DrHIfelpuQwKrLw4v+VANexySNOttQwMYH7PeAOmepjer
yXecd3We4YlRLZoEdlq+AizjYeU9MQgX6G2Is8eK6GQCYU4ZYI1WEFdRzo9qNwnt
Fx5vFZRTH8clJMhD8RrJXLaa68E3rXIe3ug/WM9hg+zB84pClJa2D1Qfc/apPd92
zVh1KtVwyhev1S/RDDJ83eanKqZ0bdjaUmsiMnaG2T72u8e5oJh0cs3qwsKsMgme
m4fqW+98GHn75d7/CGU3SUcObBMcPAdRMi0pUT9i9tKaZSS8E86NdG3EWiBm0zQ0
p3pIXTpPH226l3OKvAsdSVTMDMz/fgjcRCIu04nn4QqBSwsQDmPQeU7cB50JUkXN
klz7PoZBGXoFjszXctLtvkJI2ys59qUT25IwG/EZ2QlW0glPPuK258qrvLZT1Yja
ZHcqIpwkYgBsJAahDfxs3Y3k5zgD3o+f/tQnZFy/lGw2ub9m/RxE9BPDCJ0a3P17
mMNCOhCih8V2uwmQJtRZpcqU7QLCjMTmNwuZ1uUjUw+lw/N+yehxXd9Wo5eUwO1m
mRtBe/eePmVQxpOthn+pgazg/3AORQOIbaEbDvTysTAfEXrG5An76JHettHOa4J5
HG3vHGGhJt3UEDNniDi0eQTctbUqxI3loSJw2HIcHzXOUH1YGdPkPbVSFlwJKZuT
itwBRByZz4iOcBGgDbBWtOapO27lVOpU/cEjk5F+ae+p5mhEFoJuDX5HolqjbRMc
dBSUk2+F5Q5s3rDEXnLL2uAcJHtQDcG/6nY4rR0Bc+nQoqKrfuhMT2aIqlizFTPs
5wAnJNec7mvmvCx/zg84meZ+VCQ1odYH8OxIszMSgzP5qklHvWf9AAp6a1Rvvkgr
JhmfDtrUtBlcietpPUfCWiEvheT/qSLpzpbf/J2Gyiwb1yYC5fX3BJuhWmyODfFq
BVjnzPBmPJVb/jsegK0nyIVndxICm5L1RcwldI/fe6K0lfqtG14bYcYJ8aAnjkNP
WFqUs/FDeJc2AcVmmDibxy8UAHJTX9eK6nW9UJItw4xati+CSHQMmgCj5fHbQZDs
FL4wLj3gpuWRtvcidS25umwhYVQZbuPJznpr5orfi5mbcjihcXy97EUeflHwZOhj
D4/qqPUdmL8o7RcTMEtbNENQBw79p7c0Mrmt+X7y4fE7vTduK087uoPJW8Ruu76K
cSXG/wcakKG2ES4+AkNrCe21OlmhY4IG8Q5/Z+Z2IU3WoMPT2szjtw1K1y7fbTDI
UdYIbmljFNpz40N5PGQf918PwxhXVgcRG5QR+S29gT/0VL9xLdTnl5KHrMZxPCNr
R3lfwm45XMUAnXSEnELgUnHsZYBi4SdH+CyxXFE9eJ2Sj680fjS8gAJY+1alFuy3
qVi4sDXT9y41vfip8O4JnG0oSNHjg4L0UYKNmS7TPmUsIOws2NLMkGXeBk8i7aOD
vo8DleW6mOtFD5EgOHXrM5q0qqoey6syMz7A1r0fFReY+OixD7PwYGwgTpvYtHfY
wewGeVec1sTe1ihqCOZ/2Mbbg39vvJHbrI7AK6cP8HYVl9dzI09xsP7XKw49Dhly
+IAnm8RuMEd8oDNVKnuNn87IuJqj0x9gbahiIXg7d+T2XXgtK7C5JvNt6p93OoIo
+K+j9CA7+CHXYvp7IwGMDKtdg9+3vbDZ1TXABNF6to3VYv/zIcxUPC12arLbXIXZ
VqPApFwSCK2+IWo3bC0jDYgMXiga8MbbWa+pUKLpPKLfMXGFVqbQL2nNTvzD3iKo
EtwQeCdCRUXPWaGzW6NMNVQnKIksGHdGXq2cn48dSsLL09FUZqZL03MUpDReVYZN
Ktx+BtvPNbl4mcnso3xBgJEll9hi6FYKZEPoZyV68Oez8+2NhS8B46PnPQJk4RGg
R4rYAzGBJwAeDbZqevYIcHkFoltASYc79xXxGANNJOFuUoKAjyvYqarutQxrh9vq
jSCuD13ZxjUqTLHJTu3OUILwI60OQU7TllDfqr2xrrffw/OakAQNI2lCyFpkiDZ8
4b48dgMpKmcuHeNLALZ1w2W11uNwW3dp6eWHOyU+Alqie4UnrDiFqjXRiWvcDVhz
lYtQZheKmFqxTEsxHLCSn+HbGiIefIWjriy2uHCMQfQ92tqkbNNZd6atOx+Lavt2
6QBWvQzmyT78a7wMX/PMmmQuokYX7iWZPPuyKe5CV8Y642eknjOGf33/2bsFOmpV
091l2E84DrnkJyok0Bq0lWRxsMWPTKeHd4RPVGobXpRO/zQzDi17pKtDrlbQM4JE
Ko76wpJL4PvN4Z0rbFaTFZ62r1F+0Azlcn7VOGANFKRRwYrKTk6DKJWRgDsxBhTO
hdZ3Io9CLDpdoJITGuBuOUsIpI9nIvKXkJAAo0hfWZTcpMRsxRojD953XqNyYL5C
ojniauz5deYBJUe/itqTBKv6iJjhFFSCTyBjKb+6qzzBSBt75bRGnH9p0NWUd8pi
p2Qhd5gakupFd5LuzgFEs8JK3DBGc8ECIsqu/JzUp9D+EVreBwIjaT4Gkgs+OQhT
NMO8uYPL/SG/Ukt03aFRg6PDEX9q7THuNq3VG2RqBrWwNtKy96vU+WSDuVOv0NoF
roNuUuOg9OoTFkndl5WNMKBtmBUUtj2JpDXyBPXzUCOYYrChVO8kCTF/pRD4PKrW
Z91GnidkC5VbmtA0YF9C4TQk1dOkn7h3tPNPfKgqzgMc+hMP6xTtgJ/JLLyZHMNy
1BMXDgjKn3kfutFo5v+LKl1VKH1Bh3gfNtKD9Lrd28IgBiN/kPBq93KjRbjg9mG6
LF5V+gN8XvyrslLXoNFHFlz/33MoLwy1jhhqSOsYEWo26vQPtnbCCO60g+YK8/0W
K+9QBVivbe3KqDiO7lED6kAA4vROXpc2JXN+TWlFhPCikqHxc/3EnvdDR1Tfr4kx
RAXGVeL9YKSQFrrriilCQFAXfueoYxa5v3HTy/we1dcZtPvGlyXovKSXziN8ePfO
ekBbJ6aj8/QBWlPKBXyP37cqgjhiSCqJihoWjXFUaBC1iur/ycHZ4vuQCbIDdeCE
1d7Y0tzvazSNzkvurvPJ4RmsdXSdSntye2hI7JcvvrxUBmvOaMOzDwEGWVfJ0ePq
RTm8FARd5ilBRNVTN0aOX/nBXZW9VgR/pfvwPHiClKX55E/vu6d69wsg8kL6mfv5
5CqyaMN2gshKpn4c+9n9xn9rZyXnbCEdFYZDEvrztuiLTleUfbsY0ticsOJtEXnf
o3lThMs33wuU0pSv04q69nAQSQFHjsiHpgjULd67ntM47squEg6vbC7mP7ixRUXT
X7vZhrtKtJVArA38gDVy4D5QpqIIwlygqi+4EsRt1akLEjaGSWNsWBMZG/9YsLiN
/EycKSLTbsc6XvN0rhO9+T+si+By8/L+4okgoGl1mO6DXWqMJ/mbtUV5eI14aHYn
IIb2Z8UI5OlEodMMpFWd0Qny/t2/S4Z/m7TmZPHwzOVB3bhf/5sYnB95l8KxZ3DP
8efaTDIvgiAvioEx7zHE4NvLNYXuVwZb5HJMKnbtgUN1Ne156+u3zq23LduQZ2CX
ov+evshs9SwWjybe1UnZrNMmP/JWu3qELlnr9DdpT7Tux4wG64btqTL506W0xMEA
OgcuhQ58NjwEDoVC5nv9xalhFhjOX5qcYogt/iXHF6oL8EdQcyLc9xZvrBjxiOFY
UFKpfpf4aHHlyWlP109t9W7VN9aaV0AQcGmqGLxcyll67/tH3TeQN4CptP9O5je1
4QpCPjrK5wQ7wdDRNm/1Jak/0scFL9ytTvG6/QKNMeTG70wI4zH8ANV2/nAUTDum
dThw8/vpY4heuxGsaCXJB/JmwAJf30fR4wdmy4iEGZ1Egr1Zb90Pt/sz97dpIKhK
/sEPIzJT/GieuOwHQAdcjMHOIkl25DukSaFcY3JsTRBO6JBvYsCBu7e7HNsurjiP
go5L/U1acUAg4TK3hvuz2BdqHCGWCjZf9hnL9BVLuZNGq543Z9NW6PALNqqd6f3l
eqfg8EFqiqdskvtoneLJ423yb7EePvkOaE5ZulJE1qEmoWRLiFCEbLlkUN2k/dqi
Kn7CJGNEzZ69gwOrff9TP1TlI3hiUSRUNry/gVECW97t2PfscNuyEyzaMCuwn+7S
Jsp0Ihb29XxYE9VR09h+9MP+J/1Lp3cu5QO05ePFkpngNJXPsV75A28MoMCaP6Y8
bls9gGa9hY+Y73SKIlEHP0S4CKY8TSqayKUKPoJPerVWqgFWUtKOre6YzIMOFOqq
sYG2rZHyzSWHSBTbcVtkLhsucefJjLDX5bFZmen4Dxub1VttRmsWgu626zShivvz
6GxDlHucvYL3DhJj21X/p6QhayvHgq+haG1q7AgovxwjvPfABliy8SlNH00X/GA1
vPcbs+pLZdS5+Wlkc0CLXUHWcdHiPUWx6D9REdGUHbfDSkqlqr9LPH1O6aPV7ZMJ
qfKvqg3fInUX4N0Fo565xh3HS+XmoMN95ZtsYd3dua9C+8/8mLWfejHLftM3XrBw
OKI0mJdDlSotpW3vnP+glp+SaElszKuk/p8y2cIBiTgb5eKPKcqWeUDZPQFVvX36
cqk4NlTgneNb2001g3YvS/7cBSpZeuO5ug8yO/GFqoPz+1DhnqZN2y8cBR0u36pm
NSi4f9Hk1OF7vXMz2iyk2W1Zx5Ia1CFAYLki1HiKGsegKQYx+NUl+GERYWFYEYBX
LRBLxgRW+hfflPcJScgb93816opSbjndqvpe7xNcd8RMBcqfc2xo/JJgE8rwX6px
32TSBg4jBnvSt7wXc4z0PB5WtRd167Ft7PBnxfLLE0xvbHG3zGiogx4Nm+ctqe3d
pm3q+tWhfgyNGD9NzreqjSoXNBP5VV4CRXyVHHVVF8gha9nPE8yqyJ0Jix/0i4Fx
wCNQ8JXRFnJ4/pr/rJRA29CjWNb9pRtCIg5eZIpgLPdfraSfE+Gjhw5NhKT3neAq
nWNQDoear4LXJ1nhetBYGX/hSoM6jeGPLqmClxV+YABA6YODL/nyep+L1K9UJEDT
B6TARjxl9d/Oo98pQk5cilVCgtuI4TexUNvKApBMKgKdLw3eZHh0hG/XifOXBfco
LfjSonhjyL9j9R/ttMLrd6Sz8plIg2gPaPB2rn85cs7ptiyAfRQ6BiMp/AdWdQlB
DFuypk58PVcsAzwkVjfF8Mk8FmYdGQwQ0EMD64dkqgUUKdOI+cSWlk+mWZN0FUxC
QhWmgEz+1Hp4GNK2OV+jFVH9yxM60a1kW+A9diOxLlfDPw7eo0ytptcecc8gK951
ePRAR04dsFOxzF7waiTRK6mE5GgTOaH94h7OQGR7KyhBFZIVV3MH728NfkmFwKRL
vYD7SWdpgQZIOn3X4JVAOj1Z9Nw/7LoyBDyZyzw7z6vSZXBRVR9jImuzlGeuChYO
FuxG22pgOGWgkGO1t94+x8AXKqoGVFjIEF3wiDz1FgER9d0JRqdJAeDZRDZjSxqS
O28IJzOIVu+S6VJDRH5xSWy+rkqh9zbtL6QXPY7TatNmYFXAekiAFHem2fUg5iSi
mxYDrkZOKGDVBRuNi+7AaaTy3p/bHytzu6QCR99sOZcCVKIfF/Lp6U21Pluf408y
uIkZaj9F5L6PAg2FP3LsMD9d0j6CYX/XrtirpqzViG3R9uUQUDjKhZpMuUAGKgsf
jYN2TkXr+ertKjKn/QLcMggT9jNeT8gSmJNcn7mny0d2n8PieoIVktausRwFsibC
rcDjckZpISoZwHrl6uCK/Uea16EqbW05EdZJFfVe391ItRsUiJo6w5Df0IyKhpd5
x6MxIq8N1mRdOIWczu2hu9Wk6g4w1AEQOnodXqFIVvqDoq1FMK0RJS41/UxEuJRr
BV9aIRoDjUPbij8zkfIAGcWZBNTeqLBZCvNyL74FuX4ihqIgTdiwwqF3shllIPu6
+jDZFfnzQM+s7yEKM1P2aj5Ihii+2/EToN7jvCE5W76iUSv0Cc2mv68C5aSJtdEK
J+MwpK1VP5op505FWBP0IOeUg0GU063PCvuTpzX6D0Gcc3cshZM7BAA2wluPyrzw
v3xptxLhG/9e0SQhku3X82rV0tcWgem8+bUnrFQpAhEexkQp6z2z2tJQ+OAzramO
X+8bPi+ZnWDm9D62+CN3NIBxKn3gJT/r0L7AmCxGSkwgSf91rJD85f9HC6SmiR7j
mFLo2ptqjVz8Uq0xkPpH9rjg/002NBHJKq+PnMPpHMnIPuRYUL5oTfyoZhv61vT0
iqQw6IW5ZhnQjNlrGQrnSm0bUHrVwZAP3+eQn8OINXZ+ReHqbwF1dCO4ME21d6F+
6dMdjItSCtwuc04HDO/ZUsyKoe7y6uKZO3gcFOWfIdJ1mwV5E+5iURxZo13FUT5i
7rnrdM0z78eH8jY+KKNpm+kQeWfGjUWN3QyTD0JMgckdwK3hlxj2q2+HRiB7q4p/
uEx5DbEvbhm6fvJeKSLMgv9jDbUTseZ8wFQirbL5C+FmLlH0+TyTD4AFicxY5fzU
bRuM8aBz5wgtpTzQZtpK+5AP54/dB+iH9oHFn22meeiS5vTAGOEFDpVvXmbfI9mn
b8u/Scp6uEOCAFSW6O+kSr4lFOHESB/1v6A/TcBS9rcx3di+1hXkrg+AuPataGQE
XqnKnhwEcjTLQ9CbdWeizc2Wng7raEp6LfJGyUFxk2eHfUSHAEqUAsRUoupcIuc1
5rbY1RGyz2SX6BHbR1cCAlox4doXYZuPbJTxo9aQmRT0wmuPFkN3F5RcJsOh/wAz
4C1LIX+mZS/sYawodzSZDQVx+l74pVDdRe2S91WxyHEuS/uurrz1xgF8B4jqKPfb
wc0fF2k6xuzwA23BPWnWmCEmrzECtaSRNcf3PlVcr5F8z/KKChuLLRdu23z8mNkP
FnKbDP4yrXdZhhLlhHKwTu4h79C1aANlDoptXbap1CqSs8xhlu58ySZJq9iMIalH
EKRksGQBtoZx40M4Khi2iA8L2OD4mjVq9ER8EIq5E7yCtfFKkUxYeo6BPcNT23v3
S+8W95X5Q9unzdh7ctxwMCREmJC4AC9qF1PU0JqJXOefdsHQeIppiGuTgpAtzMHG
zZEyx/NoS/22m1hWPLFTfMdkyre/cpjbUtZbghH3oE+pAUu9gknL1DB26BBfnIkc
6kvy3WoFNxQgiD39QrdV0zcbTZ3X7iH6gdIbh8qUSPYt/Y5NC3IzSCQfIq3D6biL
rFmaxcTaeumIOiABVF9sw7glVB1Q9WbF4Y3m30F+5rmsHaZ5DRmyNPk7/GLSnR6I
pdIT8u/UvxQF0KmwwFNuEkMH3Aqjg74fN8Jy0BI3mzHYbgXe6ONu7XUPbQxRN6mu
3Ayqq2D13XDvvelyutNlX35bil+9kIabU2yZSRlesO0HNf+di1csVbaQoPlUgo+A
nIqxZQD9Jh73j6kq723p4GjAT48Go9BtK4yYbScfZGZ9kw3JtVTRPs064nAaZ3bJ
FIf8vpAR+rbyZqnI3TC1Ox5QgFl7afF317mvXhUYBjNgyxvMcHEzMBRzq+DaueJg
1C1F1SUKCayqn9wOP81q+NwHcdeNKolzskjPjt97646T8oNoQ2xqB/Y9Xx5aZFkv
XKKzxUSyuB10p3zkKkpQJrz9tNWpMCzUBSoX7LqHMeqAKo08upvjrdvZDb3Bqsl3
xL16JRHGK7PYh1NzwjbnQcIb35oOuh8iuMrLC+AgMnmju83MOVEEF5J44LjaBBIf
zz7iezticTDR7SjWcaoNiU3xk6Le9kQveFvpyHm5cgMrjKbgzauPODn02Z51yHE7
43O8GZouBfMRBSkWnFhI/fgSVinEj2xprmkI5NUXMofALO0DuhY2oGKAw18J5Kmo
punsmihTavwcrVI18jFHsLOExA/dDHsYF4H9uPCfyIACKBwXfBPUDrKFGEU3nZun
N1HKgpwjgpm0ee19RKRPC+z5Sl1ygmCzYF6PmsG01hEpb2KIUDA6by7hyYHh0otS
biWnEpVMuys6yyGJSDmqKQ1n9RmWzEgrtUKL83lJ/3AGADe4blpCmCzpq9V+MKYY
O0OSy0/qGS505KxCDSgeA8DmbOkYqVHaE2be/eEN96XckCz7d04IWSnxJl/TesPU
YH3knsEJi2F0eqzjzIV6D4mL6AxGJR9oqA/tJ6eMy1XnEVNJeG9Ep2Gumty4rGnE
TigCHNdxEKgCF+/nBWvfhEkYM9XUlwdnd577KgMgGSXRThwBKbyea/nt4HqvHKz0
HHhJBlQNRIGP4km3vfEQzZWzGPIrAcgsGv2vHfjy2Sqt5hOAbYeYR+ybQuRoR2Zb
oO8thyZwtrgtSkmM8q273HxBOuU77qgm+ontH4pbyX61ckJjVBw1MTg27raRRiVY
VxdLzhcJfny4AGTQw8vTQvGQJ97QfnUgKtzmPofV4lagRWGezn6wkYCFi8UefsYX
yi9DZ8b+toMCSiMUDID8ZoPYRADsUibAnEFGvaUEqVlfFNkXTydzghulc7EwXfAe
EJfi8JdKKVaLdPT4utrY1pO9EAMocHD93VEK4zy2KiVx5hEGrOXc5oUcxOfKOuDD
UJYmW0EWnE0/u7CVnD3VEP01OUO/nnWfeJ8T9cbSot4nRbmaqH8fd9wbAKXKcCWi
axXnFmoQPLArvovkrq60XVQ9DdKbHyePGxNTM93hv4JCX9rNvtooK67wJMkIcXSI
bnxrN4n9v4Fgj/qCgnxgLlHp28LbvDdiziM4Az4OvhvjJHg0hrh9eeSmdtBfHRzG
isA9r7DiKLTWnn/suCUmxH6Jm74psMeT7Mfaitb3MyUFv2gTFbaDNAy4tYcI/NQn
GhGGx2lSKDzTo3K5blSZB17hzt+IQpIzd7Px6MGgAfWKYM3ABW4wr8lUGCCJTmE/
HgitLzuGBeF0tIYqhwtRgXo3+DT/JFAa0IjXGgqHmF2Sh+84fZsOPHMQFl60op7u
jG2KsvFslqWMgvcVdZCDsjJLt3DbD5BWNw4EbperoZw96k1r/K1ztdTNw4GgW3C+
9zZomjmdGGFC+y6YNJSHnnKgOEds+eFuj8GMqeesGSc+7NYyIIld+eBb4M4pu+1k
XLKmY/knTIBALzcBasX5ZJinK/8uhftCGCn/AdDTanQ/35yYSld/uClY25f8/Rez
ZW6nLWM/PWRexjggWS4drHAOCbqoeqPWGYZ4szVs7Lq63OmwOpl6EJiahUQjsskS
EcwCJpoc+A2rA+ilzhbFJ3GFucXdPZ+QLTnDTjSR01uza44A1H2fxKo3vTS0NGr2
eXble2LVyUJfiXIvRdu2jhSVLB0VMCieKXYeyctwXOupiopQC5ZtVvhYzXuAGOlO
/cDmOCYJRQxq9xzW3o4tXRkMc24+RgTz9og6xSZEWGP/VZepz8/Vt078h+9FSkx5
cqugDvW6rz1fGVHDCW2FoHKHTcOIT5NfuDD3Z1NpXUS0YGf4v3a1BDlLzmlbWTmK
sz+LEvYUud18YBIKQE4xa0GGt0f/+Nc/ffvfuXQN2/mPfr4TaSsOvthw+dinPk5W
qS5VvDJ0TzmkbCCWcVgRCdsYgL0c2xdJjpLrqirvdzI13waGGycooydCZbUS1VG6
IVZ0fs3HVphk2oeSi/xHUPJT8S/zuEtcovKoR7pvojStlXI3GnpmbJoekcU6AMFh
x2CYHR2bmGZGKuslFycDft1uBcM4aaVWK3fleqmM0009zp4mGGqavSNmfMYeHu6q
6Lkjn9OMwFmtT6jd/J6f3dYfmN8ewP0ek7J58iU7YrwQFv1+ePFnyyepH46TsEO/
i+o88OcEHQrQTCh1vf0qVk3gHDmPSKzACFMqspqUEvPzQesAGSwTSryvDhIP/oHP
gw+HdK51zox3ukcjz83nWPO85GGnf29lfnVVflIdH84xUchzMx3M5Q140MUJcEL8
mvq0FFmHYuGU5ujW5V+Q8cIhKBObq+I+yFCHrK3rKG82mVYBYQ1eonL6tWfQ7SsS
MGWGvJ9AOBcyAQIk9SRIAJEqkkJIKbEwQZk9uVdhIyT2XLPBWAxGxL1rGFDk+RD4
yGmy8A5q1OVKtZ9hjdWqCKU8LpEW4dRMa/+TfMytn19XYSViM1S7zIJLCG90K72V
2Lt7Lqi7soDY73hONW6EdmPSb40ueX3+GX5pZMnKvJ1PUqYKz9dsQ42bT1Tu+utq
HuvN2bJAhUuiPC1p8yuEf4Do9eewjsqL8s1JsaJkDRBIDV8xRzGj2NvNX44BIX+O
vV6lPn99fYkeM8Srm1DgeLp/pSwfq71EAc02idMxAedDRjtwL7piUn7QzL4C5gNf
L36ivD2TVvvitC6MY5qx1O2Rw8YtINiw2VR2pIb9G5a1hggcjn8JXatuYDZ6cXel
QBn7por82B+CFunTsAv7hwcg2LhF6s7P2DlAfPqo6RZP4pGfKzoWXBouEQrRO3XU
aiHMtWCO/xye7yU4Iedg+cZ4dQZpAeOVCYmWy+ByMR9eAWySDli97c6kPLr6eFZa
bEUcCHejlNM0y3nGiPMMXrl/MCdcylsIcO4IRM4lJNpYbzKZ45FTatiwEXcjjvg5
4ullFUuT2Hgxb6hR7de/zCb/lGJcO1sWcNSMAasIEHJogMv/tB3bq9v+UTGSoGVN
PpwcvU/cq8npo1E4o4NTxt6rtYQxClLD3ByG7oYOgP68LCGjUhXc/vrBn/52yPya
gYWQsE6K+LPL4yD3d886FeN7xoBJNN148ZBkHPHCckaHwQGX/HsiSinAKgTokfxW
QaLh6vWEwcC0V9KBdq3rQvbD/YXomPt6OBI2dWQFD5ZaUa2YWUPkoMDW30Nqd6t3
A8DpMYpS/lMht1mzmY/LVhYQLdbEU+LoIeG/To4cORNeNVSzBtONvQlNFgAGkvQD
7NWxT7YRCWiuoR13qOmiVUiU4iV/WMEc7bNsqjI803j8Op4/fHLbQ2TN7oAE5jH8
vLFkaastgv0v3bZE61Uf+37/9nfU1Bf+mgMtUbm+uDHSTk4wD0YnyhyyKp0MbJbM
wczITcTJS5lT3ODQ5HhLgq6Bdl5NMonoviXwUUPy2cBcF4j2XM9eU9YJAi12F46V
4Y6WKj60bHGC6a6Gzus7czky5IGPEnbfl2HLNmBM68E0ZdyrFG14jOINV5sYe6uV
iHiV1GPmLy27g5jHv+lYjZUUn8+kHh70bUdDHt+FqM9FIZ8oaH46FblZd0/spD2G
o/cEgneYmOrbDWjPoFmbmaOEawp0detdplPzNzmfj4uLlk5AX7fhzz7cdHlImmCo
8GuFFXx/c15725fUfSQZUotGcIBlD5MVmrysKKd4kWh8IhuGLVK/4fXK+de4gBHy
S8satFr9y8EhQXFYP2o3QSlBndf7TIXF4e5KK2NvWezcCWtwbAa1mQPF+Vi9LKo8
v2B1NvjevneaoaSksBMjHodyz+DsK2uVIohGq5K1SFxvXOXEPOCLMuc0svT0spcJ
z4/bfJkpFvVMg8ydEvsfC3QrDjQbshYV5QWCXsf8iSPMDL+h2g9j7OQbcdRays80
tcKl/E+nTAIXbJ3ctX6myVk72dblc+s9TMXkGwJ5dW4KUuctb7ETST6Of7sJTl7L
xNiPoJQE3EXox3CN3hcHt9ekJDFRsJ2TP3D4p84tJa/iuSBrAcfjDzEwOS5lXLcG
7nxiFI80NO7Jfv8TkJ32HgTp4dvWmwsTSLuOibgalZngnPfGlYGLRbvlxVjWdZZy
a/8uKj7Cl9swt+5noBylslyITScHPrPvQaRNg+wtEaqRlMfUPBehR5J7cYaAEJz/
x7WJkcffwf33YvH4Je1+MSlKB3dSp/17yjo4uCCbeYd4cV/AN2mbjN1xWaWd3gxa
+tUulnzxedOpFTfCW1Id3D0Lv2q+Fzn7vT5ap8X5PP26RkRNuKi+YyyOu7m4MAKA
xabNsiJrqrBTB8SNobRf22dtgvc7/ZNguxJYO9BKytqNgwREy4lIAQfOQ2zdR2KY
66QhqgoBbhuqY0s9IgGSbHNtQBtiiHma/o88Gkyg2HqJxL+qdeCBj2mJM9lgyEQI
EB3PdM61mUF+YQ/kqrRmEoSMQiaf1Sb+NMaoqUO2XWOc4LRfQ7MUD3rhmQlyogFV
YVZine40Wm4hNJqnPMR2AXhE73ejjbDRiZ8L8JOtdmca30SS+SkltU91bOQ1/g/y
vd/3BKqZptZAxmD6+pdDbeElXY2Kcztolp8wexcLNU0T18bIE3bUFvLVOxt5Ha6o
2aPM+mfSKWKeU6TfMtBgG2BRz9Q97RRzYVwK8FBaEpT3dMoiQvOeOYdWecMsEJCW
eQJiQcIUgSW2mjq2b7aC7a2yp1MP4RrgcXsF7SAzDX6n7UwnIsdfQTg4jVJ+nA+U
dRojq+npgvRrdLhWb8h3bfvCTnVtRSVl0BYQXsnVhGtr5s2q87BR0LoPiuSlx2HA
cppslz7Xn3okvYh8uqEoAqw8qigvw1MQWt4b2SJz8QbUo/wUXc7jzlpUWDLVn6+M
MBNAeoPjfa9lK0qpO6bIp4od9R6q2cXjPx2ys60UBRK5KFMF0AuACdu5Z6Q1Tn92
QQb7C7C+HBGIhtEngpmWcWq4L620KBNaeQVZA+lrdx4AiN41Bbn6CQh+bPSfiYYm
qwzunLG1MneYegCOkrFPs0MpSDK099jUFGjHsjoBHhU5n36szH+hAJI1h/6fFfHA
tpFwljpEErL5/ULsG/zzNiHWe5mas6nsgscisI0kgINue8PRm8K8R9aQCxIJUzLN
lCABoToR0/MbJ8S9Nj5srBYDGqbl3UkrzS284o5JJzLV1HECRnW9D7R+qo8lLeoc
woIjquo1MP2Hzmsy3M6c45wMauGEdQsjmqBKojxaP0cfGkEVi7vSVTbAe+Z0HJeO
e5hws5AjxK7cpzCXEK4SiSTezVeayrgIqkdxVG6EiKB73rbsjnNDSCBJs1QRYu52
X2h8S9TXNIx+5FQ6pO4RZ5kbdBtntfbNdVNjOhviVuXMIgsZwiUMHBjJVoju/W1F
p6nMzmlUMfhXl/JDGKGAQBfmIjTBlqNjRcbhXqMeKbqk9DdKCHsAWRg8gfS65oly
vEEBMpJbgL1Hg48oZgnWYyR8EysIhIoQ+qSSmO3eVKi9rOX4XLGLCE8PrNKVSTWC
+yN/WVuer5kMP7FDVNkYILWUP+9RkBJ2svvt2bK/wE+K3aabtegdV5xBG8LkEmkP
9bseLjGRxeMQ0/WxRD3C/KEWMkcWMa2EqwvIT6j+YKyl57/dqiLYSt1n3GbD1nEM
3O9CEwSa+8m+etp8ciQIJB4vBVrXQdUcs2XVOVrdvMy4ypdkue0SLf15xhJMCOPz
y4VbZSanXOWpUMzYiRrYUi3QpwHLpNuFX9/JN5cW8ctw5yZBJ1iTnmR+PSg3SFgz
9aH4hUARYHnn0JBz6bnt7S/gqEKPvgkwJ1s/yMMJNL69z+usCEsAAuURHUf8vUH5
VN1Z0jd2e0rJnDR40VswLr+7YkAyA29/un5uEVOqHKAP1RagYShboc7gFUbMCOny
nIlPHzs5h7AoKM4H/26AzXCzEdUW8q32uSY3gLmkw7Yf2ASjbF1hEVJh6aqmHzYh
rJhtYmHvbVViBW0dNOM93qCBAeA0fRr/CrDCDXrtKyRnC3RurX6QZTI0UhLo1a0q
t6NXIYMTgy3PUsCzlnlB4x+tsCmnG7RZeKVxhrFVc66+dadq2im9/xad8i/AmuHH
70rj/MK18dgxLJpb3XZ22GWwTc5jLjWKCCB9m00Azz3oft1dGUFcbH7jH8Ye49fs
BcxaII4XWcLqIRQG2JKGKMRCVPxXwFlB7tyW3H8GY4e3REwr0RIbqcbc82r7NkMr
lRSAvFOiXzeu5RyPiGbYNuPg87uBzL40KK+CWQ34W0ABwIDbxcLfsdsahIqS7pB2
m3DaYFUFDH2jcWOO91ZAjYfWWWuyU64PzGjeeHc3527a0Yk9Ltlv5hffDUKRVxyH
ld/QgvXewq063wsnUp2QNJcWBV365dJMZ+bpwFbW0qtxmzR5OcrapuXJ2UZl7tYd
DiRAM3gb1BbhxO9MMosJIBiGTr1P6BC2OoWAL64PnMWFOpRrkYgFHWXBLC3PV9si
uux0W4uBpXmpSrbgHhSkbCPHL9cQ89K8dhZ2C8CDJrxbLr2nA22vNETg8HMwjI9i
p8Xv0lD8fWJs1TK8u/Qh26JM5JdynVMmgMfWgPW+QSYGuLo1e/W4Z3rzwYCHNHeJ
7kJebhKfxa4Vs2p9opC4okDoPrdrkE51YuSvRSJDppTLFmzW84iHHy9zqAviFVKw
us49AWvarxYTRP+K+lTXWTl2R6jps+4fZONZf5RcbMBVf8O8xY9O+cSSw2gyYTL8
4O85P2omen8aFYrKc5Ccy57S1oUG8/FuhpA8HccJ10OTFXUp2fLQ+6CludQ1cuNf
FKYLUrF2bc+/TIIYidrz9U59LnO6jc97Poj8ny0oFkpF6YLCaHjO2qKb7XoDhJcK
08yfBj5799j/h1MgyiRAeyYg12kGe8fYC7JtY+GYgeHyrcwH7XM5ZzUE7lX9sVwQ
+cMmIbCy8w9kIOpFphxQly6ohj8rpmO6s0ndCBIohCSnzTMUb3lhas1jNE4iDYSW
LU0rYXWjAViLE/rd0eerhAKAOcYG/RmscibqlUVOYFS4ywoN7wcwldaSP6kI2XDv
hG0YshwCqTq8grYgx57YxMa3e8UQlv+QP7PP4BBE4oICtZ/R4tASTNMvmx4lHzUu
yL8EZtIF8ioO6PCeOmexGIpsPZYaPUsCP41xHt9HLb3y5Xs9wl9atgMuARA6Wfhe
t6bKlttO/utff4zJFy7uEvYD6iNk9zhzsDwwIzNDPXn1qou+5Uv5Lf5WYoN9kphl
vaBNPTuDm1aIshMxP6uyi+FRDJCdqT+YN9uTwcg6Vww9gVc1bTJZwxeVA4vaq3wH
9nCdtPjecRPDBT/Ls0sibMMxeioJvHSBeUetRSoazHDBORti/3SoGvkhkFjzmBJU
r/Y/IFbSv/HRD7eZpokhAgcGJBsUXqIx2vuxD4pF3TyIGbvonFZR3fpDK9b6y92n
UFbIwKihG98PSBuISI74BeYyObSm1kMJ9r8QRkQ9QzZzRdi8U8eNMFxKjq0I0A3d
JT/M/2wTx6t1SYZcwXthqyiU97eyvJg4BnCOO5e9EW927nMX/ited0L1H6u7PgCo
G/SmWMH2g6CWOxndyZduXGgkQw+fN3Ys6tAHxHB49j7Vofj+xa1ogLMtiKtT/9Ez
WbcDAVJLXNOWNNpYuJM5+2t7Bi28lyvrE4AHEo/uWRJOUwOY7JV70Emjo1QZmro2
ZpLIlTg7BwI9+ZQsCXM9axKTNz7YwoyRnRCYLKC5kXdqoxoZU4t6zomiTL6EtQwv
pwdZMkMBBZC+3iWaJCS/S/sk8RDSbqb+UxIz3Ox7eXCsyUdls0njiY70Qs1b8oov
iLLRmdF0PWQHRD6ndlEVPTwL2ao6KsxNgRH7+SjuwfipTtbH1YohNcZXicODRtgD
REx/9it+6l9P+A2WtK20qKs30dtwRDlsHDyzI0FHLSg6zCKLxK0g7yyLlExbzDag
kXFAgHngPWzmz/3Uesdo6khH0XG+nx6Mps+OHHGRj4XBCPih4TGr98VJZq8ZuKAe
O95Em4eaB20kn4iL47UgQMqS8tWHKZJhWPtQRRaSjLHZuqVzSrLSwvB/Vvi4rmHz
Y6nDujh5UiElgfsHEWnpmcp0zUDUB4SqzUk/duhDD6a6WLiYFT9kxBFA8oRFJJKC
I9NkKTnpCxoSl3En17CFh8Cn5IBTtuhxfL1TaRbn+LZjmBPnjx+zfAzvOT9/xdud
W/LmGGk8+jidOAdg+Bu05OvVvE70LhqjfAAgTD+YK7OmieH32UKyRxEj1kYNKVa9
1y///Bc923GTe7n+jhlBO5OP4ZUDlxxhQ85x9vrkMdyajh72FYUgrO087ir2CGLq
/Z0QhxRLaF4SN7Z2tuKkMJ+FqJFN6dk9s64FQMdcNfjNyyOpPdmDFULxiUSxnn6Y
sVvur9ebdPIxI+qmMWtQK2mJXnQQa9fRd4LaEMrJlOWZn1el5P2AwvHRlDJlZrot
HLmhFspKQ5yOaIi2kK1DzDjCAQYNNHwlWcUDeYKLor0RCbmoCD1h5vzQ9NINr4rN
PegdY2vUPIM742B0SZBeGRo/ZF+ysOwbJ4+TfBmx0eXSSMczF/hqd6BCBJvvUz9w
0643HnmQJP1x7vjTGSPfPZ02FauC3ba5L3Xsfh23riIr4+lrHJ4MAcwmvtmtraJL
RPChjDHE9OmZvZKyCrNBEm6ZSrYcsL4r4/7nhBU5rCSq7mH0WQG3QmwwiYacxOh1
i2ZzfTWusnl+jG7ASS8YxUYLDTgfU4L1nONEE9wLJd05slpH74KQorQlyV1x7mqK
0ZBbgrr3vbnnhBXZchkB/uGYg56aDmIPgwkHyYglXcBAweAJaVJ/jP5UDZx8KSQ2
shu1kfR/Su2dwpEYuVdpMggDx91kTDNCoO3Ery3QLdSPSk7iD2FjYpcUcbpbPPwM
GCCAIF2Hu4q7SQYb1vFVP2649pwzIjGZ6eFAoEw2HNPvsqy9bKuH4z9WSizyipUv
kOhyCIcMWGkr9LjiN6N00Qbfx9Q2kfmVW0fJ0GRgxOc6v6GzXaEQ2i4gjoRBu+LY
rhuEv9vtkirxYCMurY8h3efY1ESIOajFr+163Y7NKy1B9dZsMZQL67IRB/KAY6vG
WkUIByO4ikN9ZgvmT4Uf/RmnB2KRK1Ko4llZD3NBNNNmemLFF9krPxZhgh4J2xbs
n3Z591AabDPN+wH7GLsFlPnfrNcgwMqfBum2utLPmzMQx20M7y4XI99Gwl1ebObn
CzQLzs0+0tNtVa3Suz08Hih+PT8mgV8cO12PUwgA95AfFu5mb0ctWITRuJGrFLr6
Q2ZHHWMa8zt+IF6Z7wOQ6RJtPCzeZw9ZAs4mO1+llGcBySvf/vlMVYpVRlPiDQmM
uHcu0n7MlIGH/pxFYVJFlVxIJB1FidUcCBJNQFkjFcOZ4TjXWJDbJV9GASQcJLAu
ce2RWfJMHTyUbQPiPfUwrWfZnvLydFi3U5zmHz4i98rt7wBttTNY1D+c7q5wEJCh
xNW7moW4jlEGQ1KT2yZ72PxhT9p2i9FMo3ILMNKZqetoKimXAS7dfAyUDlOHv7J0
pUtC4EZNu0ouNX9t8/GobPas+FVHQebS86E35lb2FPlcPUR+JGvAyKxLqhCopS+m
3CSGSx4AAjXUuHlJq65cu7uw81SZ7SnxVreAIEytIfcV/NuI3ecMjQn4lJ8xR8zy
ElIXApOo0z4f7ao9GvltjlNhaP+J+khQjkGLmbrAHS3iRSIW814t5cM4zxyyQHVS
dzGPH+wZrn+9vql0d0TjoMGlmv1hr1KVXnfBlJE/GHKdgGcGkdAszXdJZYo4P3DW
48hDr2BmLI3lkpWD4YNECR+4cDWvgbdhF91ZtGRdbtjDeZGfLGrxq4vOid/xQDze
ZMHXFmQk3KJAHwS9kmI9MHGtXXkdiTL+bmjvtBIon9AbDw7Pd3ylV5MW9y+vOY7v
1JxV5N+bs4sS4hx9OEcPyMf2ZM7C2BA9LCZhq7eHqyIsfhAdcH/w9CuTxkN8WMbe
MHYNc9WrW+03tqkJHgOR1s/kLigSzcUZreShggLIeM/o3p2YeZWHKir6ne7clcgg
A7w+4BaTxc5VeTd49wfjUQw5pcIOrsXn/A/8S2TB2ttfqiZTKMNUKkztN9gnYL6+
cnPo0JoahVeUCQPIORf/4mBpR5+FE8uuXs/vjnC1ChAnvvXiPdSD7HqTo/kh3T0I
lePSHnPW9N88EYSD8MkyLIDpHA0CgynuxxSdFJhd19y9Yrm9G8FZncdg7o5i1uYW
VyevWcR7ZinZdQKw4kP56cKlfeM6QC7s8JnU4+7+ZJj9uQGAo3+2GCw9KJexicuX
7crFTT6y0ekqUEDztIyv2dL8ZpAE4afNs3QAnsGy8Feflb1ytoZENnNffdNQHfoI
9YDcK0XAdG6mvuovaAzrqAUoiVhIMbSF8ErCPay+Shr95XljtwFMZG/u5oS5QUgD
QpRQcBjsngTS5G65PilmvAVEJklXFBcr2c6/fB3gLGl9FKFAJIkigm0vsOcJpSfg
0tBkCYYiV++rl7G1unYdPT5vYcKce3SXGI4OmHiARW97Ocy252st/UDkSE5zd+FY
hTTyp4b8+3/5S5bYOHDGNwcZhf+jTnQiWJ/LfONH/9eRZxduK+ECPb4+1iIXcrxP
wAMyJuqAgoKExl4/AJWCt3Ox8ZsHbyzFuzvW/n7RqijK0jAb0MHO1WM0ChQCcMzr
Vlz4OYPvl06Q5RhCdu0qLK7g3Dr8z3M0suXrpQgQgMND3+36zROIt4DCE/++E60o
+BDmRO5+GPCo9tQlJpco/NeqWJlFqu0DzKgKGWjE00/kZGCwlVJZx+Sm75ti+8cc
MSN8dC1z+UcOTVoFUOpcJy4Gcl1rcqtS1mUmvH6kT/CSIgDoeGp1wh45ka1h9GEl
K1aR8onMviFHvH4GoZGy+M/7HBNi9oKF5QEmTMjK7aM4GvJNtncaoScMdtKseeMW
VOqo5NrqHKGtXEoLZDSAWwohLxHeNHxTc2qpAtY9ES9PrbD2KxDrKySbfs/7kzzf
E5Drd79YmuB5SLcuBnt1Fs/RenG2MIq6uF7X/MTQQcntU2qzIvXf49aklLk4X6JH
ReTS4x1dZ5faeMqwQaTbmcKKSAXYks8d0uxe13NLbxNNn6P6GZdJ87oYCVpz/7hx
o1ZkdlbgpjHRgaAX+/PYE5ldgGxrE1qWB+KbqxiyGc0ZDu4+sLgPGA+SxQxaAeAQ
+Y4Tg8qOAc2Z41pC4BGe/L+3I+hTwsT6rhEwAU8rfIhzwk7D5YrB6YnkK1GYZYDh
1oH4bxeX5pS3gSzkHx+wMJbBSFrIdKPNOH7+fbjX2wKykixpJd1SsOV3YVQwxeVu
ZOFTmfpjKLXY5c44QlGEf5dSB1gQWpeM//BpZjBlzJ7/VR1jE+BtEDfK6UHkdPV0
+OX/vQhCbgs1YuJvYrW5ZnT4lu/bokbOYbCgu9680p0ExMrUs7mBlmGP+mwBusBM
vreTT5SNifgIMamfa1cd9T9MXn8ErttfmhR+JmE8Y5zYpChb2ehsvuTCp1LCIZKu
sVt/AMICEHC7+l/1F8zUot/yRSYEN659+oc/Pnkk5PC8m+g5/hK0FAuXfq+dXASq
yalUVYgqCJ4iHfcrSoPcuTiWYcKXNKflJNpj80QOQ4Yn4cMKIAc+g3Q7lODicZLb
tgiiIKpNTccyhEvqQGrh6NmO7yQhNMTaTwJi10BYZsaJTQE5CezJbruSJsRs6XJO
GSC/8vyTVMEL1FKRYuDPoSClYGNdWDXnRcRwLCw05lkhOXaQenAZrvdEK6OP6Srn
9cX2b8ooRnjB90xpqh2w2XHPIzaTXx2WsVoDwlgXzDH36luLguVv2rJpePIl06QK
1SC+nAZ/E0GSXrQ6n5p/PzooDoY/38diE4YqmavP6kd+yR3A0Ri9Vq56At43SMwN
Zr2qk5jlKvA71ImlckurRkZdFz3kNTjPA5FvC9g/gNer4HPFCRQ4C9QCZvzRrL4A
suq12qaoMjYF/GzkUEmEV4eQCKs+FP8eDXKR4qhioF41+iMXJ8Ou4KE0iViuXASE
yj8C41yXuXiFa1zORV89dh9TVZaivyjojRPuWS7mARMwScIz0E7PupnlrAe/yr2h
CEnmE7X631+wqibh0PIYJn1lPzyugrHt1wQtj4cBzkJcHEXpftscqhx8V2489Hfl
ln1nRAjvDOBK12yomMKLAhY1liJdmKRLfXs9UQJnDFPdh57pQCiXXMPl5/KwW8we
g5ZCjz34Tp3FZUJUyvjRhF6CHEVrkNx8kVR2CBUPw1hQwuN9RZC8dcOM0/SHAmqv
JZHaAhR+bYyAA06IhSvIUBBZCbInqOH/rMt+vu+uvI22SvrrYmJPZYOLrOLy3+s8
pRElH9zQsCg/2WQ8g6rHjsavkuBo+wjGv07ouSVGrC/0TvE6a1curepoL6MvOlIt
eb1SgUjRgtCsB9RY7uFPiZUiEYjR+H97yZjcYoVRLl0FJB0zx48czu94Jigc1tD0
3wb7JtzUsB2NNdN0k+G8lyEkwx/Zuw3bdiHr9aBz94I9UyrQKZwBxRSdBP7q4odj
3Sac3Rwf6KE1v8slrI8sBrluWj9FdSV0dZBqyZPZR5X3qRNUbiY359gHdPBR5slM
uBqWC+etZnankEEVxb0DhP1ZFsUlATDFA0HvAVUZ4SLZsNn8h1mXuBnD4wZT2jgY
Uhl2PNC3Mbz16+m/24oONDKcE6uwnk6iC877BeNc++LxTYhVREd+67M1Qj712ENQ
gAuuo4MMvNeaydW6sy0N1NHvUkI0zXK76ABrFWLa06j/VL6iMuJVzbhg3JEcFvFK
okA1UNXxLbTSYXDIlFR1v+DDUafs56ra37t+ETd94DKe9UQi98FfchfryRppLLJa
8mb1sspVZUpUt9b+mfuln8vZN7OJnQIyt3GGlsRg+oY3JY1OBT14FdSGaOx7EJvO
MTOjQsa05pF0pfmhJbp3JxErauLHJXJZWPKAFuMvbgEDYTdg86XnxWX49peUkNir
jLFIKyVPegjKFvMOrX9ZQLt3sBvZaDA+yv5DPMk32AUY9nvpAoqEND3pjKGXCgDV
FsTwh7YjuuaSi4QccqCUnKXdIAV33kQNW3JHCrt2WbDRQqdYMXjinQzPddU5PlU4
j55ofVGad3lso2s1YSexKuE8pm4HWu+zNyF12bzO+8PyKreqtYFdFilQmAKzHzAf
hdNpF3WlRjH+3ypt0vUDgjurRwKaDDSbjGq8TcI/EqxAiNRZYA3Z24zJkQcb1Erz
JBChP4M7gdm79g9VTisbPZPDZxIZsN+tqNnrVYK6O834x+coiGZUVscPWjezU8GL
6GF608jjvyO9ShKVEivv6fYhRrkYP3jO1d/oo6ZwHNnciTu+91kSyVLm0jS1tPjx
VXzsRIiitGK0lQlC9ocae+LtJ8ir5Oi0lmDcmYYvrUSKHHKImfli2HF70I8W2H2j
AyI/aonLMDe3liDucqfKivPLlGBdUuTx8ZykVP0wyQ/pKGB9/ox2jjk539ZpYFR+
O7a0YCAwazg+Dqc8Jq0cj6xMxwY1lSJd+94U+f5GFvPlaAUQ4uxttwEYcs43DjpY
FlBv4eq6OZ7pCtW1v/ZxneevTJviag+j7yjhvM1eVmX15lpB3f3yrtguXsVYHA4+
70hU37jtPb1ECS2AxzQYxcPSpuF/Qyx+QHXdn4wN9GQyg1zBZf8LmCCEXGHmH/Rv
YfQa6r+Oe9Aigu9B/CWmkkRssyNSafdNPCqVeWX40hYjAeJIkT2S/351nlxUAkcf
pUaI/Aq86uCUZHsGGOKLtBWbxidQrnLIUSVrax2CHXwiIIhEe6RhA7idBUJSaWXR
yccBbqwFtGdmnS0HjCqNs5T+2kXngqoTnOAYoyVs1Ymxt4OQQZg+uh2OYEE8zfDZ
amVRVvAi8WbrSbnZfnzAv/PcR57gwUPJnHl6Vpa0qL44/7J4uWKD/fqmRoMKcXPd
PdQChRWyEGe7DU6ZubYUcJqMUkR5ELdJd5trqpJYTjKeor7+oosXrvxrXybg6StB
WVM48sOYKkFyK6qOVJYleomwwHeRLjRVHYogaQG5wxQAUdsy3lDSTVi1fXTvKgAB
M8OEKHo3Vsuz65kgXSiSm2Hry7Mfd6VuMco/dmSH/BezpKBoPAPpUxJ5KO1irS2y
zikYGltz1cbX/q3pXM9zq3UHwykokXYi7ItQnMxwQrvQfi4vEKXfneqK3OOcAUC6
rgsAOUtlXnHGyh3wvkBN2qyhequxlVAnbrSDkTcDX3xQXlVy9PrUbimZcyw79JH8
fIHNUeIo2Wa2mwpd5Enp0d2vFBoqdXbcVCLD+QQYw2fONoxVs7lByJVyKTZ+3djY
T+M6LfsEGbcYedgN2axBjp9IBeqi3whicu0Mxac5o/hocmvDu85J/cJ9R+cYyAKW
E5jw4/w5BoVNQ2sXnr2n1Ub7lspVcl3XfVRiXBxD+aZY79uWLJtplAK6XQrZfHMv
uecR6zbIbyhewTyaBPAOaA1PrcBwi7tfECdmIq2c4vUZk/ES/3FHTwdP9dV3yah6
bwh7/g0JivYmgy4cXF8+5C6ASJyEvyyAKwdityEPOHwQ5Tu3oOEGsO7uJ1Is/nS6
qIENFKMYriDo7tWpXamGANTT7WQi/qiXyIBCfjT/7onLTLL92L2qkNGPvB7KLnOS
4Vhw+MvNMmyK4xnKLaaIii+PXGnOd5fgATe97/8LOalH/R7sCktUZHEiKJypSmG4
9hvxGphm8iJ/P5ufM3msdTbgo6pjOFzIGnQhyYWJKHG/NLhriz5M5VrdUauPl7tA
KQBh+2BkZcYFvEyWpAb9GZhC9G7HvyqIzoyvFFh4Tc2xMoDx1LLI7gYRnExhSV0J
Ofs/w2GhbU2dRBchlEfUsKAQvSF+JYXa1MxLf3gm7As6N4dmMuoISvSI9Wvm58rY
6j1boWjyeQAgAdn0SEzztS74rhrU9ZwO+FXfgQjsGmIG1/A0RuhOirPQjWGkpb+v
1aBcY6LVoDCiRXS8Jj8Re2nr8tXy/5xsPelHJynYjYeGePMBDj0jMQmmUtRV//ur
BwSNplFZxadmze96s6QSY4U/Ow3+T7AGHZmwtM5zIU17nBRaiEJuD+uqntpG3zSl
yz0QIRdRApwH/8WPuaVH41J9lGm7/2hnbCFNEhPUv2plfNX9Tlk8HAA7ATvv3b+5
tE+5lIgil6n4/YPcR5M0lPEdcFreY4HpfMiDHvJRVmhavpnWH8UvtnkpmgWujwfL
ElMehUcqkMbT2qcNaMO6X3jCuk5Pj8YhTNXq/JIywGNIqcxCeM3mw9WrXzhW5KWu
tzfGScrMeu6GLDA+BJsguBxdqp7cAIhybd/+yf8NGgfx3fU4Ob9XGUsshqvUGBai
3Oj6CSHICSFDWC42I7ykXj6Yz5LwuZPTkOjPkz8ReobMFxO/AZzsdQo0j20rxiY7
S4LuLcttbVIZLwG3xxKRA9utepj9YFadr4jA2BXbXfK91i+XlMmNa8baWnNdLbcc
QdS3Qyo/oX4CUF2S2ICBbKuUeAGA2c//kOqdIVxugZtlhi+1N1GAQMytkmUtbBom
rnv+MbIdBGZZKPbM8voBquhJFYy6CxopVsSTfGkhKEsLzH8zDAZ50JXlUnhsTw5k
ynY80XWi7AJdst30C2Fs3xHPCV1asmu8AcGioMoKhNPwhD6ne9DePmpBw2yDWiCn
pr9HYKLXVoJNnpwFp1KVREQbpeY7IrlCmHKh2uOxeieq95zGOqQfjo/jzepVDeyO
oK8SvbCyFEeMuRBUPfdJFJn/3FWn/j4MldWUar6PkKKvun3OegfsGJ1mf98bwSAe
uMhOG5ddCbMh2AFvGH3Xi11Jc8qSSTbuRpJ8AAGDzZyX25O1WJ5LJzmpMButj3qq
DR8ZicSr8ac7DaD8m7PJ29u4fmjRaKkSnB+jD+cCEJF9KPqhXUD7wHP616198u7w
WyvV2gPUKmOto+61QLd9wKDU6ZPae4XMW+tmYuNFfOCBmSQtZ6Q6TCZsNGhg3kNY
yYoC92yqitK0aW7HTICjtqiTmpFANVocBEga1wX+Moj7rP+aHF6t0lKj1PrdVq/P
jOd/YbVkFXSH4a+c5wZHMJ/tek1hf4TqZAT2w8OtFW809kPoQ7iXR8/1C40GQrYc
6dRpP71pkT0igMg/KUuIhMk1mn4BLhLzzss0oALEOPJgbPVeTIfCW8oyiQHybPNA
wAMFPRVAbiheK3W1rT77vN9iONTYm7/IAFAXpKJqX6KXogU8W9X1BoQNzcqB3HMQ
GECMR8CKaCp9X4155wfKnNiXZDvZcSAeKgqQd4CmTpCr7OtjXAGES+xIoN6OVRlV
asi5Ck9+Cn6/d7XfMI4o4PW48Ekm2xBXdVRorjrzI/xEsmP0Qs9aJ3Let2J/k+XL
U9gMb38ORmKVPZDGYlbWqoGFk2eebdGHGzbqTQ7eqsDWv2/K6TxdoF0iPcXokqF6
sWd/tEgXPjwpEezMMillAxz2TcuH1mctx5SvXW8+PRRJFSPN2qK77Oj8dXN2U3KD
ZJd71Jh7DZwebzHMLbJdDGiBo7jM5e9ApZOHeaoD0hsdPfai68DOiZzaCAYQiatt
c3JED7A8QODxmVRpTheMo/6haWGJga7EvdnZLqPreU6OBZuhyVxLnoCTo5dffVUi
iHWYtFPptN51AXqdQUJ0UwVNWwCMeMtrq32akOX71BB2DrG611z0l68k65marHRQ
ACVVQ0BZCBTm8pJ8kILcVcBGK++guBjRybywRuFGMzGOTC4AjIeLK+J5Kl5UwQCc
3L8BOzGi9P31idscBeNiCKiUWW4x2h1aa2Uc5iCJTzZezHGj8N1K79ZxahdCBvle
lb0EjuFAxN2DEmV2ND0XQs2FPfpNSdnnZuHOYHndSyU5jeJbDrDt0svaWR3KQ4Kd
3Z4s+czRg1d1/0Vy66wD8UnPaWKkkS0Tdod3nuUngf2Jqk9TX2L92no5REOMqv72
1IloWBA1ay7YiybRq73BsCIZuW9yi1bbxN6ArytK5LWxihCYjTeKvvY52jxlMi+k
8FwGC/xWfuT0N+UJqMpzPUHKMvUjOkwTdCoxxG+4jZ120XSmF8mHmV3zClXd3EeJ
2FUDEyhLnlFR5xmVysyQxkguxM58Z1lMWlLgQraIimOHTRYbFNNxn6b0bJySRD5g
UukGic0t02zSiDe5CJX7oX73UHJsO3W3d9erFReidyKBnL/Ek7PQEWEX3S37vlvr
Y1WIbu6qAbTxtEhZPvOWjeLiATwD9ky9of9pOWVQlbUyw9ZK3vcwSPG9+QJ13MlO
MZoJDbl+YqnH3smOo2XhKGEOnmojzdZPBDO6zGSV/P6UmTCrClfKziUs002xOquo
Ug1hnkqe/Zs6dd8FIF+LrsNiaEQZSY0SZz44UQA8ZB/tXJFyS12xIEBjyaWUsR09
W+XBElXpL128O/B1mT2Y9HLh0NeHkT7ItfDqauzNpLcs2Zh4gvOvB6wYNMpVaZb4
mDIq4cVQrQ9fUl4TFtA0nG77Ek1rCxaWr0iDMM78A3TRC7tG1vKNsws2UhHGJhUu
bn4b+YScxg+UT+Mr4a6zgZdjUNY+KVDEsYpP6Q23nlfwwaouvywnaL7+2HHh6ZJb
Ph3WCE2ZlfmwL1NbZCE3IDGHrZZFeZIyReBIAbRpzVX2Tgp/a9A864qQWJEHTi1x
vTC1JdS7CSPevUB285J0Yr9OxHKHTR+nNwBmJJUQODvqd1VDb2Aq9cnOz4GC8yW6
Iioadb4i6LvkcWyBpEKetA02sgeL3wIQnZhRHcgdU/WEbPiRGogx5AdbBuemW/dR
J8QOk5Pv0oCXEJ9cTyw9oDS4wo5lPwsAlYnb/EsxrGSi1lmMjyai+lzW93s6Wz0y
NoonGKv7D3t2HvcbO4XbBpXoZnX4p6QsldP3Nm8+VoXbAVxfqx34mFELvWpQhtHb
/zwnOlB0BcOxOAnlgg3vZMV93tMOd23nelHRE2jk56w+bseoJHFvfAmicIu1ucKO
l4ynmwacEvDvzpqif2F8QsEbbv4KKPwQi+92UMDv2LS0sctRAkbttPijTtVfq5Tq
NKp15DqEISjTFVC8nzwxX11sYehqYbrpX5weuJ3Z6PJhACELSDUeqB1lszMupMui
kQ+cuNcpDv7QlDveUHpAzi4EBaF5MVUwekKqNesWT7wqqzfVQ7wfGd3smAzccUuh
pLSly1LBaZBFOf4V36CQkfNX+kmDs90sicPmX2Vaptf6AevLjKhVhSBb+/BS9B1X
epPxoGoSt4ffGKj/3034OHM+hZtydtF/3FT9txtw5ZkW5bpmYruGsukqfK75qCHd
/GRRN8RVoPmrFcR6/CSpJJ/s77hNz31/1QXpkbz0sccHulPlvfmiZwZoXEdNcUcN
r9uDo3eD/lZryWEN+xiD+xzszHn8x/Iw8b6IemDSLh2YYxZ3A0ar1mr+OY2TA629
fMGqtfOivQhVXyz8iwPk95Xm37G5RfmWeZUy2tZHvtLP9Inxvfvcuhqw8W828RS8
adgMIcu1JGJs1E6EZcEmtpgCA/ozl9QumIN25ckueWHEpfZIt8gnIljC+4Af8dR0
9ujEQUU7Yxu1BMpp59RgZ94MicCx+x59hwh+/hpnB2ab6sOYueK/MnpzC6hCYmPB
f/IDMg9KsXSG9wSDrOUBz+UmQ/ouHY48FoEVIlDOF9lIhpnOi4F5fAutUXgnVfeo
KMErTd4QMV80Pm/ZLvaOWCH+Rsz/9HuL/DICUDzzzO+bkcCiX5BGKfiBYK99CNH2
Xa8CZMGKjMA0yhHTYjsAfUR+jWj5tBrvdRuto6KywgKUhP5jUAuGGfbpru/Vi+MW
DNjURS174ZLt4f1+eG/3o9zTFwAd4ojVEUBJKKhXI90rNZq17jHJfj1JD8wuufy1
BFQR9oVIBLj/ki+nVQIYDf0reibYtW4L9hpCB8RMAfbiprs1db9IUt82UMdSwHzg
82n0w11pbQ5/qej7k4ak+AgQbS42AdVSSe1MVCkSG8lYi3nmAE71zT/9EqfmXsNT
8jsa43HvAH75XFkV/AEMTeW8ZVbln91byUyKuTlTQZijUsoS62S6n0LI81MIl8RM
PfjzGg2xAvC7c9XvdCI/nq3dpOkVqxuEuVUovC1tRe1Wh5QJf0i4KzvPd87wzKEH
e90BAgCWbWjfiS9GXV6CehvN/+4MZA9ajz9ZIo3UGnZv+aq85j2W9b1AdY4N+JXw
WqnbQmX2GzcCq7rqXAjwm3llpP6frrkhsSwjNlVG3/p5oc3edTinte6js3+NKoHs
3YZH7dLxOBH3uI4bvchwPiHyC3fMwhcMU5zyLpM2S2GE0s66CjtqpO0ZJ4zmi8ux
JXdD+AD2Bf2G907lo4SQDNv+Yp9NJbPlxXouFYXdSVrbbztcGkutT+h9hqz8dm2z
EZuoFelyw8LCKgxwotunfYNwlqcrkkSHoxW1E/HQvlo16LSWbwVuOGa3+ORrpl3o
6vZS9ceV+sNBGIW5Dizve7jZ13KyvAoAjnWX85Fltujc4IACGE7awE8k7LWrrScR
alQB5MtPWFtJ/gw+iuG+IkGpJPO4AKI5rB7ajxXtSjMtAARil0M5GkUkZGTsl63W
0MKgFhNTFYtt/tRdXJmUr4oCBmI2i8PI9iGMWmS7LycW4tsjVG8Yy904Dj5MxOqZ
C7qoWiggkwZWz+h4T/tO/uj9DNcMR0OTOTN5p9yGketKQIW+Ex4KE0bfUJ2ryJg/
jOIeJY64sBJ990mitn+yBmRiznwtcX4nNWRYB37ePYdj0+uJ9ru8A27Ep+47wEq9
emO7NVs6NdvGstc7XQHu8aFCcpZHLYqk4vv3W3LQa47B/NsMNcbhWuUepd00llTY
1s7dTaiMbCdwzp8x2lwOCYQ1H+xz0yzqTdWRUKAKFWpaO56ceuBHbNEwrPxMpgDv
36WuPGR5aADbdfoNvtSew+MA3bzOGScLs+V9gN1GBslie3KhAtwWR4DOgkc0BcU3
gW+teUTHHnfEFObu98iB3KyGOn/IVZNV1BsKv3Oiy8XmbvbIwLWcvsHMeAsmatEV
hIpd213cctiVgr9pVKhh7X1q6vABVx1jKKXHHKQf22AS3MpUPK2IXzvIBE1zSZ/L
z25m4dJH5dmG2kDH0vZSNlA/Dp0BWI+4qHQXHqA5YUSxY/kB21HBKVYAjIToG1Mn
zKukGdrDAic0cYdo8KZaH1g2A8TpWywWooRb4IKUnZIHp5A8xUnGdPJLYZDDmoWC
mjNYaDTqjMH4WYeD/p/6Ijp/M52D1OiaYTy7zYAS/5S2KHKou3NMOnWwI61w82iz
Lkbulg218tzNsYUEw/peYtnE6MP1yXG4yYm8c0lDkSKblLLczf5nnWLoEUFnxpMi
ZCjQ84E39M083pFYmEt2GLtz3BO8i4TRI6bp2VQif78buX0Gs2EALoIIhOlCRd1O
svs7zlmC7AgrTpwNoNLvQ2gvf8QSxVfY0eZWzl31A8T0jwqjFEIgMpz8jc68roTS
bUC889yT17leZdATIuFmGDS8l3UZeR0LzXB0iWP98Mu2A/+0WeJ3CC9shlp9dQsr
v1YePdXfrtSg9PUM3/BDQJR2MkuJQ4GXj+o/v9Wv8RTV5nargYdUm2XC2JsZM7Xj
l2bCCAhb80aaDBf3r6aKZgaM+j6hoJ6geT9rMVtQSc8hIYqhntD/QItGap+bf1mR
UPYcgmlGzZpNgfhJQW56g23ithdF+w+NVhvFBVcPByKD0cz9ArvVcLjALZVeBCeL
o5QAstPKeU8Tq7gEzmgn4zRm/C+tKG7zdDWC2Xn3iL3FmqPvvo1HG8bh3810qZNC
85Q8PobwvH6c85jrKWW4aOmup6Yljs9fHbGOZ63xQpGdqDcwi2WRapu0QiLqjsAj
OwHeSUWaz4soPuvlZokqx9wYr89210cJywHHetMHHDyMaOwKNqogu6AxqPZqbdgv
jXXokjtJx6dLNO5aug9w3jRXVJS90hlk7uUlbYyGJIwzuG1GzQo/csTIz8TrZT0C
TeZzQf0WngZzhVN+xMso4vxJdV9fZW+VVQ75C9++l+DdBOwxjkGgTSTYqxvQuzif
6NMj7c9hemtwWQjnELD3UBvMS8B28wn3/Z8cJV6XQxThed84DJmZ2qaDnh9J8CDq
PtWTGbjtIHsZBtdr92Jd+gqBTryrec7FXqtJgbSnZ6HZMHCAXA+EkjjGqSVALqCN
UH+fTqyEDlyhWqJhrJXh7USoL8KBYXYC4TwLLBDrSCou+O7/sBTV5uO+qHZLBrDl
HbHDc6YrNzVqNzYv3a7wQIbkGiETKJVUmsIg7KXucX3zzMjjoOqeJYS1H+vxgUtG
8LI91e8tHaq0eMsJitOvxE75x69JhCA3ATpvKTpcmYqaWgJlVuHX+omzNlwWkPJX
AVR3KVmYleqiwvasxU7t3YGcqymfDaAFwKdE9P5dFo0p5yoyeiqft97ez/TR92Kv
LlRLQD2866bM2smRFgLE3HJy1nfRio3ZCYvu9qyxNucqek33Vswae03jm7XO1oiO
pJF3V82SV797ets1XJONcOmjmRckWk2Ybv2FCmz0oNpIA/rhJpZqXbN/m9Hl+od8
YJ3sH4AcRQ0Z9tiN/KSA7ylHhcBr4c9hJE9DE2A11cynkBdu1eqS3esPBBbjF1bg
0Gp2DqQwTjIaR5kRMUs8CUOx6Xl4eLdOTIkTgEUOz1DasnRj2vLes1x2TRYFDRvl
waglgzx8HLuDH6OVPtFddYq4unHdI0+eakeEsPIfFvxH6pFSyU/uJOxg1/K5VXL2
uajJH7vASJm7UMORxEDDXrtfkgbmb1ZIKhFDyAoewAdbM6htrA1+Z0PlB5oasS48
AgFi5Psw8xEDAyGX5lQVWFnB53bOldZMZV6snbGtWuNkK0pHqZ0QpvoBVrSVE4QR
2SF3OnTnxrIIS3OKR5yyv65GIj24W80O2GSmWojDVvWMBpWFNhkADb76nNl0lXTz
qQl8NRLou86M2Euod8L4/OyTXs3eX5aKNRPLjuO8aiTk1Z+gqwq47mBvCwZJ927y
mJzhwXN3B7JUUQLW+DuGSyryrsnnnTypcuhfApm5bDm9R35MNJP9QR8tkUmRgRLZ
aM/b8rw0prdSyaFmzc80QPcDi4VcTBEf8rDlDpJKTBeqMPTILKwsxaEWxoF9tTAM
zJ3tJj31y21NmR2jNw34wsDZ8YTAR/RaDlUlZKHQ17WzNrJ0QOSeIv7EYQ08DvNq
N5KX40A6zbZsJzGBB+CWS7K/wC/+KcAviGYPBSWAegeUogjHqUA7t5H9QVIOPTGa
gDrJ+G2qTBwcT/yb8gPEwVtVR5RFgncROJNppTylVUKitabgRJrAtOWAAN0a2n0R
BSGOVqwj+ARrfg760ivx1OMK+qxVC3BkV8SnPttjOoNhMt3GQzc6nqTS5kLtRd2J
+lV+KRJ50HBN8BIgnV5N/TZDlbkPEQVuYkAJ4JbLYZH/DwGU8nFTNx771NB0b8MJ
vq6IQB6CVuhagzzYaSF0lWOllQ463LJxBEgsvbFYgsqv43IXClTYqt8oMCwlhmAz
sQtsWnBvhyHMSdTs7rqHGgf+rIMSG3Ze3nUeriLEj56mhMpxjJsOkFDFUelrCUt8
hvQUD9ENxyyPdtXrHdE5IyMiqfNDd3Q7QlMsalbznlhSnj26TRqckspMSsozy0Dx
7oHjcu3SaG61ZqbMCdUfF5rcZ9R0t8Acd2ZwFX2uMzrLBdCtEH+Qkg5sgq9ZXDMP
4e1BmRUIk/xJGjYPcY4/wy3zewVFpANV2EmVPOp8+Q+p7AcJxK7F5YyZiiU2Pt5h
Q1Cd9Pu/MMdGgpxxJqxD2cXLYpfHbHGgLI1YW84/UjM/EysbG32G2ZerIlPZxCSD
kTgzWVZHlBBhlgfoaQtypcSCjpJgKSf1d5TYZxsTNaTRjpjFucXr/UDWbZsZtnfu
IQU3zNBnrVtLUId1toWERnlkLIWTYFJ31sYYr+JDM2ASpcoDNA/ggp6ZJcbju/nE
rI1hy+97/7T4hbvhfjMK/F5xgwMZtDJFhGe6oqp7DWhbnNwU1hDQoQDNV/RX1oAZ
vx2y2/LOVACcTM2nGMnTSrqUFxPVr56wZzMQuZcTc/JVVEhxMu7fRkCaCiSfCVaY
OjMXUYcIwwIOuALRSmvSchiXavG2jQ4T6rv5mI+h/QbQO095AHPYW+fhi6NxlUoK
+Pv1H3IW2G1qGYDDiiv9zzAX0BhU9CgTtyA+stRqHkH1g/jsWyXvnfNlHri5IP6J
qrlvNo9iGaYxzcB5W7u/JJF7lpQ0EyVCf2/bCBcJnOGTQcNHZdDzFhTSK3zRWVq0
jtBabfQ0cvUgbOb5fTcPhcfmhNy+LjUCETNCj8Pj7sGSKcem+268DflC0uFtEcYv
yPES4PmPv2QQpUtfkdCgHCOat27zNx6+NnBzwkErqtStaA9yX5gwKOPH+xUYey79
mysYAlcjc4lUsBXXcjvX+3U4ZCMlRU/EwoLeFgwlAle5pzvGf654DXL6yg2yQCfv
+zlpjVDOtgYxLnuxaUh8pSb5y4U6yOC2vgjJO3JmM4LFxR0LFRuZjRk9iSQRXu1/
WyA8A6H/o3YDY1vAQWZbhZuLB0TcSqxEBKMNbBvkedrdFxGBqqSCFvrMZoPLrJc5
aLLDeey/6qAgsgAHQqOikVlaygKinuYfTna6N9If0ELvavMxqWZKglkWeXy8lPhc
oDKj4lYrUU+ezndQsTblFt+0CrjJQ3Y9/WeCyzU1JKTSifzavi6B4AWKuj7A0Ly0
x9JyHQc5rNnNm4Y8HU7lGngNudqAFu6wG+ODE4UuNw8Wl9G+mgSZBwthYGeQXwHX
sorqsIKortc3D19sJb98nBtjlnHmxuvKQVwvCvaKw+J3Os6MawcfaOuds7WhKcLj
VFnT6G7lbwP10bpx5JebHTryFCtSPAQzcy37dbqhuafAqUIUSoWaSCwQoSfmnsjc
i0mjmp05M74NnTPTui1qg33ex1Zu0Hddw7DBuqNcJW+fp/jxUpE6qq5UGT/06yIz
dBPmsSqGMakPF/xLGgDX4sy8x5hgTDlf/ClBF6V99FajAU8Z9xY2G0wK3i8Ck4RH
PVsGEq6nuCSUu4CieosP2cRiH6v8Oyb5OSaHOQJAh4r0Tm7Saj1eFnOo93CuKpDQ
LH1IoPB4u75mpHg7q5aKurn3y48kpKa/Rhqori76S3kY4CR7+YrBb+yhGr+u1MRt
/4woFqes7DF8M7pthyvOzgvwRiUeSyxw0dWmsGlfHUkT1YlMfiJ5cnBezVQiw6wm
ci0293aovUT+62tvPzgIlUngArDz9JTIzm+8f0Eqw9LVtOVSD7akLFN4zEIJBM8t
nukNC8dqJBuhd84x+kW8eGfvO1EH8vDQmuSYeQm4fy6aamNnM93wAzP7EKMoU9V9
a/lm4Fcfkwclfjjcq9haj6DcaqWWMHFXpsloDF9gUICxVzJDBBjtML41ZhShPClR
r8DanfIpAvEtepL/SMBLQFS5iYk3ob8ugstDNr9KXhQKyMXeLxEKEdHocQDppRZr
XbANXBfPrUmVt01vToRbwDKg9xx4MlOai1uVd1w+t4pw1XkfCailOCkwoS8eqm49
gAcx1OqwqT4OSMijp5zCtRkxVlcwDJNTT0+lXopzPJ6gTJoI5Ew4WWdI3yShPVHG
YdUWz6XDu8uapzl078F7iS+bO7N2NiN4x+Ezh5DcTOnTpnXVtK2PQE0pWOFbVTzJ
/yY08rxNwRgfy2nB8rgQxPUeFEXzgNBQqHdPyapsJaIrrDzjVMD2oMLBO356P68S
58mh6/HprbDlHtScnoaGIg7Dj+5rk3QOVQMKYJovs+JDPeXUTyhke7oUIeIuetXY
Az1EtGwMdw8l9xDlVe7zpUtF7OSmKsJ+EjVskmPwP4X84sXpr1I3CeqzP036Tdll
ONIXl+ojREQ3cmvRFqZXW+p2rCH+JwKv/OFz98Y8+5f5A9xTWbEOqRt2JRZSmqqm
poe8EBC4hF9kcpuUbYLce2C1pxPyaxqetwABFt9JSfXs4VI9QV8FTDPcpOP0RiN2
p/hdVeIwTCoLSkiYZEDjItcDKRnBImDabmANI0UWvG+qN16C3e6vffEVX/AmVMYi
jJJ51jRJFe10yi5+M1RWsut2n8jjFSQFfc6qb9POY3hn7AX95OpV4OuEDelSrD8o
Tqhex1naCPPIBLDWCD8TI80bfkE6R88hhegm3o2tHI//5vYDlJrlpPpr1p+V7lpS
9VRtLoh5fQnPs8nb+2i2yyzlUaPo+ovCbrWWHQLsIy3G49KavXCERyUI/1bwd0iE
QeUbrQC6+lzY4oK37BaH6kcWoQhvjyvsVnzN2briZtNXmjYpsvOTCuQb3YHgyG1N
NotfN9fJzn2npQkThEtntCo7BB5JFWNqIYmQXwQGOaz/8CgjL4ZGMLRi6nBgBoK2
tVl54XQCvDMgedoKxHHQ8UQg7QCQB3aN36FxdQw84N4C9X2KrUYVbZ53znwZcQv9
zC8IWJCt0v+ntkiMEn1LfTvxUrlyLVAUS0W2m/h67z8Fm+Tpwnd0QysVd7k0zXX8
CcgLUn9cAucxJSf6IRwMGmXa8Hh9BDpUEGM4HVeUX9fryQOrEL2EAz/8LpF0jM41
/UrfJbJi117zchvFFj6BHqXM4BYENAsUMd0onbmgs6FKkkdqz/qqdNTOurqY38rl
lye5yCmytHO1hje6Keb/m+MgnG5zC4FwKSao/EgtLJRxcXhg2j/qrYqoZOvoOK8S
rm6r3RhPuLAkkxj1xtvWawr7Sic/KIdv5LBO5f3wxLalXWxVOh2K/ra/RRWg7WTe
b+t6Myru7CSPGIZTGPNs60g2iUknFk5+OoguX8RTe5u3z0oqfiCG59x0QBGp5txS
FLr8xOknHOn+9AzT5K6P1h55B13bNelWNB5EON4iYwkia8jol1KJtNb+LebUj8Js
Vur0hYtMRr9fgbNRhFAXEyZURkBDXpUg71PGIPWt0gqc1ym2yjf3Cv+EXKpWl+2i
x2NuEhcGMUPkeyzpED96NS4L0SGkjErou/lGxbakLEHc363FIaNnfMdRJUJ+VrSc
l0eSRzx+PV+XZTZhNJgsdvSJasZi8UtmTyhgAWrpH/v3jR6c8PQzmKy41ng61dHM
dqvUACDwAXN52Y9HnbRvDC9YS6ibtm1LJgYug/FHlES29y0hlkY28SJckBFcFxDi
z3pDtSPqTrZCLNpJaSmPFIky+IUgjkr/eB7FGADY64dkS96hDvhbKyMwPftUSqrP
EaitkF7mMBxr5TedE43jwJy4GN417YdhaB7bIOGP6i3cPCRdBMIbTRvkYxnGV9QO
sVyGfUlEFj9CQ/9bN27l97QJ+3vgzKt7/UFRzqKn5XDcQeEUfJWNWWXJCtnFvz2l
o5b1gxcruUqkQGyeB/wH/+AS49siIwp5ERe+wS+SzKSlv82S032epXWM1Z1720va
otF87rybVESQv6MVSlZyNk/L81WTVJhiZDcdjB/TuTkjcX5fxS6oFnH6fxTYEIr1
DJOgcZdrBz0A380b2qsOU47IG8mt1kO/kftDII4ztUxNBROzFroRBTYjFrUVNy8e
PaYwA5UW5Zb81BWTNJ2+GmtxYs+w6DBPNB15EvMdl4XgDPNj3m+0SaA8Pzi7hp6S
ypmudP6ikQVQ/5GQ632RbRUnA65QA72tqu5yyplWPWqoQcb9xm6WSJCmCNhXL6r8
jUD61cXw1+lKnrAxHCwg4EosA3gOMq2WmkV+GARXb0wZEJBt1Wi0GGycOPKxmF5H
46bNWGt0fnnF9aJjNitUwXeiAW+gzSHu+zMP7lmPnaLvFMPerYasstBBIQip0gRJ
zverhto6gqISY9KEploFpfFNpBhNHCW0nHXI/huoI2r7dwkfh8vAKGMbnr6Mx/oN
s/T9EyTdKifg6HWIE9izP5RksuROMQlJf5biQGqVzbymHhhaLho5cv8zFgZ51AwN
A8AWm9iZLxNT/bvM4g5FARCVeebhgzdgUX7dkwMwUGgDs4Iycm4Hrx/oo6g5OJX2
6UHvhJm/8rwpwhOaoRMI80DC5Ct4m5KMo5WpgKNpjSux0LRl3BsXKqmQ4hokgPNg
tUrAsTJrjY4y+E3Av+TyInbrS3LWd6xnFU17TCgl4hZYy0wVYx0Lul6MaQgq2QkC
oHFJZUm6mYjGr4ZTSIFo/SiFg7rb6gT1ONhHRgdIy40Hl8lKkayrjD2OcwGIyQtX
BwbC9y1KnI/5Ta6LKw08neFz5vRA9ZLipB+w6g2EcxDVm8rsY3aTpV/92vMODgk3
fo6nlS5sPaxg6+5WLLys/aLFX32FFq/yOU0q9LJlNCzR1RyHQCAIj5NB4IjH9cTB
mxibuKyW5JqDlsr1K1puK7tMTM3ux6ouCXZn4Iswc9qXC5WVsSGCDq7ATgy8Q+eA
Io7JK2CV+153ivxNAbqcho+iQVfQLU5NL1F4p7DHW0M10LO7YEpG+uLC/8OOjZ5Y
NITJVpaFJf1HIQAx3fzTcLGM4we8OUV6PLqjcdomTupWqh8SB9NNQxF+gTCmqns/
tgiIOecif+x2jyFyzrJ0Q6yItoI2jigZJ5MRhowkTHGlO7fGdJ58naHPhlerwlVb
UsxgMp4g6s/YTnVgLrK5r6wqNLnc7Xr80NkJjJDzcI0PpJ6A4wc8y+ZAno2JP8b8
ePNXwkIZ5eUzZ6oRsViBgj73bg/a+pSBTbtCEUN58qAwevcJF4QaKanKcVkB3iZn
5JXVTscdO3du0AHPD3JBL9LdjdGgLTv78R+cH/KihIQidlGRg3HiyzfiWpP97L9c
hMCMBryothD5m3KAKkzOKHLSVuzkErQJCjcQWLUGb4TQhKEpmM+W81Rtnf6IFf6X
+EBJC0v7dbh3HAhX70YGBHV6UiME1rof0CZOZ5M32u1jSzGZaNP4vStOLn/7anog
MD3r+A38wJbjWxGomqN2ne4HO+ldpt/XMFq2C7VvlA8VcW9/v/rQxsjFBchA1oY1
XbzMdr9NyeNRxQwbz95cM37EXT3KzwPx494rrQ4i2uouv/CXO60IwGSkUBh8bXsb
xkYb9JDGQGVeCa4cfrK+LM2Mx7FIMCNOzcvz8t4un2ZT/rgQVgJFYe0MSUMdXMQu
ms5THdf6QoSJXPclnLJFYsDwDQe3Bq7duyDtB0tbD1+oGoPd+aZkY4B38L4zAYVF
D37k/mYQ0bqqyNTzXwQr7Bq+haRsSvrqQc5vhmzBwyp4QacVNuqe9FgTbQDR0lSl
JBuH6YGnlyfO/iZGVgBCGqx1bcZYU7HKTQnSG3jDCQTe9fdo8fdODI7ymNQ1m9Jw
/QWA+QmXm3VcRTchptpFJNVQZ3g+YK3fcVw7WA3ZDmfD+QuDFZikz+4wgBk+PFKI
FObgy/+7EpS2KHrxKEvuNmGrnRdQNIfSNn56KmQJ7HcBTzaMHcbXxP7acHlRySh+
wJXI427r8f1Sj4fhvirHyIq+Satq/NlqOhhnOeVLBl70jBYB3utEHEKCB64xAI6+
cnCI3friJfjUVA0GSDthRfrfp/mIZM48HtrhMEbRgxeWkikhovyKCwbBW4SmuTYD
8g33zontQYPYv0BgwSQEcZ47UadGIfSstgLBfZ9l9NufYDaaBOJKzo2n52G5oVuz
+jb6GqhhehBE6MKKLXR1enNCogXRG6+kNrqQLBIl0FGiRAFyiLCKEvKgteJ4Vgbn
8c6YAC2DWolK0/fa2b8h1+Omq56e4i2oPOLa4/Y6yCnLcE2+oYBA0rfGs7EzpXqT
RDOAuSS62BCU0HJ42GnpL2XUx5XJc/+V8eE3IJzuTaEKrOdmbkk6ei/Lbggk5KbU
hDHSlL0TRpts7DjvqlonOWAF8W6TnxoWBKWPoQg7MhQc/oV68g5G1T8QdJFyq3Y2
RpUeKC2haDi7d6QSZL/gM/YVbSAb6J/8+KwGI85e6aCzM31nVdlYVscfmszhw1nl
mxWLVu9VlG4AsMnEuJXoyiRbNTj6Ok5n/wxVgRQ50cqUQKZWluutC/Skc4jlZEGp
wfAwtSoEYIxF3MWGd9OM54VY1hIjgyerr4A6CGlNrzfjX7jzHb1riLp3GwnAZuap
aJ8tgVUalC2mu972y01vahP7PHuLR88T57oVUvdT63OT4Vp6KYkJTXOL5I7gwvGP
7/nnwSbVdOBtmAD7rb2DF0SV3j0Ofev2ZWDvAJph7/wQvl4HjA67U9d+sQ7CXwdn
DdWNpTFCmPIPs19q3Q6YQx0A5xMcpUWPxaNcsDmacwXfzjDgwv6xr7QTLJ65xwd6
YjXoUJ4ULGNyTCiXx/g3YKpslsMkCjncDx22MhmOdM/pfajLvBH8cCOiEFQamN7l
/SHtfw4bd32rRAXoysPQ107XrOPVWIRAbkHQBfvLXuTNvrVePUzijapePKQmz5NZ
0NhdRkN1N1bs2Nj+cGrO3rtFhIKsfkjYsUGM4gW4VAqmSYcm2IsJgmcsDSf23pbw
wq7povX9oj6T4tjZLIJGLZ154rmSxiO+V2noe0INmAwalirRBnMlcEn9Ruw8R9Fa
brL4b+A+Gx75CRLgf+AeEAPSi67EYDWysxSm8AX/TRWM9s+k4nZwZ7wYqkuMmHZ6
quVdd3my+69Kqb/xgKgRJ3BWYxpB5OO9x938jcFMOImHJadopZCp4ULMkUXDMdpJ
F1RHBpwsINd1wPKJpvBdOg9sDA4IiOWZkz64kml7FqhTPQDRSOu2UwFz1v896FBm
QP8+Xl3x87F0nLSdbANCFHpJsyz6vNw3bJelduR8PQ2RbO8Yl42R3pnpYw6G2OtL
rPO/uKflmmscxEGYSe4KwjhBOB1nYmIhgCneQxQUdbmgU+ubWyxm/Aj96rzks2Jw
73X2Y8CfdSOUH3PSiFVwm39ThsY/oEAyWsveilQMHldNVTEcV3r26Z83tQuWsZxJ
VEnbbmOKdjLyMm66DYdQDJkpRsrvbZCpql08xSXwk4tG/GmgOSa7XIsxJgBPeh+h
vtZ2343Mmjia24n9PVhBUeWdbN3ZF9yOuv3isTnScB40s9z9ZpfLP0OaJcCQT0CY
83EglqQWrelA6qS1wZoJRpNU0qMLQX0WEW6hZCHVuU6onE5HqQSfk/4BZJhImZWr
8/eD4xRz2aTTZpZGSSuTraltxTOyRbW5q/LoI9qauQG9Fw8uJ6987VQ7szJfijo6
JhGPTyqFZ9dbn3oQztQf87ANpsfs7rP3HBEpBMoa1CPFb1okaHXoJXCueOybxadA
fXmkkzVsKHlggzjn4ygKqnn/db1LeOle6lZxMPxIzgLYlv2NRdDEsm5kNh0HdthH
kcQm8d4Z3f4YILbKGFkKC3PGXD5MRwfHziCyiVBFpK/uMmbMEWfXjDAnuwwqnp6d
SFbaE3qy2adx7mbWglzPZ19oNsOsfbKNoEcp2YIo+nT/SoPK8X5CeuJ+M7Y1Ye7E
fy/pqeX6xJS2zzvWpAVoosVfe0ysN1gfRfYnZOKnTVe0jwE/197KrHnrncqRqN6T
9JFtbeNF+TI9mOiZiVxO46hmwaqFNatkiCVaQrcbBtFdgg1jcvyjhPGhhZDv0dUp
tzBxw3ES2rwrDHukilZjyV9SpYs8yezGmTQoUSGgCrP2af8s8G1JARSei7IOfVBI
C8qZs9/TWm2VShUPpb3HJCZS0DoUz0EHh6pfKM9iqhFpUJpHv0OCpRrk1UcfwdI1
sKXbZTVrfctHRpCbKDj50DSMzb41Ldzrn39TnPp0Kg6pAEaylhItNX9OK8Q/t3zS
I/t5bA0ZAb8JGv7CkPNvFIe7DvTvIq4SxnMwW6SHXiFNy6+NRKTB+mLzg1XUBGK2
sAU8SpwsDXQ1drmO4/27YsXOljFWV7wVOcFMmWVb17iNLvUhzXUWV1aIenbdi3ul
/lLPae6lkoFpfgnzGnoat+XYhAa/BJAC4LtABsljF5cAA/eI25kvVEFFx03OuUk0
bR65Ag9ANMh0xhLqWH2JcxJ9tv5/9GtbAurRZRiRQ8a3JfGb7ir1aVzJmlOYdgZa
qvbJrlp1fskdsREk8bgkTruanq7I705NBR4lPsGJnh2F/DD9EHQonzNS7peXjDxX
wzBDFkLL9vDdsqLDUG5bOJpIza9O1Ae5/NsMx0O40wW80VjD3RojhBd0HPXiTxqF
YZ8nbuwRQKfgLKmeYwSCImJfGWtkwo2PQ6fujc9mghdRPlmehomuh63I2SbkUt3A
/AnHXX+6piCO6v0vXyMso0ODY3OQTXxvdN5oJ2H93KBa4rHZmbT6LWJHiZ5qSQqD
mfpFrjsIhMa+lp7xg+gieesgaSVkHvk5TqNHaxnxO436JwocQfuyczx9GXq+NvHF
v37OSn00t64XEjEjHqMVbnZkOC5VBeNIZxctb1KH7hJPOVJqTVGVJUvee0HPDwuE
xmlKoI2M8ETSMorOGJKl6OAy7VJa+bDFZI9BKsOFCgAIf9hocl3XcqNWdxykZ2Ec
bKMlQ6vAc6qAxJmdNzgr2Ipe2HCmaKY6EvpxNRgQHFbnqHsvilV7YRC3IuOxDQOH
oUz29RNTY0Ll1ghrkpU0mlLpGVCTxsbESfc1rztuX7TTsjBm9n4/eKHfVHZDCHap
PRzHbSVTK0kyDnXVjhjUE1bgJWo0eDxOLoG2F7e5pLBAbbGUijQJ8MCNdRE8yebb
pY3/Xuw+k9e2Uck0dvWpXQFi8mRdqj0wwnZxUpseXOki5mlRrkxSBh9R2gg4hHGR
8l5Nn6B1lVCjRm1cXQ0XkDJ4M4uRQDXoplSee2a2kIVXK2pT7opTB2Dc68qIo14n
BvCsMuxf0z8iIUxbHtOCvnjVWr8Uihe0RvFDr0/PMvCNGl5XnuPJAhwDdU8Vc4I9
OvbogzJ5zwABvF8pgDWp7JPhRqbItEJ/0xw0pBqw98UGDZFe3t9t3Zpm8YKZNymb
Ea2nrPB9rcKbt237G7FlorARrSB/+IggLcKndH+IQg81gABIQulHVPyMvcOZ8axl
HBC5m21TGmB/fAnwSs9qbtwA5eb0tPrXDXdJgOosGT7xd0tGKgQDa9mE3uHEPMS5
jp+UYx232Au5sRk9aKbv/NrndVrNDZnnnBnUH9PCnpds76BOKKsRy4NW/kiZanUL
eMv9qO1zWxUvu65wWlnFQfwXnPGYBa1mAUSRoG2cOJn0wf523hyULQGAGJajolyP
aI1h7XX+M44UHmbvNdLcP5JkuxqUtK4Fw+ENW/DsXHmSmTk8G1U50YCvKZIWiAZb
FzaWKUwQuvsBpympiF7Nu2xPizJvAUezuT05CFNqzXOXnD6NARWtXsMgglB+y+Fz
1O9qhKDWf8t0MgBfaD7hCz0LeKS/YCs35qv2jETsbbPJq3tUmOLwHISHrkJka8Xm
ljKVlgQOsehsZK2EQvBM09VwtxvSUqB8FDfJDH58NyuPRTW7/katWyYN5F1vV/ZY
uVMTiydkxqTrjk+NM21Qvxl5NEUaLd0y+8p7W9nb9WXQrKN6iRtapy8Wk2ho36fb
OMn9l6mjwA6Pk8dM1FqIagY/bUBrZAgCgpmjJaloh7LHH64Msh1iIL+9gtHev3/P
Bv5k4yfIOoFbHmQcXgBXgFJ2BLL5qUMbv023KV01yAF8+HRfPQw8f2WcxsU3zGHq
eUYfS4tJxnz++G8R0eAMV4lz8ZfR3gm4OvcJy98usXPaUojaOWAlLFwnYHoDN0wa
4vDYripVunEkqisdONq6f/yylUWTW41FhSDPxDQ2M1aB6oMGjcyOofqiDbrO0g93
eXs36/werCrohq1FSjpdE5J6VkLrlZdzh6iHkosG7vLtRIrY0Erpjb4wkW0kjolH
UodIcDZHaQFxsvFLFKJArrjLIgHzxOXgMRTr8ec0CkxUF5wAqkFgbfc0fEYRHa1I
oDGbp3ybEeMA9+HHnrj3lViVxS0FM/MglGPKEvkt9Yi3JagC7SBRZxQ/eoi/XqyL
nL9K/iIIo79gOvI6uRRvQgLlUsMzvPCCdx5IDZJEVwOu1L2TZ57xm6/OazLsaygz
/9rf+cZ8/xmpgDPxMmXuU2V20jFrOdGix+2+1l798Kfhy0gxu7yCKT0BT0ayGSWf
06b9KgCqdu949IZQsMe+s67ay8TaxrDXK6RCDOhb2mKkmkxMf3dzQXSMAp2eOsy/
UDumS/4ghbVVHfj+JOyGLTnhfzN//lR5gXyiwJ+ta7GE/6Hf4Rjd9a615b/xyBW+
xO1ADbA+DbUuOx/xLX83RXOB3SNK8EuKx1Yghi3st1mfmNIWhledjjKr+n53xr7y
sS86o0ehp5TBY01RlyljcmVBlZ50DkFgORFG0IHY6xrEz2aizqeHjZUBR9Fuj/i3
ELobCtJFbAzK3TWBEAbaii4ctv8S30Aw4QvKeVE6KfuZ4LSnG2zsZJzW0Ggqx97L
3CmRtRNNWTT7eiyFJGjqnfvY4cca5Nhnqk3bebfHIyYdUdAvfhSOQxXHSBEbkrZw
t2bz2U5XRdX0SZC7hpCS0t0SMVZjz9TqpKKURGxeEHuY0BfyPvDBGp/lcL0CeKhQ
zcV6lV20hRzCwdcvub96OOfv+A53JKM0vtJGfkgO+h58utse0djqfvN7WL/mQ7D4
+dUH0IDIcbPedTw8fBzMCb/CYU+8xqO83kWeIRACxR+EJee2bXESVN1ql+G3nQvf
O6keQNFCtmk6cMcGrK4mLCaODuw4oZRzL8UofYzJrIySultMZFQgdDCcv7MbnC86
04kVQIbJ9nzQRJEb8jK7Fa1oWgpsHhZvTAizNUCE6NXD7BO6GiLQ5qidzfHZ5osJ
4FCOuvzy3TL2B0LnCzx5h4EyxgfxN0lv1YmVNqt0EMthVaRFrjDHJwBeaNNOlbmr
+geaNV6ZgKWBbr6PVwUd6fHYjlUG64thdpDIUwdR9Jglo1/8BzkOmjkNtv1iSVm+
sbWqFOIroVovZBpctLJ3MGBdWX4PJFMyAkpPJob5nkallD+DlwAKmC43nEvK8K+D
PLQ2zegxd/DkdqbFkBoZ7/ZUXLFGfnw/9kPlziR7bHnY0UMbcBmpI/4HLgkNwewa
jgNizPt5sDi970x32znVQtFCnci2jERy8PQzcbn2EzEyL5szrBwUBj3IDGoxXZub
BMYo5ZPtxpExNB3c/I5WjFW71A6y83tQRyRdxtN2J+pp4TSjbll0hOB0Bp0lkjYw
Y9vVf35KTDuiCm8O7tvAXfMkLIMZGw5ODRI1sIOL3EZ+26g5Mp0nsgOkERsRkIdH
PVo8+ZRG55r5VxuQ7VnGa1mG8fXCE31qRWhMBMijI2IgC+TyYNIPSY5+ith7ZBwU
uixuUjFDJJ+l6e7/reo0g6ZddfNKFwGHfp7hGOyhwloQFRRCHyF2QjCNpQ8WK2qa
vb1AziqYjU1uQjt3cpfjQxqlabiQw+lBnTjD80k6YEWgKPXGkUgb88gJO2N7P18k
qpzj4WO8pcJ8M4rrhJnpe2L6gfViCQ89jtqYgRCsc0usNFo81xsf9iNqAnIKpCs2
dpUfYcEa41MXHgp+SQ6eXgXwHbrA4lONOmA/a8rfViSDPIAlJ4GlIaxTbGyvFWjW
gBnILPH05Bn3uB9XCHLrNZnPE9lYjqLZPkDHEapbQOQMcQC+3FPohkGQHj/qsR+O
jCRa8p42qy+o0QvuGBUUUTVx+S+ndRsU/wY1/5Lo+vvf9eCsiNUc8XpfH9MsoX/m
yerXuN1Nitd+q3uIh5gKTQPKOel88KmJxma/5QnGDj+PMgwGHXJT7V3NvrXuaZje
rnkxpgfBWXjBc3IRaszDpMz80x/XEZrDcGIoj4WPY8V0uwMr5HfKhv/wWScteLUp
XDWZ5UK1C6cyvzr/hImus5R/CrhO0ns3vOlF1T7NN5hnEctYnmvfZR8gGG40nVu5
owH695AjObr4LvgRqvMHhNfzPk1UktoSEExwhBdHu1uvoRf3IrfZwqVWd1A+LgfQ
gEiTqA2LkAHlNX0LZcp0/HbktEdyKZ32qZTlZFENK+8XRHtlPOVRh1nUccs9be2v
vbw1pzGFgPOCjDy/UMxnMeJ7wnpMJLF2huqFawCXcY3IdjvP6/uVnxyZrIZOclDO
IflME8aeqLb+tNxoyOpB6hNXaF9vlE58riWCq5ODjih+sO2S3LrfrPqGziKBdWEo
VqW6+w5s0SfK+dgXjxKHqscjiRpgUcWrmU/I7nsB43X4E3pOrahFmIrr9/U3x1us
5SmGceYJtfef2XEutRTtbgvUOhakAhU4mDiCTpoeCCux9sDvcZbUWyoJVlcUvgg0
Zl25TfnPI5ZtHp88VYodn2ICnwJAXgmjh12GR95iNIAnLHlMjT2WHwZWWEA6snfB
M1gzC4+oFe11kB0YdRmEbdRo5Q8jHe7/FftXbKLy0lx6iI5i66F86rY1rjVzatOV
LXqITwkoeT9iGroxvOJ4VVe4/QqJIUzoxM5dhVnp5+NW24Oq3DlHVm/qr+edPa1O
bH5YYYbPMODLPtMbwYh9/+kH/7yvUe6kmw9459TsBFlugBcYIH6sd9ukDniDF8Tb
9q5DdUruxawnLyzpnMF2l9jlkaewlo/M0Eg0QLYdSCqdMw1yz79xJUx9QtouTMuN
jIQGYUs4cPCPHgtbcewkeQhIyLt2U1taX1XJEiRCzTih6ICN1mIPx8K6/ET33tor
EYwDa5W0k4NGDAMDdDR4ddehbAoTs3D+Mdf5nLbo5lXJ+Gnx/bsGiKjXilEekyRx
kP0AkXBuyLe5UWoaNFt/2DLoUjjwEMRYc0NQBsLe+wAGeIkrufyaCdIojagyg1D6
GlNcYLPmanAHDPvw/7ehpanWQUr4bk5M47Kg3NhK7cpR9R2D7m23ls+GIeQH5F5S
tG8L7wVSUTPnjl7XDn/74KktSWvEpU51xl4yUuUyUz81jyW68R7TXJHFRNS9Narv
AU7y/v6Qecu958kuxhAE5UzC0pB1EdUXA5AkrSXWhhWL6+zRx5O7kN2ZG3aeg/WW
MuNWsp8bbgL1404/1XZuVZCIeNmZVOi8EQqJE4UrjzF9x6E96mUtIG4UVcAPUkBT
auKz/S6yU/EfALRt0jfR53FfFS5nLSqv2e+QrCTUyuDZHirws20BL3z7nBpVw+SM
wS6c+tiDYj8mvpmjB0PQ7mfZkgJoYFGzCT54TBTfh3rZ71tRdhG8VFaHSApg/tnG
Vm377dFdX8iosKj7OcSc516kKxNDrWkw2QJ6F1GUnbC1B7Mo1vn3n+rIuAiZIV9P
+UQpt7Vrbupj+7HspQPfZwUN5otLDjKJ3DojZFWXrJdCT+LQjcRjw/xrovzW//hS
oobypAyL5JTkb5lzD8uz6E1CKEb1C/6cRB46WOHxyv821kxfA7EkSKh8KwZDEvK5
LQBYlfiBB/r2bk1Zbdl5yd+gzoszapS7MrCcCAf6diMZMQECVAmVm7JZQrkD34B6
oud4jFxpKA/VyV3pxaHu8X9V5G0ireC5gScISGcyXQVvIhPkrwxpmuELAyAwX9CI
t89Lvo8GkrUjdIv8prZvmXqxK1OKcZ0pjbvPCZ299iFWvdM/OGZ+YqrKwirf1Q3u
uplsnzEhCR3gm0pcS/LzwDyvI2JepQlBK+0VUbQ3hKKhRD8WvgZzJucFWlUsr4gg
zqTD8fnzA+l+3seAu76S0V93d9jzp4bSNtv1ICZXkWOrtuB4fv5bki8gnLRb8Uag
aSOPYCo/Su+UO1zOY5vLTYBGE0XcyB49D3vIwxmyOiVLKwRMKMuL6B3CCEXHi2Uy
W9GVF9rXnT7xVBL1xbnZkyAAWr+/Nrn1bidvqAk5vEEr58tk9lnBnaKP3BpgzVEM
35i/NlZ4RPD9otcKx5vrW9LyJ7B1upPQkM8aqED+/6K3a2ohNJ3Md1aperr5Fqy4
W6IM/WzQzvV1BTetRWGw6doPuP5G8OA35UEVW8K2NS6W+2/O69rmcNqa4aFTK40z
Nj02rtN8Jf9oPbMFYDClw9CtsnoGXIwZ1YGyWJwpY9YtI39K8XyrMOpsL0gif/x4
Yh1J+nXI6ACabDBcZqCSGNllZlPRS3fLu468RcgpZbWPuAf0VulRSn3/hC3UsiL/
Zfx3itIH6iH+8Huqgt3lThhsNe8n+6ATuB/cVlrejAGbIEkgFs6ES15eXXD/YK8Q
SNOoToW65ybvCmgX6TGPwYb/lEv4DFdpGAbXSh4bco8PLOZmLR+sPCDaAio8gFra
du4ApaE221VZQlbKhfWbQJHv+klE6UFdlDQM/6wUmllURFpRyQJjnsWNwYrDt3sn
mDBsM4el4mWCUlIgj0tir5HxpDo/qJuH78WhNZWhHbx08CpWrAPIS5TGx/Nkw3wM
0vpFBnv5T0Flgs8vMK+ZsPCqfiFhgl2pkXP3gpBOUoVs6OwBtmqvyHfMk5SMOQvE
SPTsfgdIxefkXAeuHxgt7sq5clilPHpmP6zuq36WvXh1mvwUJSrTURFzyHmAlzq2
WlNPC0hTVt1gM556dR7Q+5pZWlOT5QXpGohX31JG3mi3+NWFA6I/MOJ+eRnwklnE
vvDMtdrTR5aKvIy7ID9I3nle41tMQCY+QieBSI8FJFzqD1S+DYFL91z8oQ6+k0FQ
JvZb8zCbDrsLnMJBsNts8KNKM9BmvGA7AeVw7J1PH8dPnlk2DbhwpVYZOxCLG1ZL
TpTN4YLdWD+ZT8WG+axISgaamX0L9tVIDEEUalpay4jvDSD/ZMqYq0IQpdwfWJOy
bFG9z4MZOk5QF0ox2PjEyK7NJSQlcifwywCJ6M0/tkLjSTk8/II8k2Wsp7F3zchz
MQiUdDq7R1nQ3if9i82Z29hJ7NXvh/r3aqFR0nkbLk41GX032ogkak8Okyqlpq6U
klieBjOFFE5d0zmYPsH3Pu9VagXF5dpZnz6WKQ8klPIycI1kD81jgDw+lcWL6c/k
GjHoGzOsJ8SEIS1jmXnBD7XDoUS4MqiNtWZcgeAoF/6FqwzeByWdBB4qRSurdsLr
29YV/6c709f/ik+n7pGj0PxkK27SBJC/Z1Ng6u5yNMvjNYFqm8aglCojprfbBaHv
H/ySloa6uao5LWxMuAaWhL93nh4xVdudQLCBtTLpQrIyhqCCNVmvB91qDJwC/pft
UPsvUV3kgvebrsLUDXpKv/uPHPWqwtHXiwcl12YLKd/e1cYQq7MrqJ2NyRVFnRGV
OFRQc/xFnnvHtoHrCyiZVNqQOgJ195+MExYblzIfgGmoY+UDi7wYufvjet7zOZKy
PBaBhcj6QAL6Fzw76BrCW+TX7bkdVdVT3IufGb2FmkCCFzRDv8ECRg0ZYlt3k4D1
X61wVKafdkXNSvGXG0zps48CSLjIFK2OdpbO1s8wGC8UPuHdubcfwF7PIC68uJgs
gmNKu+/ri85Z9dS5puXrfPm+08v5V1+OSvKBFHx/yept2KzYIUgG4BrJruN+St9C
wn7y2/FKQx4Uu78ZVcqKWkBI1fF08ix7qYnFX/PVZxXy3FZMGOt7AfihCYrv2oRs
/xHImPe2LtscI029YW+ojabbPfQsH8vZ6wWD1dpDUhHyxnEh3qazIG2qzGwljgHV
4knAKuNQvDpXSO9Zbwn5nK1eYhEN3OSeQb48k+T1BkZeuwX/8pcSTlB+a3SYha93
cCBzW76SLzrJAouPy7jpX+6JdVXuyUXHjun947ANOXyO8w/vztSoajvzW6rumNcD
gPfAmb7ZPOXVuBya3KoyJkRoqkqD7tJou+aXN+a9J6L54MKYIYGxfy+aKY0gXlFV
vIF22J0EERQwMavEYWoVNI/HPwwJPfLj4VgPaI8i+0Xa6jjiBxsVM4d2IbPY2VGq
svP53BAFxIEi/vBhTtIYBApsqrE3ES9myh0gqUNOlWYNyOX1demGkhqjkP0yRv+k
VT9HhqkMIorZhle951cttwdq7T41qakQckXXYFzbSQrWIP8IYuXUJWlcHeUBy4J5
rEhPntQHX6d1iJPJV1TUjJzSLmjNh+cPpdtjNF4ZhPtGOV94jdYbQFbrwVt1l8OX
2/UCS5kDvN7DyqJJ+JhLGLkW9XitPSzI77Bm2CzZM57rdEL1dAERL0NpVEtbDE48
9PhL5Bgwi9uBWA3YHLRiRLAMh9x5aDhzo9wJ1YdLdibjMxlkCDn/lZT1eOAZKx/w
4F8EFNY5d02sDzHSo6wBM/WlN2ARbdCq3VUPYtpZg73y3n1/gXCIFgEB3kdqYsFu
fn3128WOi2MLhbhsPIlOKIF1WX9z+LvEdG2x8fwexxbE4HrzP+a1KqpIxaw3Fh7l
RNr8HnMRbDmo38cdeYhi02R+VKlYlxMa23twvxsiqZCikY5hr151o7fhZinJ347f
zxt2d782Fwvo3I5qfRXFVVi8jf2MHUQcf4G7AhxKrcRSPV+Ug3znL8I3jbDocgtp
1XIXESxbuyjUdtktZ3BJo/4FPaNua34ZZztFH/LzI5qF//+XwCgWmKphq/WFhGSl
/LBn6JmjXTQ+/tsMNTGUX4jiVCzidVNffGYnkTmx07VzrdqR8CwCuULRykGhwblT
ppMG2nTeUheTq7lkzfn1aOhloCVM4LM0MfAbieAkgEVAfp46QGEMy8x2X+b0Bi0e
SUmDuAi5LeTADttsDwfNpEwBSusuTC7syQyDPgVSVuIZxPQ5Q9eLIucCTv1DuIGs
MiXDVBjnyZy4S5am14N60+VGUbhdxGkLIFzi9VsCB7f7n+s9D/TiFl9oh0PAGSRg
HYve+ZLriVPY+HiDFSvYbpc9Zhv5tzW2fhwDDbgvULW2L1IAKFivxPTA+q57U7jg
VivPVEax/op9UNPJV3LHMDdiudY8NNQnNYdkDrCh1v2b7K8gTaU6A02w+nVgrQBL
Jl0UWVrAszV4+SQhasgaRNaqXf7+aJR8Qe+iJnt9wDuz9BDvxL8CJlFRlTpulbCb
wMXnspyGd00sfGRB4KYW0phxC0R9tRQXuKZ/m1qtso6eTmkIoPwR/FOATREQmsQg
MaNmpZj2A7VIRJfmIZ9Jfu019vrcCkBftqI1byZZAzukcz5XOZcNs8Ova3C61Mf5
geP1Wq6kJ/vGmMRS7NMWOfuMuwZAhUtkUeyWQX7bEXkb+rXZzC+xf32/AZCwVhd6
dG5sl0lV2EpTjmRh9B5haR/i8w1MhqgUdtX3bGcr/Gq5cJ7XXR3mrIRijevqrmED
MuqHM+Axr7HWvS9I2oLgdJmaEA3p08C/NkoqjOpvKH2bcOe361DfL3xqfIGCZvT/
7uUnpCsALyZHJDTC09jJJNvHVyOhNp2YlgxhP7OF7Mi1fzvfds5q/cIPyxf3CiyY
wKcQWO3Uis9lbo5WzKYS6zWyU6UkhAmOwyzOWGAbA8v1VSl9CrLMzfxxFn+/aFrE
FP86oHND68jI8dWgyLKe5eKYk78e0ZEpKDSY5e/GUUXMe3aMQ8TqKPK2/KJBtekj
PTGE9vJGZ3uTbruMb5goIHHymsaNzktky8GQeiBGBivvGzzXgFOeZWAlG1cEJvMw
y14nsK1eEzO2LTcMhmxT4120G0ZskQRHNIjJ5NeKtpezyN73mrOp/i3oAcLvtsXq
PbgcU+IKO+DmuWLgVUIUKhUYCD5M1Qd9f7yxyYgl+36bZghdUCieEAqokhFc8EJZ
5pQ/4w+dLvLag1Ra61t9pvbYRceAcw+7f+4+fOZEMcOz15iQg/BdoonBSr0CrrG2
xAbSG7NMK/i4fNSXw4BQlabajnYGZhXXDYifltoasOBkSpF3P3TDpTW9GFoXxp1y
VL+fldgwIQwx/8UyI6H/XrO5e9xgfBsvvAtgnav5Jsbusin++g1aKnMb7mI2TppK
Ol9I8iJD4QsPXBjUA+nQkai+dPO2Gjv8j+rB68DI9iBChQhp14mnrnCQxa/DbYE1
T7gFRTrAQW8BzLPJcxZjw2McbL2K601Wsm9bqvph1AsoosR5fDaeckLiQfqcpNfQ
Z9sq3sNy5+OoPyP43VZ2F8xkpY5g7FmvkIyro3GlvkXrB2WcSPAVrcOtJ/bMiNSF
0/3fMfZj3OBovi9VeNCu1OZKDARb9HrKFQjCyIT1eUX7dWbk1Ykx2VRctsa/+SIs
u+hgCS2kPu077VcpMwl8L+88vJVWwbM9VDtAiTqM1Y7UJVMIPtUudlPPXMQBpRaX
MLAt/ceNie0WEgO4s27VLqVsCuiLf2QevDV6ruAJY83EzEgvlLzzx+8uY4CzEzEm
zlg6TteLNQ5OcIMz+O/ma6FLTz6ykEG1VF4UAC1wUaT4ksJx2DIAzFiFMNWM4K0O
mtJ9uSMGivCHO+NurBzpUReX7/+zWDJ7Mu1+nZxF+JCdXq1wuBCw7zfU1aarCZRL
S/vXESsbKeGcdGnsvZ59wwb3u2xEZbMSfuH+R7aiHKDhVsK2Nb/7yGpxEuhqijPN
IuU/jcQ0j4bClOm/mD5CYPdMJUeTWctDxwvxkPl2ejy2QRY4o5a07J6Eq6IOqHwO
ZHKLuF909LP9uArJWS1hrCV0bCVMNwT9AkLyExxUpl8sRgrCbHBHX7gXXr08PFLF
WipNldENxrSj8uayM/kf+WlUjyegfHzvJCC2xNDupmh2V3uakOvRK7t1Y5W8Z7FM
SqVB1Rja7Mngc38ogi2liqPJjaI2mKKugPlwhdKS528ROsuxCyH5MvkES6lM2IKC
yHiN1JecsNTcu0FCZPjPGuEdn1meZy2mLHCOmYwq9qRwcS+TDbfQ3OsSWLSMmqzB
I0Msyznv7Sis+k2/dNn6PsyNPk4RsdAaZoooRrW/JNGxkwkqL2RsWHIgYfNurml0
hrxOHWFychtm6f4X4UnfoGVKMN7yZ+bKzmp255Ps5OoW1bCkxAuNP4SpYtLq/zO/
HyvICgmS5AK2emvmuhDTHymlOs6sYbFbmf2IK3FhaYw5tuT6hVc670lDNTGzggtW
7A9iKjpgsOt1aCM/Hjl3FfgbRfZJDXO9LrwqRStTPxkHhDInrplfgI15/KUcyXID
EC2hOawOE/iVntOzzQYXIjATW6EePnJb3DG5avwB+ALs7I332KbkOBdpdQdd00Ux
FnWsDWNTJp1fsAynh70STa3sKispazIwojcd3EyHQ4jSXuWBSrZPjsIb24dnvUXt
O3hPiIiP/wtHC2N2QNX+Yf/EbzytF+9y462pr0JcKEJ+wD4TD+tZhGTHZiwRYc62
wW74Slw69Q5AIA6mkatHh9W1G1Y+5V3e5utPE8Az4FxH8bJQ7f3lD+p2TKvEZoAR
2H3pXbwiTcsbQ6pdiYIeasz39QpXLVDHph3Cyf0G9DW0uCh4EuBjh47sLgSl3Y81
JH7HwogTepT71xyYFEhqqtSsuFMo1dJjb6JMRITloilrxbvTXuOr1LC9MYpu4L3j
ryQ8hTqGX9UPO8rv63d3Z+rf0OVWX9iJ9/SG0XRPJg/uFbquuSiaKXLT0W8ntKFI
COAX/CWqNSglj2SUgWXk34PdXd29DHhuuw9EcOTHBvL1PXzd7eNO7i+jaycbF7iA
b1EH+wdxGL3HCZHMLRlX/Hjblrkkpv1sZ3kYAZIpD/x92gzGJsPYK1wH0eouoF1l
o5t/dCOkLt99F2mgKDS4TcfYoT8k7OzK5QgQ/yW3rQA/QPrRC6qJDc6HPkXHujXl
rSxF3QknARcxQAPtewKTh1LJwAhF31vA3tEbCwnwQGG3BNHUreFKmt/EMsFqQyQF
H70FzZJGlj4NhMkgmhUQA+ncwVk8M+72aN0eTA7NVUPTwWeQd+GE+NIXDuHfzCPo
UI1MauERb2RfblZkfclpuqaw5ougoeXvlrShKgdJN3HBjpIkWHztyYTMFacWcLA+
3Tkf8BONy9j6hIknEUNjJQ3Wub4FJDDjnY+yPQtizUQmIDKa4AvIyjXGsVUrTHCk
veHbUIS/e/tn3gniN63iAPIGDNVhLamW15Oz6pA15Vr9nPNjLZ84AWr6Li9PK7lx
HzeSfpO1nQjqr5LOP225XEoLox/qpYL6cBs05MNQ3maKUE/5vgNLlXSJFP/wrS/B
FuGE/BY1raalxrX3sqw9g5rTNLrX2Ltdgxlq2Gx7B1YEMafSBseuVHIfRhNmESRA
WKfOL8JfxmCgZTM6t1Wx3c+n9v150d/rnJ2h0aVe67M5Q/t3gdhOxXeausZ2aTFz
we4uZG9FhSoLtVSKmgiHfZTHG3vtw46kHRAZ4/rR8gzIOfs+RljTNGn+qkRn4WkS
6GpsPOIGMoWAWCvAig7nLNLXuVatDXyKvQ2JdX/oq0ZhkopX1If1bxVpqO0Ok8nt
scBYwUHBiJukDT9RF9WIn8pxX2XTabK5+rFlOXdYpz/G1DQ+pROxUQk3s/t1D0dX
r6qyU3cM9gUkWGBPtvAg8p6m0zRmT1tpwW40L7diO/kMw+NpqZncnhQ5+G379mh/
QxtEJBbHxzmVzKN3L3xGcbtC15ixOETyUzW2H24n0qUCLl9dZdG0eqAXxsjoGEQt
X/zGG+A+uVI02j9SSO7iI2F1rNbO62HzH+9Oxhupq/YAlWXxUxdZYm1/TcXfR+F7
88fjQHUwCOhRQlHApsYunl/3KMzv0FzcQuLVKvol2kQypSVendshQXpvGzAqiOjo
7NUuxD4c/VHZiPs1XmzIuWIzJmeLe9a5GT8Xp2JRIex6pRx/+mlDTiTcVX0zHwdL
/6iJdl3GFKQd2LFoWxXEB33IYeCHN/74Fs6P0X4Qlh89qVy0VK87hkI5QT6uAQ6g
OnD0IlK9DiO+txp6PkHACrLN6r6nq+ZgJVMBNkha2ZfHr5Z5wv4WBm7pbKnRHfcm
112SB8yTrQ7rssBcm/D1Wyhg5mgj+iqSq+UZwIKquJGZObMegy8FLGjZE/naozF8
bIJn0oOeMmGB/GPw0kHD5s+hRI9kcq6APHUeqUUKVjoz9GMjRn0TyzD05QLKIULS
p6lKLFRNVpbmNnmZKgZJf5J/nz14m5Xj7hc7mZRUViw9SeBfi6sX9NvWfiKpsVl6
wKn/B+1Gsw0R8tXpLKniZAKnWlu2+Be0SC9lPb3ItEs+vEUumSfFMfTqH0k59yHb
b8zTV69iEOp15fsSgEb2QY3aT4gRMROChtl/UmkYvFfKo5AWDJtn15N4a1ouTXAF
FqHdQBQSEBm1S1IBqBy8yR2xmG/kFdrQG7utao82sdeOt4stUYD99pMMri1+1r8l
va1qilyzDVfpJ0nuov0KuPyCB6nBqVU63aK4+8P3Q0KbmbeiGSHAKic5epEDz/8m
8JGYu+9jfSYvUiyg4vUwABkSMW0IoOx0LzrLV/xviN1gY6UJqCmqEv4qcbRNLQ9e
dXmWaONXeg5dfyiJ3bZU/N3/uVtRURUNy2vfhzpBYOkaw27U3AturbPeyR3G1OB8
60XrUNc7RLvjlVQU/3ZrJqiUQgW89qrAJEMO1xj61pBxp1RG7aToZg11Jw4hklYl
WVKLdbgyFzsB8S4yr+WIBSVR9cWTLL4rv+A27DUMXoJHddlS+TjjSQjJ2/7MCgQT
xQfDeRGZM+nbvvm5/zrAb5e7ExsqDajkP5WS2tm6KrlLpod5eaCJA4ePax/3nzxS
IlHDVdVox5w3Q0mdmOkhvg8tjYH0oN2oBO4eu4aK1K0Grk37hyqjOszM7pcVTup+
zDbsZojBkxS/O38PJ8LTewPDE7vDiiUA4KvcIRVj4RMTtB/+U44UNQj2q3aI5vmB
cxouoZj+1fqdFP+CQLWYKh66/oyJDL8tzhbxrzCIX9VbY8BDjj6WL6k7iIxYYUNY
npd9OsFj0ayU5kcWTFcqsQAyA98xpEL3FEyY/fLXBBxbT0pAThKvJuaAuADIEDgc
aSNhG7URxxDwrloHxaQHuxcCNTYQkkiIeQGzg929GdennrFLquVjW/tBiggYHSom
WbESgXfLtrMSR0jmLctfDbU4/xPoL+EscIcyQTiKsynQOWWI6ctOTGsO1nHNE1B1
oio6HbtFjDXX+jvtpe2mlYV+RFbGnZYhDBC9cg/DPlS43qzsDcGqtexwKhVAu50o
SS5Asgmn/iAWDy5WPg0RAjV8bTL205464z0YP4ok/ELSr884Sc31/ACi9LwWOmlz
itD2a9h2z1abd9i5+lM70P1BDiFL0g4ZOwGlWNDZWeNiMHhtmLXRU3gux6lDgKYY
I/E3Ssk6LO//o3QkaFdwP9ByISPXEnPKBdacfFlOJq5Us/eERpP819dV367YqWb+
MTAvKLiu2D+3MQyyQQOl8/xZhColi0z95jJBV8n9Y6rEO69n6df5pA9ACj6NpPaC
ev+O69LyMch19Imn1om6gsyPXn7HFVTT0tvQubqcTdsnPbJDzBFs+C0Gq7wxgFez
2SlXY/qWwWeLMqbFjGW0pFDvelBM+vWPGS25ql7qlq7Gb1QJ2j9aUeW2n5+vGQr/
gTpVvsTdNXjRmK6xmaNFzKpQeseHKYzwrtIQKpQkKLCArRxs3wgOJwHdtuAWMRsk
dB/yw8ZRohiruu3orfW+/gNayc+0t+VJZ38oEF8Bps+Np5vIEOIL68YkqYDYFDfB
kGXPKZ9VoyXypSYoKMtxQMpkIQF59g2POECTUNQOOH4yBErsMTewIcrrSBszzyg+
B64dQz43s4lhslPQF6PYXSiejgI3Ek/trUWm9nndLJWFlEelhDes1s/La37Yu0YB
7aPdOJntetYaCkFTdWxkz2p8lKIhEUK7uiW6ookq5J0i+B0cPi1aj75x2Vi5lgHy
oUyfLMKbxPVJSKWPycxLfRRRFzcUQWu+GIXSu1H8O6vAY8wM4H1TQ2Px4Tmuakt2
NFKnvDJSmHk2mK/2R4IyDCcK7xI1uSbmqV0Rmpmk76hAvorjhtcBUl8CprNcy06S
TAVzQzdoBUCkRFaY99EdpVT2b9ZQR8GbRRVJTLpVVBbf+9YSGrifnrIEyRmHX4jz
fWRY0/793+L4P3FAA9744r6IkuofTABqlPqq17HOa8AK2mxiC5x8KP+spD2O8Y+y
tDAkI5sGF0uBLbkKb0wku6M1ogc9fCSpYY8qSFLYX/PPM3o8Qm1k08otvHnZ6ZBk
VYW1eeuLA87YyflABiJ6x0EEZSiyAUG2aniSZGRqflUxpt5Mzx899g4+FNj5yaT2
+5K3BMst83Ds9fpSTcKDSENGP4W/D1VesR+CkydmiuNPFlRtMmrDt3yc67uYXUMi
FQkvMScNk5DYQoSj9idlkKcBDZmA59mCfS08xzhl+0jMwjl6ekErmfZyYdzb1obx
xyTWnnVztLUn4av8wCnJ6bgt1IxO9C9FokID/Q9G4dM6MqiBEwq8UWUeprfnOHg6
4ROIKc2aVzZblEvfa+AX8y/Z9P/kMscqSNRJs+YC+ZyvvmbgQPJ/fZQwp095FSXR
+Pq96SoDAQ5snr9WLlAeBMuqo3kqbv3AuPj3ZuzRsUIjI80vOp4NmC9hvUoFFVZ6
5BrYla1J4Vx1mLlH7JkQfX8nh4B65rUPWqF4jgqjaVCHvy1d1/4LwCErRzs4UZHi
EOm2FJSXvLHNpeIWiOLIYNV0CIqaJoMi+RcanxTKj42OIDdBJXunwSF7grn8cbKq
MZURYh1aZmVAtBCqOH4hFOx21AR2s6a/Z9ch1wa26EgTs/c1T2Q8/u5NmBm24TLW
QlUueuWzk3a3sYWtWxpj3H38DMgOkmXKukVZtMnDRagaxlrWPFQZ5v9Jf3VcZ/z3
raEtMI+FmuJCI9MTH9SRBVjGnh1bFIOOGsRN2WO/0VzZTTjedDLY1A4Fav2Sxuwj
kLVJAsLIVKXz02KKZpOYNwv+wk6CxzhJwXEXe59Z4M83x0hp0ZWcAcBZeOEIlVoG
SGYC5DgSZDHNiKh7/X/NHzHE0183ryu1rDIXqSYdDeC+OnJ1cekKTUZNTFwpdLG+
LIcv70hJyl9wHgYuHzG/MIyCZSHvKbTpakTMPszyebkizxPnom9jhB/fNXo783e/
1wQcJ/i7dAyy0beezY1ny2kfqtUphWAoiHbE9xWlHIfy8jA9XKJPCrdcRHd597UN
/MTfl+pTFcdrk20nh7aWXIqBsQXBPUcYiwgLFW8DmkhNHbnG90lS4v+tLMoMCUsv
T4eY84yMNMmjWBRzkeV4cnq/h3FhYxWvD5bGXPk1aVxad0xTuthW2sVD4RimP59l
0y0m/MEi0k6XAyVQoVQDQQRcQmfChjblPZORrzOJvk3UpEQt6PoxYB+DdXAFvsMr
4fotFMzxDcXiy3AK5QLA5uaPWeY+V25+VheN39JLIOjFI169I/Qvj/VbVrhfdxJZ
j4Q9Wxe4bCZs0ezo8UViuky1FG4Hv72wrSB2PMYWrVskWNnWA6QSYAkzwT9ERO2G
liXy1xLKiYMiCq3rOLtVb8RsLFSGev5NPx+2ngCQlgkwjfpyEXBzR3X2xo4hHmm8
x2kP2zvnOOiJ/lVn3aiNlsbjO3d3yRrck5vinpExv8FmtCj1qTmjYidgadcfRy4R
xtQYiIuV+OCwC7fOBrXByMYXS3QvFoFenqq+Gj6sgMT1XzuRvxxjDOzXrnEmrG5N
doj9KVZNJtH/TleMWNu1dNXT9XXTjMk3R9cV4QJ/4ak4js+ZeVfEX4ua545SLG6r
vBAUpTA/Sx73oj7AN4zf3RYe5wB61E1XoUGvqb+upx0ziDd13rGTymklLpSj8SS1
0xlg77XUcH9/XQX/nSYdTkFEafapM5H5X7blINuQdtDmc1/99nvwEtHlsHW/4Pzl
pwa7rRLMl3DTgm0z0m+NqFSwZ5q7L20mImuzIHO+zz0Y9GxKkoehuyc24aBkXUIa
dgOaZB8wxegmDDMnf+lhUPFbGfq3/95tyd1YayqIw4Dg+j8EvWA/+EW7MmsKAJXz
AhPEpBwGmOuz2vV9n68Q2747pt9NT86kT99IaBVrFzuU4Ne0Qy9tnDtyAUMYxebP
jFxnC/Jlnc6B1ZLX7xUFMSF+OVgOuWxQWEkVX18kvyjohDp4eEE6G6getF1+lcXb
aDfdM1JqkjuoveJioeV35bP74z0dzeEfxyFcdV6oao0Dy4r/WeYoS/+w+l622MuX
kGmy1YC07Z+Pyxkfh9gV/vSCXjxhOriZIBctBaVEwcpkltDNEJKjXWcy3YLx9vEk
A9Fz01FJxisXZmQbjwpYQlKk2YxcRhYg6/YL5UJF/mBF/siATC3pX1ZsEyGe8E3G
46S+gqw+7v8xSPXMKFDCTqGlkLVsszbxaSntC2GCWshUaGpGMp7oqeS++kKy5Lbw
0TOsDp6jE/6nx8GcWNiVDWW4RZ266XZyY4RE6TsQuJgVnleluB4OACtNnIs/sErg
8XDYjPOl7mNyz+OZvWJDMiaxt9HHrrx/hEXQK0daPyqD8q0mprTkP+C7QxlqQx+1
LxtrC/lUAt0mOHqHsu3OAoKNMjMX4pC8wfQYWJX1GcbehWSVFSTt8Qcme1L9pRHj
cik+2yDkl5XmndFAEFbGKGo/VpQOQEqafa54Q3RVkjxhhLiVSSESL32vdMhBSqTE
2vyEyyNlVWSUfln3PDKle0fSSzqzqPavj/4G1rleMRoSwrbaGbv7PUPP1KFrmV64
BMCOGalrnu5r2uZTJxNpY8f7koFRAlHb0NbtaPAhRMz4yufqf0nA4EYDFLVRG8FX
yHrBbdSJ5OGSA6HimqjNEFif775u74TNdUr0NKwm6B/FcteMJFRmFvA4HpZJXZ4a
+YKW2uGbEXK4efGdTwsoPqfOzM+wEidhIVV2LC5Tt0BXHuU9oThug3saGbryxiNu
zqolUuxZixNJYgkCP5gtWsNznoUbVvHyVhR+V96h7Oq1JutT4h7QQmejVfA+Bl5i
BfPrQfPB3cR2YYUHs5xRBxmOzWgtusg7XJE+C0x75625EAao5ds4c0vlRv00dwYZ
QSHtC0Lm2SWmKsjiD+PGFDHEWPg1RKyWk+/3zqvkmiOlpqZxkUDk2zjJbBNy9gzt
iHWaWpcQxhqKMSe9RMWpNu3N4pM0ceku73Wi9hC1Fa5tMgYpWQCTqTnWis//FTfx
Kmrijs3GCDmj9sP+jFju3k9RjNEzbeERuP7a48ERPhgJj4NlGug7qGB2k1WWIn9P
a2qjYqzG8vch5xaDfn6MiC3e5qja39vPsTGwkhSy84dJ7ohIj4/JXaidLSIDGE90
cDGUwEQrNlp9flq+mDhCEwUSEuhDChvIEi4JRU1qFzHrS/DL5rh34yAFRKVdxzDU
WhH8GKnFW6s+fqxs8kko/XtyGxRuvQN9Cq1sLlqxFKZVo+KDJSAEO1BYWT/L48sv
vAhjmr0aP75gI+3pc8LDRr0cl2IJFvRseR9gG093QlrzTfPEOb51WweUhEfx5qYK
9snmN/7pz9gt3U/5zqC6PgVrYLYJMhPzJIiT49jGx5kj9wmzafRyLPo2DyQhSutR
CTTkmb9XoDcuacSLjtCcq0ODSvI7OpFncR6bLYMO32B/9c+VfYG4CdGRiNt/vAyX
wTkBrLH5fhJDRJCbd+UGTX0k1RhPOD9IzY74mmaw5hgiId1nHd3b/fc/+A3gsKHp
fF/8ffujszGl4Jqua+MbX41znH0itsZO46PDRx2YhB8tAy/hAlf72qeViYo2kS/l
664tnMt1n0aNqUEVA0nBIhUMA77brh3CMXuPdyZ/fOKBwqn/Vx87FCfuTBbZ7Iy3
9xrBurseubURtJ86NNkQuUv9EYhMdASDOBYgXZScK2hFDgqpTptVTg1Opay8F/hP
7MP/peC6cLx24XFxep7xLRr7/IG4U9PPY1c/Zny0xsC2NlYJ+ySNiqpx+2IxiyyC
1vvk3+lUnfmZTAumoLDlznfrQa5ap0R2YLEuzhK9ttYag41i6NxyIYRQw+GDCrPe
LsSXJG9KE//E27k50/PGosstwR13Ylx2fzQ2WJ52uPqw2GGWs3bOzfpQ3LYHHgxD
0ONnhYdyRzHS8trWm3cTnFL2bkAJ90Nij6kTSp4ifXP7kiUcWFrv/d8fipEgTFXP
sHqCBgDYj7JfVwKdG/67zsP4BAArWtOcHuC32XnYq5BSRPq8KT7VIxuKpusOWOaB
n/Ry+mKuEPtDKMaz0PpCfR74YiyGFx2At5yTnAnaL5zPa5rvRRx/sfjwFcuxvPs1
tleDfkPc+WjVMoVLuZwjuJNAx+HCVr/fbbYdJ7qyDKFGwmXVE1lntkH7efztnTnU
rxZHuKPlAnKnmA1V5fIw7sE324qbCciyFCxOtsLSy7xONVFmnhAHm1Vq1SMl8dmX
fRozBYPWeioBHHWZ+MAhd1GlX5VFraKBHXuhuGiE/D/a8HXSiGOng7Y+oyM1B8mu
J1ruHrdnRJM12GTMOMNRLDzk8MU0oUII0Ps81jb7oBAkSeeWz4RksEB6Piq+SztD
ACOMgUtyAubfaLOsrIoTjcbc4rvl58POUZRY4V0qx8+djK0hOL7E4g4U6ojk12XT
Ry/HVga3jS7tKouAo77n9keytXRlrVaEiXFgneSWTla9RBESoc5eVKOOgxst4hza
+0bG4e5TO2oRnS/skcav0shGy8VHlnWR9P4Bu/8la2SOXHS30V5F+JZTl8nCzLFX
zvyRbyDVjfCKpsg0ftn4gKHVGQZlDgsAoIv9MqDePDQO/yudhFVeNtx0mTGDgMo3
4dd7+rtqPyfE086w+KIq6Uk/5g+ZBMsXn0bEUBMoMaXPEsePEy0TsCvCAPtOsrTW
Xk5MNCr2/nm+96iTWUxgPwjBkXKX0Ako/KSPh5yze6UXsRqoLKIg+2zZiFR2xCjc
uGN8I0V78K5kxJQc0T+VNTX+YgJ1yRIQR93yfeKAHteQLCo2O3GZQrxAxLHv44/i
/9EEwT7pCSLJyMX9naeW0yXulyUDynZyxitHSn86a8O6FrzbqnS27XytOx7LPD57
m5kTtkOdvgYP7caxA2sKCni/A1KRtcCcin2iy48iSp/FTq0Y9YdB9757TbQe+ueB
tp4vYK4CNeIo9EfVghbL52UgbcFP5IlL9NE7RMSJK/ViAsaTVxASPek+1zYnOx8Y
9y/x6+c4busvK+bkYBcW3B1pbzV64iGLhcTGukoW0ShTaIoQAhmI0gsjgjjYFgjv
FTM39seTgEXPhfzJm1wfxrAPcu6/aZV0Ky3UAJ9et+cMKYQ+97oI0gbIL168KjjG
RpU5W5o6YVBe9KOmrhZwXv/iEv6epXRoymic21PfDo9lyOWYynUXdgO7Cbas3TJh
6U8cjNm2p4g8RHbTLFHuVXBSzRW4ah89qvei0z08i/OA8qCLPTwEsh9ezOMI+FkY
qH1HRnNG+hv0PZabuvb4kb6/F72TlZJRA2BJ86DX2Gn255tk3iW/7K34T9RAyDpa
Pk+dcheLaFWJwPlX24nublPewV6S2S48W/nNLhdhxd04cU/FBo8Gl1x5UptfbiXh
N/44Zu0ohOs+2yGKTRHWx11Mj760dVGzyPfBB4zvWDJsbj8dBbm+Tuxr/vs+61ng
gnqyaEH+dNdtn1eNFTYQ0DoTPoMjhPb15TtPspblTZiyPCYwN5cpNpPNgoDw51Pl
CszVmIQN/NSHkXbJFlt46UeXaYSwe2rfC2FOIcKVXc2pW/TRbtHz3BZwVjfkQpe5
q2NsHLU9+lvlNW2f4UxDCQlsemOjmvZPFpD95WldGzEcrBL5Zw6mNFJLAFWnFMgz
kRJOjS0rsppYDvf1Ke7cz9MafreJc3VNNZ+o2hi1W+nUNAKCwyzXQnowvm6DWMQz
2ogZafB4OyPQSNgLWxM7iWAOy2ILov2iZEHizNZNA5nPZr4112r0F8ym6uVNeSWa
YJR4UnQUzI3w0+4ArdwrR5+p4kxtZrnMfp7/ZX57DR4ocT8+NleOF/ruh79pPKpl
Pa630xevJTZU/MWxwV65weBCWBHWHCuWw93H3vMV51yBm3Hd6LRNurAL0Wv/1Y1s
Rmxs9PjWuc9saDrlEtbtEr2q2K4tO0CtrRXYhtKmNfbhoX5nt/ssi5EjRNkwOcDo
cdwD71Eudus8zoA7eCHg1n2dRtcrvZGNXactgd5WPHOZaVb6vYFWwJFgyDEka84i
ub8jjLSQIn4Jx9Ty9BKXp9BCe5g7TiQ145jP9QSU4xNQuw7hB4N4p5U6c6BMBK8Y
w8kg43DE0wHIatf7Qpt6ggbmlHHpqf7zuU6nmo0ZBdjtecJReiQAvODTFHrQvMv+
KO2ds6RS7XKha+zuDpCdROmuPlZWA7kJPL0cqnY5kRt9nfN2TlOn2iRt+qYClNJT
xoN9NTWs7d8TiGqQa1ya4PSp9QdUga64J2wUkx/q/3rcD1upO6R8onEEbU/NKXn0
y2vKy6ERy8ScX5jPHNqP9UAyi8UUmgQyi6wsaomP56cagb0Zuc8KPnlnJrriwIDe
ZLFWcFNjrY+IKm60vdXHuexDXJfQvZlXmYIf5dhLs+mzfMLBj6cGMcJx06rhq3ft
HN5JFPJRPmLCpYVF8qh1tfZ9rgg04cBSc35k16EUWjpqm//xlPTO+GFDvhZDpgTf
eRXYZ+v7OCFkKEhxmXchCTFvYLP3YVC1J6rwMYacuQSWwyIIXLP+pzM0AqFK4yZE
dJrhWBYQJTQ6Y8CaOK183btNgcXIh0/2lzw3X5uLCsvFT2MUhTWIR6CWb2GHgttZ
Q7aE7RxNcodE19icnwAlFkwIf1SYjjMOnGZQZ87to5WlaeX054MC+9lkTYPupO7e
9RnG7UJCj983N0CLZI4CEB4XsEPJbliek8ve7zJs8uBxZlfYEAa7mbKfmi5pXPwH
zlRVs4LT9yJObpGMY48JVg5i3wISrrnFV3+XxCEKBkCosJuRWlWc5HpF5LKkWDuu
H7z0f2v9A96FfznP0Au88Q7DFX37EUtGnUKjWqfnBSWGae/GvmubIocKRVWYMLq5
5DZeiuieQA8f2PTbmrWtu5ZIGjHKAy/vJzHbZDaq/X1b4ZmOxbEkujc0pQXU0JEA
Om6GLrOQwjF50qN/I8UgNKptmdZCn91oMWeIAm6eekKYzt7L2uOKl+b8ds2F+b6r
9azQ8v9ZLUe7DZuBCI3DiPbYhsHePh7I6T6qCfLQvyulLNINU7+qWSR+WBlvvR96
PbtjYMOxo7QACE4IAlOoU5RFhye/xqF+mDbIPaE8Lu4q7fbp7+wVv6qTjovXW544
StCoWoVx80UR63Hx/yWafE6J5LBASj82icCApt45edvtBrx2oA0nuSkWA0+ejmxU
+r3VejrWZue48KQmDMBVruFZnubx2/EvCG5mP4LeD/rTycrWbg7O6lr0qL37tOFD
3JP7MQpyJy9SNeoJoAdxRnnH5//TNsul29Lq32Fq3Tor5/yUAHz5flD4NkmbrXjS
myxu65KB4CsGerLVUv8Nkver3wgeIGs0N3TtkJ9WSfue2b1hD46RE0OjREp5kDYP
GYXTWd1PvJ1gnNo7sPRks6zghbOxtmATs5HAtyXg52cdi3LQEYsArBMQ6eTbLgN4
iYJo9DjLp4jnedtHBseGllE0NAv4m/pRUqkqedf2SCwwoYY2IjZd5ZIaN+jZWGIB
xWcsYqW30IRNgKbbaWinxsqWjxdub2ZIVe805pb7WSFqYh0JWKec66ilLv/rorIY
BxHhNjMQx9DBYkJSm5gdDRTvjp9J+qovrWURyUalWs2v65tEvoLMNSDEgE7pyefV
kdG7X9vFWkx3vylOFz5j4d10AwovCBCplFaEdTtqi/Lik+swZUu2WQO7bMtCeHgS
ZsenDeqytH84U2iTioIwgP9tfe5gWrZ6k2ckOg/HrKXd4hgCbeBN8sbOB77l+8Ja
Va/aaKHJgSUPz1M0cnUhzhw91BLp74T4TnUNl/eDs9imWNyg/bhHelivK1zkL929
K+8lhn0XbIQm3gaU+gTU4gzTjizhl+LxXncVZYHl4JV4OVPFceG/azX7PM2vCTqq
SqMyj6GlS1jbt6O6zhb+ImL93TDL1GMELkcgox/2C6CYThzdBDqtkTZgG57zAulr
c9VRUySeS7I1QDO9f5PyK+2ne45SYYOJF8pWglbyOYpwSBGgTHSaj+beBd2RVYR2
GUY1mSEZXRXwJr5NPalbtDCrjhIg/PdHOEBM+9nNuBkqJeGj42YCnkRfy+u0/Gpe
q7yhPBVv36r7inOmunf0AwNcSIDKBt3e+uwKq8YKYQYVxbScp6RgoY8/EgCLPW/f
vXZFiWpSwKVLGzBzL06aouIGtIzwhl51A+7yWm+8hFvB0iMoDNfDSg+GGRsa/cUd
DbAFR3U1LbIFLF1xxNsudQ+RxH4iYgicM36hLL/x2aQHdPBxKDBVM3ZOJ9LEsXD3
urs/xPmwOG2vanf8Sv2sGIFfz7/FwFkL29HShoikYtvg/tC/6XKhF/eCp+iiVlIV
UpPMPK7qQn0T9e6KScn+nDRQe3fSLzuQWy+zBFYsDi/560hNd3fUK8dOPxwT1o9L
pUb+OPSIreS5JWQsZ0cgGJHZ8I814a/CIgDlzv2cRrzpIVlS6cpv018Hj08gsr2+
VNSFcIMQTxECF5+M+aw9InGv+rTSundbT373wwjPJPsaakDBHaV/kkilth+oeEti
MPPMXEZKYiAW4IV6nn3bk2GjrgjfaJrMPY9rI4YtIaiijiXcanjKp5MMsQh4juf8
Ao6XF1Vu3fWRQWHF7UssUnd70uh2CcbHyxetgwXAl4xkQKqI+eBohW/xM35on3jb
MpQE6O60hrKjtrPMuA3A9NWsrWDi2Qe6m2M1P3qI51XazlXiBWQgNnahzaVSj5T8
/xdNptxAh6j/YjKXDDiXKtfhbkPFMvQWv6w2mca5tnk4wz67MnSuLFhMY5nI2lmZ
pDQPcfJuH+5eSTK3nZGIpL9/SJFMo6Z6+GFawsnUG3egd6de2OUv7xu/G/2R5XKx
wTFo3+gEjqrMvyOfumXiPM5Fa5OPc3JaSnnPSKem2L67NIOvgCPXOXGBNI6wSOj+
O6KQhk+YiM304P/1iVmc1zErrqZkGIPQSaZDYitOYS7M5cCbRss0viGIG/YbCpJA
H96hDNCovK0aJrxwVLyszctfo3WH/Azwm3DgRfrgZpBrL0jdyavLvw9uswN6DtCI
eoVLTPUuBk5VqB5Uj1yHXHQEyYPeawfBi5SdwypQHODGAJFVcxlnvJnlQhuPOG/L
ZKX+mdQMsP38pDN4UGqCaXuw4Mr4ITIXUVYwGkzhUrPlLAHIzBaHedR3Ozv6ytY/
rByX3XAv92Pzuu6/H91rERZ6wb4SVF1iIP7ETpKiNX9xHobpW6BF2CCHutLg8ZEH
2/1TmVcAlSIJ7uI7hv+kdE9DPyXQc+PD+SPF+Cgh/ZfDTJfpRvNx4Elw3AEsN9OS
gOefw9u1cMj1Z9s7JZczCMhK0/913DVKRy+YqQ2UsYOr6MuoUwM3kC6/9QuZ0tWg
IqNKbBj+G1yMVJ5ma2HDHHrMG5yb8uF+7FQEcUTcpC2EmieqJeTktNlGdAS7pYvy
WeND7ySEoijhKCTe3HF+CRk++WWfoO6EtDzMsGHEFAJYPP4blA2AHh0DhqKrRDOZ
vhc7s3b24ZmQMKrQAMcsYcqyRhyEUDV4NKIXpF+SzUmN7hZMRuHCoasY0eKJzzlf
JAyE3PlVyvbGVAJYfQE4C8ICyJH9k6GLXIT7LJm6EJWNgTV6GMC6orGiNOb0jzDT
hwzhi7aUFva8KDA/RtViv17baYuWEcNRqTUjrRA+xXb7iVcmHRJK+mZG92zngoBA
GZbF78j2ui6uC7ZRYcxZSbiz5X7JijK1eaevWBra6CseR8rlDPa5wuE+4GISoLjH
+dVTlRG7upgc+41Hup/G25U6wWGVgqjQg267+OY0wBpi+/qwoR2jgi8ycEvCPJgQ
TXJI29mjqK6EnRVstR5SLBkwh1LgwL9NsvwqR0kFLhDnM0D9RHfYGfNjzGeJhxya
6/QHIsiJjdLMfpOZu9x/iPF3zw/p5LCefnb2RRSLaC+SVvhIQlyYjAnWqn4Q0C6v
oDjPYfG48lEfJt4FblKN7raUNXdAgBoXU0KSq8Z5RoZxZx1bdCzji45xrInQR81U
UHI8bsvVrpD2yFiaO/t1f0LF1SizbWBgo4ln7+QDZNaTH74l8s7sJjkZ0kF83JVz
8bR+eEqZtY0ipiziV7GCrrCu6594t0HbYwDS9ee79RzQXwCdUQjVoPjU0t3NC+xI
YhHkmjQUr8+VLmWTCdCllhuoGkjZhOBf6XClL1au8FBwTmkV1XwvbbDeWCNeUf1Z
Sy9gqaZUmRk0n16FuwNvICUoLH6dmeeK4VKWhWT5+IdL/4kv+Zdg1dZm4qJtELGR
1tmH80sGtuonxx6X7ZOOsf1WLyKUG2NvRESvxwEt1c29YDB92YzhnF7R0f5vDycy
q/iKRVjxS77Rc8Duh4gee+EGCs7+fUlVwstj/nxzoYBHzn97KahURqHAM81jnQ9c
l8rS+Z07toX8+A0oVoWnGXTzq/kF1ElhcHlXStMQ3dDFTtSnyjQV2plCWMyq1BCe
POrAzJIX0cIbQFvVDn4fY52sYqC07kPDQFbvUznz24HOuuf2SyWkPfSTqZSOx0EN
FJZ2ZZtrKEQW6joHvfADchG5hUjcLu24wTG84hWAy37GBp0a5nOBrsaSAwiUc0lx
MYmgRGX+2T5YYM/O5HGgRYksmHPCr68v3YIdRfMj7171smiVdkO3pTmT2lb4c6KN
VUQV/umYDlB9Y+iaapuuul6o/ohZhbIpCr7WfGJTmqUt92jGxdUVuPbs2A3kML5w
ncKixn59f6FbIxnDKo1Oge8GoF113FdKBAq3bvZ5YhFtQJYQZdfDIpdkTUFCXrCU
Wc4WPcTl0gqUvsWxB9jkUJZ9qStMvJKvGVmjtFfw++qbf3ejtHcopezrJqgMjupG
b4/xk/gOBqfJD3UE3y+Vr2gWABZEApkc7JGcnqCiNAtoGqUPgj1j4GNa6215yee1
AmTtV+K7bvV9LmkqtN10/llclUgWu396WbjfGVqbS1z+1ey63lUPfyT0VqzteXRk
TmZLj/hskIhYUAi4Szj5D5qEZiCPkawwIWXHaGPHGRkcTO4T6hdWQvHyNHgOvxum
6cs3QYrNpAxwuPuUVTyi1M9VI3EOInVBYPj2Qjod/hTbMYFS+OAIcNwpJxKlmLas
rTrVjXdjX+Vhmbc2Z08VoitSkorgIlDhAyIbnMt37oWv/hBLLSvKwMOyD6Z3f7XR
dW4jGY5P2+S1urGl9rqj9V/CWnl3+BOrW+Soa/XeKDossdmMyHi/xy+UzbmlIxmD
GYZG6kgMAAMBRAiyTrE0vHIFaAvFsECkVBfN6gOX+szgtmsAzSKiyJK+rrH6jfPd
4RN5tlDIjz+hJqr8pJBfX+6j9IF7HytE2sVWLShYANOeyyaw82zOtOL2jbsI1D1L
Flc+OWr/CSuU1caNOyo6CDH4jn2+8iPEbg4FJPoS8x/1SaDyP/ai38iFoa2Pj5Tg
DMjndOP/GnQYD3R3sldH9BareQCOmq6zpcyFtTDX/ZZyAHKzawnGu3ZunSizxJAZ
W2xwncMgQrSzze/7ZnImJfkAQgQphVY8lW6ZRIBxPoMkYUb5EEhq7fGPS/lWO5lt
VcZ+CPNXmzTllvH+yRats17Ziygo7ImFZDKQ5TmjohbiQMWnfdZv+vCTfYCvpcgQ
YlG72YopZGXlWayMh/8Rkbcm07UJs4qyMf+m/D0FLfKXASyg0LHKlHGsHAeUk6MR
DzUOXrDgmWuDRSJpnhFEXRWWYo475k3v9cD4vNeOMfazLxc4o3otRIwkneKMCSTR
/vPp5RS9f0guq0xWBRQ5b6DTQC7ahUsl2FiGJ1ZPc+svc8vlknMRamvVj/y7+hBz
ZtBRROlbLGCzMn0MQD/+jJQAx10z7GNvL6483rpRzpyLUDpOSvLroSbAok07b9wH
FZV7xzzEPtwcOnd6s2ynpF+xR5y+aVUWKNkqs9zuSuGoAoNuv86mi1utOxHW5YyL
dS0+BhgB/GTqy7QRK9M88rmiogFS2eaa2qMcPpcMNxAdmp22tbR7qzCbZfr6S0Wa
jkNo0MymHCrfkMQT5HeO380/kfupjYnkRhJtFwHe9u4tEbCviULgkCjnrKzzyxk2
V+TlWy8LL3NS+T1ZkXpRVOheAEZVa11dIBXJrkIIfi/GwR4NJzrZtHS9ekHcYF2H
eB6zEMkSgSBuIlAjoIznq9vdAxm36Z/pwYhRwwt0NYe7LhaItlxEtlSRGSGFZAP5
BM7POJ4z6bOmZJl84OA2t+wJ4gzQuAPe7XAAB/Ao2RROqVXbJdkV2jmALtfjrCcD
lWUUd1ETw+jWfQwXzyt2qSjr9EUTr1QjkbDtT7l9IVmgt+iU7vJxk62HqNl49Pge
S+A5JD61sHaBj30OyHOYwmXTWBmrAbhENm5CkGeYMlS6JY9pPxV9a50sarIIRcG2
q/aViBqwlJhCNvqqEgR7NUddTvKyEtcELjjVrG7R7U6+fQ+Zs/oO89pruBx3U6jV
jxcO+GQwdNBR+zqeSkLHv7hOcP3c13Cvae0zk0QJ7HgSTRRYJhu8d0jxv82qgdf2
fXtClYs/wsd9ojsuhtVaTWGZWSh8YkOCjusfM52X4EHQAbmg9f1KO2mIsjTTSj1l
6Ynf3GC1Aziled0Y6zD0R32vqSjsPg3O/GTdYKrZP3sYYcu7z/G3/X1Uzzuw1sNv
Fw7qAikXR67aml0gXa9GdQwe+YT4QWGZhSlqf5neP2FFqLAnPKzTjmILC10miJWW
Klghqrn7m9syF8y2YLksW16N4kEPH6rJetyLALW3DPI39xlxkFFEb3YqjHdRmyHM
byl6WcmSdYUhbPYblKLhr+1dnbkKJjqecZektfi8n9QUrtuAVwQln5KeMMwBIk4E
h6L5aE0qBTLsgnmTgvzMxYimRkZTm6AYHsTRLQDOVOrYMWfpzrwD79yka//VbF8e
jj0TnyAmGi3gSAc5SwcsJ9+J81SlTCoIVlIILbzFSuxJdKolTzxXaOGKba9O7TzE
dpqGD3iNHa3makivRvXzxIY5eYIH/PuraVD0vvq3YNfC5Ggln1gqv5frSN77iEFl
C09nmdZlamV5kZgJKS2usVDCLY/WwjUXtg2liaM2LmHdjSQ+BbCyd25EKyzUMcpP
SBGCQ08lOfgeB4TiFq42fc5+OgsU2VCMThkwl7xT02fNlejBzy3A/JW/LeR2/bZ6
WXwsyxykQiAM3udWxyrHW+CnUR0B1riv+UzPTJnt5iMg+kUUbh6BGCcuXbGunQ2l
cV9zDBw+M9hTkSovZY7kzHihW8JsVh+tgK7jmHPMrf8mSGm5Ae9R8S9zkWg9q2ev
i1r8ed8lp80LFgb2QVJSCHXPOVppBvZR0LBsTGTbDt2YbZFEDOes9e0l2s3BJvBk
IdQEqn4bpEuc0oqnl970QfcnrwF/KjNW87xrBDPJin10UpK4RwyFhT+MchK4UwWs
0kN7VjgKOBBbj6Pp07dxQHwb2+NqQhbmRPKPGu5SDF7BLPzuyFUo65IehCz9FwDB
SPyl/x7WGAj1cXk3l53XZaPYF8h0oJxI8wp5nY3Uentl79vxmcPh/BtrKBtKjRUo
Lkkzx3NOxBrUa2u2pxSILoE1q5bfa4A1B87uRAcom4sSxmGZtcc3GOyHYYLkho4U
kAr8jA8keTzgHYapegdnNSGDgQhQTDeX0lXu+tFr6GQf4f0RQ9Ogc+c4WpDfBdti
38TbBR8I3pV3Xmz6P9i0Ho1hh26IQ+8doW88UHJIu5ldg29OsGEe5k+Y6bagwhCL
cLPybeW7RdacIMZOU3JrzipcUPzd9b1l/N2CgLCmLZQVxMDwe/JFe1ASRzTiPXtO
90v/YZZOHTgxcz0pmmbJlWO3AP8zJsyvL00wkNjzYizUNkFWfqREiiBGLrIkVCVL
5cS2MXaLcTXK55NBR9SVEDcQRNV2FcUIk+gIJwnvaAtlB+Y0Bg8qcvN07RQKmXni
pXO+A4SMQlqk8cyEnXAMjqQThESsH7sZpMTdJhJTNPxWYpQQskw5ZMY5Rrq02PdC
q32SJwVXOIllWnlbcZvNfLRa9RCR7HtZLNnsxpUxs7WxjOa+oYX2XCT2C3dVjgHL
CYWzP3huz72tRfMqqtx1Wr47S1FWL7Zw/wt0kZJoYsMNpRutrRJavKNP8JW5t5wp
1QoQtB3YfDVfB+YMpUpRb/UGhuDXZ2gTKWy3CF53GWbgtFgdrXxVp6Sj4h9r3uKO
chvVEW2oDPfh14JWBOK0bdIf9LZgcPoCt0ehsEeEl9BpM3tOC7amkFiFYge35GVQ
v13PMpCDgApqm4FwkW4uGoB/Prpg2lHx86laHwoooekxxbftj9UK7zZGLCVAhxXX
RK94JNss86ZLI00wyBe1zk84eQ9/CSQU08+Wf+tw4E/aeiqLcyIaGiyLJhcAiIFk
E8rc7tnzXT0Y6JfZi9kJ/+FtX7gKD/XPg2sOWIZ83tVTyuOyJz21stZ5KkBUrZt+
KBJIsI3japItgUY336uP8gnt9kVcsMxzM3H9pHp6IucET8fieyJJvSKfz+V/tAm9
9QikZtuc/q0pmQGL/RVRbWXNOo02/3sNq9P1FOlGDYefqdXosYL/tZr5rHfvjvBc
W3tL2bSUnoP32K+xt/Cax+Q/Bf9v24RbL3XfkpRy1g3D80GbE4HiGnEAT9Q0OdPU
CVk26Bs0573wW5U1b6nP+80QwRyeLyQMCydwKaSm0FFnAL1BW2+973axnUWPdkgk
jVpRsm95XZdSU5dunNijqjuW+kDUDlN0XSi84n581Te0IYU8W0MfJTosJNBoc0L8
YkABdl1E5Y6Ysp07l9eJYCXDrMGB5sIW2GcCegeI/uQ8ErDfzGwY0qIktOCgEFcr
iY12nYn8Zyjof2u2NbwOZ9iomi3+DbREsGTvl8Ng8s6/EZIXr6jgWTXLQ2FDcn0m
cLxA8GhDlSKv+8Eq1sk/wRcKhamlHMcjgBQPlTtI2RA0VS7WTT/YNP6lXSgA7TVo
dugwb7gD5t0TN1G22ZgfUHDQissV8F/usytgCmLxQKOJbeX44W1RwXU0AZo5HTFA
qS7+/KWfjguAIPo3G8g2ffGLQz4aRGzrN1hcvulXaDMV8NOEuWxdJNnEhtDAJEGr
6AbGkRWCmWOmVYFXpBZHSHOKZ/JZ0H3or3jgeMg6MnCB9cGjMxkaUR10PFgeuPWO
HHpfEeE2etbp7tM5r9D+7d90ObNwg+RD17nT85Okwjp6eHB7JOwRA19Bsutfjhvh
EVQud0HC8tTR5i4KSart4+RrTdsT9m15niAGe9da+Xo3w+pBErOjBJqHYopRaY7Z
rKf5iuDh2QRMON9NLP6osRC8Cu2FCji2JkUAmZ2R/XTnbcQ6Sr4mSLqY3/83uSxq
nZyi95vPlomPdDpE0TDpac++FeuURMhNiCCBvcDbHEfxmSD8pRK++skz7ugs/b+V
b0+ZDFflQKci8QN++NVIfhyWM26c4FjGdMVqDm+sFT3ankoz7oHmA/4WoMhagZzo
YBRhqToX9URpjXTY0hhyxxGZ1t1b3Tb87l+pQbUGG7FZWH2fIQvKlBkBt4+xebyO
m/VwcUVXdhEs9pvLZ85l3UjsxC8CYMJdoh0TFhaebuLJaweVXlRV3Qf4yyKP8O9g
5iLHPA/2+dgUhCWvjza9ZJYT8DB7pnMsofLi3Uq8qVqaIt5eHcNYlPgZqh49u4Ev
NqzMy1Ocd2PJ2F8hwHDX+XVTUXzNmhxUYkliZ6CTW5I3IGTmIboHCJ3wj8J1rgb/
hjs9BDNNameyCn90REdnzlNffLSqaDfqmbbhLU8F/Zo2jqrPKL6rJLjZ1Bv207Vq
crHEbvxTF/4kStofVB+Adn+jKpxRNabp+Uh0gyHcXAZP18Zd6WniYB6rEQtuAeLt
JO/b8iJwbypkJMtLrD1zFEPzA8S08uMbXADMZ1pPV4Hrwb/HzpMOGW1+FIK1FG91
JbxPo7+/4hLDWKTIzbUAD53FVBCFC/TX8ww/y9QUrbUnYLDr9Msu1OJ+mn1Fi2CY
02ylsB8MYDovavtARQ6gtwqtH95FoT72czKMEjcYBZw7QxtJM5PFnEcyWo4fOG4w
m0DQ3FG7kbGbcRAp8Z73NeAzTYmJyCj3nxTqI71E/mcnfyQcTylEFpgZcRMAg4wx
1n4CiVxCT2RbOqnsEulDVtoVzs+43o/OAMzQ1E/D7heKyk1oFPwgBc6340GyhF30
k8/23jGWwh+6iEFxqsGZ2tmw+Iy1F5B1znjCbt7zpn2gWBP3OurizEraYNln4XCe
6kZ7+mdhRi+ZI6vy0S+GPE0/SdbjmH2ICb3Tp3aQ8lSNjyhOMvi8LMVaIvk0/CMa
wpfDxc+LAupWWB4kONkoGU5CGPLsdveeidrVrRuO/eXHMZFuBtFAY36AFNWx7ob4
H52GjTDQ/Ovb1Lr7xG6tPgyI18PJxxwmxjyx6UnA2jd59Qu9VYTfephqvv8kkoIy
akXz3CWvtloglu0BZ8JkPh3PFXIAjb28jy53hY85SvTkqW/FC8KNQS+DzJXNdFO9
2Ku0R+/tQhHtUUhe7aq52+K1JPGz4YoQOjop/5DO7+BB7s6RZrN+WFZCfu6lQEt1
LEvPRzrFu2XtnKrQW8s8heaB/rMwVnNOpV7qXllMl6gj8mDbAw74cB0WvQco7pK+
bKngGbBUTFaLCjDYYPeoCAjWIU7J8+dKeeO39g0oUKc3A9WawQoK2s0XP3EPwDDa
9/n9okG6MLvW28tulaQdk8k5UOF6aDxgKXPFf4sNH2tmp/7l6W7q3P7kjqgjBCeu
t3WHfHozV4bY3oUYpjEillBcoG+EPVf4OOAOX4f7UZDWKUZZR+HgmZBWcooUGi35
90o5D3oB1ZjmBja4Lm9W1c4QVPO9qufdizTAwaOAgBjobkjPUxUyTi9SGG6ReKgA
duZz8oV/5EJOAm+YzQwHnLlUioSS6ZOQ+VgEjbCn8Vn0rwx0NCnr1PCjitGu8npe
EuDb5h8Z7XfUfb8zoi0hROlWWwJpXiU5P93h1y8OA5jP1hfLaGNmK1o8zYEJowF0
txfe5UBu8CMjYcR/0FrocUA3qGCXksAAWZWDfIMbuN56FW4jeowaMxmJN2I4hboE
e70V7QQZxZmsYIak8V8UuLl3HFX6kT5EFJUemBwVCa8VyKJoEA1zMJ0ToB3AlbFG
rcR/n/9Ld8KQ9n6zu2cz+/1jOGglDaeExs03n2/HOgzFCmZ2UPsGj1Wn/cjpP1PP
nft6F2PsaBNQz5nTBaskwmMm4BV8CU1Gra36bArBZaQMOPY2olSwMe56M6SFCfhq
Pxsdb2dxNEFWsyfZrTKMUJDO4uS+bbCxPO38LI8tqQa/rFD1V2VaiIt5Sx6Qsv2J
c5dhWlMheIl1ZoW4vlc6rJYNsu9r8BfRdoMWCn9pCbmhtM24D28s6hL7ZR0gel6t
/fS91c7N1yLJvKymwIwJ6XqOcytmh/EEYXwB/UyCx1bkvz+NZP7SBPrancoHLuaN
nF2eugAqMjZAeCXF720yOy51pjr2OxjcMnsXK9FHsW/KvFyXSZLvf2bKA/cx5lNc
pbiYmuzU0kAd2OQ1X4zdI8aHhLWkYORlJXM6qsiqeugzeu0+RG4YprXfzD5tLQZC
/LdivLNkq15vX4oKIEx5qKE68zMJW73X6QwHDHGr+mPT0D1XFsnXvgKwI4+H3Cgp
pyyT4zXjxvc6fsmZqmLKtIIHAS/iKkCo7C2m6nNgdCfrdaxmug1t71xNP95eV0bB
qv4KCKlTDWytgNdYdS3j8mXnilD7hpqqsczn3ZGEEu8uICNqRkgkwnnRuwGzVTO9
mZJZ/IQAp9cR3z+g5Xb8tgYcT1gZ/gAh7lPu8Vgtc9nixqmQJS/RuqCX1XpFDUgh
R1fahnA4EnbOBRu3eMGtgZ26Evl/D1pIwS8meUEdx6NquV9urB5Wh+mI8S4t+iXY
Vg45OoJsCFZZmt74IYMMgS5ElLtXPAyZk0l7FpXdeTgDgvP+zXSOEILrgF3K483d
bID5X80Q6nV1a4y0DPIfdEIFdZW/Oj/B+hZq0NhNINbdla0WbM+06NEEmURFhJAn
ERdl8uKvLuRT0v331+9PZItCHrtLEpVUV0zNuoKsnPd1GuqPddaQY9r2dhEmFksT
7lGF/LKTb7rNm7v4wUeb+lfYvMV3/kEkyLQrlAV+Q5xctf68SbktaTuEQCAZ/Ac2
SYYcd0LHIDKiPRkZbgWrWIZu9jINVmslmxAnU1Gq0nPqaKkfkoPO7++be6ZW9i0l
ng/3dOkLxiM4v6jUAOJT0gN/YvANfApv11eYHjL/2CT2JKlLdvVczmkt60QhvREW
9dderVpkSV91kW8RXndoI47WbncNxAheSvFrED5LA6XhYtYHpV6zvGsBZVV6rkm8
vKFUqxrgNu1SC3xA8UikDnEq3x8qYA02RmpoRGWeanqhRyfiz5xD/DkAO5UaSpyh
1CEXBcL5DfUxoYE5qm2sJLdHdzxKw24MJbBOvnyR8VdIRxDDNCZErdgCPBOMQm2P
0nwKQ2qk7VRVdHLBBXWAYLZKmPuN6SrF3h+dooalaDsmayIhAFuoeSfIp4t8GYbX
iYEBsYkbR8Q4FQzmqHkEbnxnhqKA8kIWbamY3EfJW2e9X6hVtsVqv2d74oxDQDSi
jRSuWYfecDc/56juHHUUNhBVKHwbpgsCC/RvCP74T5IQ3j+MxD2y3TNykbpHPnMK
DzYhmsffB29UaBgHFWh/bDF6TIVElbkOEZXdoaosgiuW5SN5AOerLs6fpQSFqWzl
T9yHzxkjlJLCrY+axa8QGbHLWwYr9E94fOtVXwLfdUVVnDugH7IFOJS9v1FQKEFU
axPp0MdYR3gp5GTXjN5SCbcm8naGb55JuBmKrlWS8wDolacCRRQGISbra7Dt07Fy
a8z7DmOicuKFHsoOx1YDr5/T9pm2uDMZCxJlh3w9INFC8zs302AKDaBcA2ImU0tQ
sSdREdRtUqldCbvd9GYyya4VyOSSt/i9KSyYdcl63W7rNOxgPAF5aXFO9xG4S08O
p/zXG4sdYz9TjxekRt7/ogL0EapYcESmRrLdagjLNqS7XAYuZ99wOyE1+ib0r/4o
BEATCxi4iVaZ/a1SL5ze0XGi3YtaGbyNX79uuMZNlaxha46kXQTGzzlKql9I+Vnm
X9JwqD26aU6Kf4pfc8cRnl0Mr+QKQf9TadsIUxPL66RxxVyZh0D+nYoc/3SBWhKf
QQuhHLO7gvbYcsZWH6wPt0jYTj3QKKAWpxpG2SOnVO5ZXjvkqUVeaahBWdyF2zOk
vLmo0luBl+dsW1gH0L1NbrtfRDjgezmaNKWERA8tLIglrGcUDxga0US9BmqX0rkY
XOaHhRr/DTOzE87oy1B4yVHJ1knC8Oz+tYwbTGiRswwVOpir76a64wxjWIcfS8eV
735Ge+TxRB22URqqyPj7qkOByM1UjOegzQdBVywnm/m0RtafBgzMS71tQN9Y5akN
OWyXfU9KBz1lkKuT6kRS0wYuJFER/otRp6HvtbcWSakSIl9aZ6dvB+673/YuOVvf
0w4GeXdHKYtSRdOc3JC8JsPm98FSIxWz14Rn4qnEn1itABmrkcdqDsmAxVcj3OwH
s69FCAW5Ru7sYugJ6EULunfkXMCfkhe0ObmcRfj3o1idz4QSwSmmVXC0qZksIAv1
5bx8Mg+o/jb0Oiz/R3rSa7iV0wx2dzO0MxPgVgDbuN9FHPMszmmsAkXGx9mYtMTQ
T2vrGdJd98+E8ddaS7uzPuYNWSua0N0YIxTey28r4Td9l9u5h15QTNiDdaSs5qxn
3d5PfhHoSyuo5Ep/2zSDv6B35MCm9YtYwT7My4Qv/SX5Z8EkLsMpjiPkgqdCg4vy
28w0ZvJE3JdavSvRf2QMSzIhQDc6+mFJXyFQ0ZTUHxXqHE5MVDgUCIQ0YqedrZna
cX3n1+SKT3cH/HpwrOquut3HJMu8WwB5dlOGDEApPspZDpEz/CWczO14Pc6lqSgK
f1DEUpTAjp14Y0Q9vciw5E4VWl1BWbIe6FBwBNxU/jpVVCtThkbbpPfdwkb09T/w
Tgbf1MY2mqKFtrwayTzZgp95nQAXQyZyPj3XH2JUiqN0ZMgQp7JG1Du3005AlJRZ
QPxGAZHUmrRb7IjwSdEZYw/hMLlz1xIEnU42pOWuTrIyXNX85mwo121PJ0ccA3nv
S10tNvM8/JJfKilshqldtx5uhP64V10Z2noNMihqStEnWD59u6RO0hhOTY23oIh1
UcAdMTQdBMeYmFmFwWH5u4zmjYh9C0howC0Cj0hDnJilsDP1Iu0IzcfjgTPFz429
VzV0gCthuN9sq30mNhzEaHmMCGtdoUkU0/bvtue5UmhjjnV/0Yj3XihFuZmFUwwZ
4kuNO6v+CxGbppQYq4XSGPIjCPvfJzZLPPcMqeDvx12A9nvihSYOwRLhSkY+OQ0C
BeSoNjgc2SMKwKGSnwrZzd5H1N/g05XKkwT4zuhyO6D/OPXqj8fmmaU0tNKps9Gw
rCA511Zy8wJ8f3cuh/56pw7vGFq3s0anUDeXU6yhjr6wcgu0riOYfpkdiCAiiugr
RvB2jQPqE0osAtP65GmN35RW23ftY0aXijTEouvzu4C5NJUe/UsYjo9LgOM9BTPe
BjyIUJxF//oWsjm/hMXpCQIAGHg0YnK+ihl0U1a9+eQSHk2GRxgO7MzDQVLiOz2J
dyD6VbcA6VQCKD5IASxyOjTki3f9SZp21uOoM98RHfsS+mp6g4VuBvDo/R5P8B9D
/MzVLdYT9iUUrXPI4azv+IqaBMhWZakSRucZ6H+hhfQg1vgGQX+5E1VhG6k1beyt
BrrWSoExMmEXKPYIa5dSywTYXwqSsMmCePbEzJEBUa/qnh8NVd8kWfPo5uoMtaQw
siwYqHLMidyJBqxFjnjZjcbQh/TQks0hDHN1iOHF5J2jlaLG3TP4pinVkrI1icfS
DbkxFGM5NNtQ9t35gp/yQo5rXyELKbdjKrjns2k59Qz5XLm6osIhONlCaPrIdHUY
ieTj+3UJsMWGvYUa98lyYmTM6fito6q3z/WmJ5nxSnqvj2MgBFtUUvMR3HV19U9p
hTwSEL+g4LrqRTT1b7a/6NLlzWb5mTJdprIczV+nKWojOWPKc5UTCOlyyGBXTdyR
KZsMqgy+k+fIkbmYH6KfX0pJlGN1R4sW4kDjPiD+JESmB2sFI6m+gyTOfEnXg4ia
kFKMUx73vThD3UwuBLE9nuvdMcJD11b2zzsqkc4Zx7hVNZSzQVpQgMnZYcJlH8R3
RRUV7oYTE044bkiaYG+yEkdLzl3FcaiKEtXk8ZhHjLGFIiLh2UZ3XOqSuWZ6DihE
KmpIa0nq6P53m4GK0QnN1vMFwyJNLdkGrLxKFGpIunUd3uOihBcxDuFAh007aXEI
R2W7l30ph7qVxD5m1KU/op7yct7epihX3vY2KvYcKtvxshY70o6NRrAafGbiVwKY
ouTL9u6aA9AVSPVRvVUeTn7J8f7Z5ASdhCv2+mBDxLT+yiWP2zlUTvRvaBTynOaZ
Zb49xdmOWRYAf6hIDnZbkcbjgpz5N3H33y4HPd3Cf9RpQ+eHGUvNLhMkx+uP2wYU
v+Rn9CFtdX0QMKS82oxW6tKhWmvg1TM3PIltE3Pbgl0JpFwJ+wv836kOd+kQMQYE
SZ7q4B9rmEFtEuxWM4uyiP7dOCjqSLuuYkhS4r9Z12OzJPkV3fBBKC12hrf8Ke2H
xcgrSkvEk5iuuZfrq8/DYon557OBRJOynBm2f5NARdaKhdxsFOkzs1rl+RJUdzoB
i6pZ4aSlq/i6s6GMJm+5qMh5CgbE9ym+lgsMSp75+iU59IObv8P/iZbHo8kNPZId
aUwG5sHPxLGu4REzhv0x/Sis3vDslNC69CsBkvJqbDHOPo4KrLXpArgnDbj8AoGD
OnM9L+eXpieib7SKal36VeEqZzixwAp3lJgukoe3OCw2SuMIQwrBhXBDNxCoF/Rl
4YJwtiiuWwmNYJEkWRVQ+wuLf28VNdf+TkBB0m28enBRILvNB8fXrvFeipl3OB7Q
iQA+6JcjP8vAoDAeGJZWO9Uf+ISE0q/fA6eMyscevEYeBs9Lc2/7KilMJPBaw/Hc
5NHIRUKsHdJYYiXW2ie8bPSEnc126s8C7YMPynW5hIUP8qhV0kzL2r/hofPGWgVK
NOlyOAJX2ScejEQC0xqOMqHlagCA080y418+mJkDRlN9He4/WGr8Fwb5RWkFhDa1
n3WV+GhiQbgXm+rFTOspEDG1E3ZJydxaUSe43VSFBaIKzUHRqL61YJMPNJCzA6ZN
3lA7ventS7OzMuXgyRpqsRUXgdIodDjLU5qgqcoH0kbXKC5XRngsHcPfcZdVJWt6
/6JPLFj+HvkP8Z/2QTQWnxbp2Omjih3w51ivF+UCSYaHBIz60/Wm2oxDP8mjKuXQ
tdKh8idD1T4x25vouOLObq3PVWt/N+1FVsCZFcGFjRk19XaScUW6zM6niox06WAR
mHsHsNQ/ju/DJnYonlMN279uOP0mODyPnYB61XPtll7G2Bk5XVs5NjGA+WUhyKht
K9G9bWZMnqlb47OLBhOvGbVQ0iviDVJYbhSXMGp5yLBeICKd2T7YaxWsGrz+2yef
Kd7f4qaISU5vjlVGmQoEFKKU7B+lwruhTlkgPoRb/BnIa/3/ywLoj75qx3EFH7U0
pwIW7ZqSdJ8BI95VoM3PkBTDlOI6kAwD6Rnz0ruF0pYFs4raBPht6nHunTwWE0eF
6r97QA5hOD3N8mfkr2R5Ski9Neh9GbMJsfLH6occlb44QatgcJleC4XHjcW3JeWA
GBkc5vmbcve3IaD2o0VwHPLIM+CXN2zgbVnfOYkf6FEHddClRhWFNCtIfpX55pbR
Wmiv+gDzCM4FbA2RfJ89LZ0EZTm+Y3pwRcNsWE2qND5Wkm3gr4Gquw4HsINgFDB2
ubVTcvpOreH/7I7UIQdXOBxA4bbETKXoaMYobc/Jwa2rlupuplzFhWk/Z4sOd1Jp
IeRasAFvpE31+51cRjWVM5VSMY8QO50iF+mziLwwa16qv7HrM4CUK4XdQWuSHe6n
88AEShtMEQFz7U5B7IzFiOHj9zkaUxRrpAePbeKPktEbVGVb7ez2j08rQPe20NbF
L4JLrGl+fVAEhgNeh4W+bqyrfW4/UmPxh0exsGM8mrdrg8emtTKieC4YEwpIQGds
dPqMVA9VTFMATUTPs/0b4c48jlKzHkZsAqgxLdkGU1zQwnF1/3gMMw2jjmJzb1mx
ga9s2isrpCYXMGjqNV1BixGZkaQT+z4kY9TaGuBAiynRZ16Ms6f+p8urSP/k+2UU
3A59tYC8yhPaM4wGNW/i9PoclnZ0w8p9gdef7xFdtRZqksfF2IhM+NUTEJktVT4h
+o5rsYEFiyA7wMAytilo/1LqgCd8FhMP73qe82TE95GLBeJh+9BiKQ98webUAQtk
Zb8wCdlenc2nYXbhEiXxCCJiospHdV1KfYXzne73stt0HST78DKo2zJcCSJ/itJw
mOF/6SxqVv3WUAskV0opeFARVHw9AIXDXtqtFChUKwsye/8MericvkwqDLwq30Kp
TxfSkgQgXTJh6zF7nYG9yL2DEVq3V5aVWYcwHpLN00zePCAd03asSP0JkGic8mpD
cwY0M6WHvr3ywoVeRh1fh90G+BJgFzOg/XyPCwg18Wwc4/LxGxdHyIwxU5b8lIHm
Wj76tCRqVwplqOrqu8UOWkCs62ciXrLioFKGyvS83I+5Kz6trcW/jhK35hXAWEXK
uCsBZxY46DClB73RrEnVYvCcxvJgx5Vu/UZ1/7u9mA+6bn3pm4v4NZYCImroP6nM
r839A26fNtYc8VYCSsmaupOBJnZWRtHlhJI+lM8d3FEKsNCQEoirDp23fiGqeCXA
P21D03WtBWkG/Z/1yQ75axGgvS2YL/7ghWGfHlOHqx+5pAVdsrIPnHnAAFUPMGhL
DR+h9WZSHpYcW1/RJBRXS9SphmCk8bxRHIJrDZePMySlo3HPCP2+/hvPgWtPmsgA
AnODw7/Kye8XF3hxOy9OlyUoHy0v0MMkzpYPF7yWhObKka53Z9+591lC9kLiNrBa
VYEQGQWcfeqW7dQJ5C13vufnhYb/2hip44Z7EcsS+a5gpTC7Z25zjZJea5BlcAyV
4g0S7fKBRQL72f7z3tZ6C4J8h/yVcayALqcqNLB5PP1j2hWrwd2YVDm7bSKQPpal
FXMp0xHWOLToj8Oa/nRcVkzqzOSuI7i1e0vUQF3E7/joicFomDzUQ7sUROwAiTz7
/+pQXafuBqcFES4wv7detR7e4LDLWi8TI1mJL9HSaKEoI/jN6AY9kfiFGVRBGcx2
DuJ14VNhSlhxLhkofkbqsBR2dH5nGOS1D9+nfsMIE8RvFNTq0TwSBeMYr5e2CU56
nkD6DbZYDlKuW7mXWUK8pG+DQO7tlnHGmDFMtmSYjiTzIJ0i/gdTYDUCDEy/E6tu
ycx3ddPvtbiA+RSFeX2HLdejl9f41CXQRZQIMxxgSN9M7o5vB7rC4mqzfyfUiQjb
KaBZ/vAwUdvltbUC8+nLsvEYoSVUaUnnjxBHQ95y4EGkVIfuJrGJxvF2jxKV9Vsq
QTOGLgTqq64LmhrAf8D0uNIZfQBTDgAd/RstZyf4GGXzLaiv5PvRbql0z3ZAQ+tq
Yurn9F+A3eaIPFijnWivYtu2K5bHDbprvNuTFA/pd+zj9c3LNy4rQyGLg4W9URm3
yj8fkGi/ZeWe+ILNC7O78+L9LNzXrl/3HKfGVAAkmzHUhV3nFpmQi4KujXQyfnxz
8wq1HswrxHE+3S9zHfy8eUsg+S/ddQYedO7nC9MQEghEbFZGnrMe6UbKNIcnikuQ
vHJexFSynxIMiuP1Mb+5VjTvvWi8ACzUWVqAefP1XJqIavlAdAPMAtNeCaWGcc+a
y+G82iSphJApF48UImc3mYyl05nQcMSK8laH/9doNvHX/Wkv/RSZXySUtyMy1hS/
fm/r1nGRAxUlseoDFoM/68LxqR5VxH+2zgHEKzv0cDionbIHBGvL2W2zwoF5Px5l
f3yXh38ifPzl9a014+znAqEkU4HbIcQ6/o6hG20/hQs7isl/Wt41Gfag3Zt10unD
OqJXEbr9uPAiHOlUrfkc5pM1wY/5aEsfCsDzI8KrdGVTDP8h9L4dc0uo9nhDBrRo
7+6viBzrLGuSxZVHo9l8udAh6L97NWKcTINVzgSQPftMedGNqDPlv8G7/64dbKfi
V/86fmT5o6Qi/Fgyf81bj9wRaUipzJjapWIZwMbiaMZ7yUh/yykhNHPnf9wfoPFP
UupsGf2WWwunjv5ABmRXMb1pdnNxSXLIfoJju6pb9VGgHTxEUrodz7H9Z+V8d3Sp
YYYxv05DC++0k4lG+Xmu3oq69EGU3ikD5WXMJfJInnPyMkgjQqpUXji/Vr9eW+hf
Tx8S6p4QL0H54DMsqphOyYa/1QS5CvIXPTas7arZXV1cdfsnDy3RtvPA4qp9AXSt
s9sGYwDZBkxPVKskDDbhHqiPB20kA0pnFJEuNZcjb8J6jGgYwdyNFPJoeM/tMW5U
SKC/rW5evXMtl/fF7ZTc7BpdEiKiapNFVv9bbXhSNKgYm5Iz9JIY4Fe8UlCdtPXG
RGUlli/sHKwb1BwTh6f179QFkA8qFGzOQNKQLLjoV+TyCol9gvwy6ndanEC+EyPG
AGI6UMVejUMMxWQ6i/Vy6RpVB+0OiUDaVhJ1cDEKa1mv/xELF6qJykKFNEdZRfWn
tV3y0iyLyS4YMusr0GhYzx8N6/PO/NJIS8gzTDZx3v0kn3vbgxcEkT4IvsF8YkLn
mFs7EGN9ESKCz3l2ePqEw2NlQjK5qhBFcabBdCrjl2D13KiO0JaYRlc/quO/6pgn
ksIfzAcXN+AmceQAH1qtafpzQSvuW/VtYlezo9l8P7Zxf723m7AGye/6t8yr4s5O
DBvDNrD/hFKXSYXsJ8D9sEPl6rO40cr5rmdA5RNi20POaYRi/K4qzl2Y27hu+hsE
7iVLs1x06cbx27m9izgNjXTelT+Zbs42whuI3HyTa3R4MQ0/N5EDfYxXysxbbMZZ
4FJUG5fzXr2HGK3MBZ2qyKICT7fxXYIisO/hdb+UXLpnVccVCbo6RBE8kj8J9SEZ
KzH54JozMIcLTFH/ZJVO1CHJtnSl3/9eTVUE5fcA6T8mqN2qnYybfkWdXnfi8vDp
UGcJ8678amie6l0chyJkoySmCvJU87lzGMbKNmPRgKP9hLzO0SRb6KdKpNe8KLMe
dEYfyFjJm9lENDpYWPEQYSMiL+UT9mZrJGV3vVEy/FOXZBTgIzJJ2F2hnpzltF67
/iLDqnJ8LpLCtZlfmLyMlP2CeHQuSEWJT+hH2p6K4PaqCPfvAegOcJVwvF7ZbMe0
+eLhlTBw3hojoZ+ZCaYv//dp0tLEaym3SuF2Melqq/bXGYf1D/y+3K90WmpXNED9
wD5i6djnkCBHMlqGC3m89/fOxWFDI0YBi3uXWHtk4TA4Vm0R1FiNLcf/Bx3Pujoz
Dx6E337e8Ku/qQ5ukC/MfbNTqoOyj3WwI4tw7logvRm+mhH8ePkUoa8g0ujoCscr
iJZ3hdIy3VQ3euNOLBlJ6A9+o9m45ABo+04aD4cVnpWCxkLsxkB6c2ROudtGgdn3
uCw9HbOBCO+062qWH2LY7QdlyZjdu+lAT1+t9ZmwDdvq866AQDPgB85+gzvTFgvs
J2sJzj/z1zF4IEOH0TaK2DBM0zBnWnKi+Y37A9Xj+2LowPvyauMAOoY04nfnFdUD
siH/YfwT+RfljeHNiw5FvjzjmowQUka0MCOFSEc5CccK7JY2R+D9om5aIQHkeh9z
8O1//G1N2eM6squ6bRyHEwn3aYy107c3VUce6iVwDjHeNhjW9X259KAavybEs06a
lfN8zO0zddp/RZTSmTIDHmZ/jiz52tdLsoJo29FI9/wgDQZRgs5QIBKn60qi9qmT
5YWzf7HMM8nmRnTBCeLpeizbZ+J/zwXn7C15IuyKnnlvkwq0pIj8DZQY/YnYwM3w
EOVMMmFQWzTMyVu4Uz4Hul78H47JBvr3Z4cFjY+fo2ST0D4RfxNfm4fKTUoU3iTl
ba8XoFFsRSaOLZSCTBIOSUbQrm+a7g3DDQWsOxSfwmo/sWstvuNxOmKPOAMX2imV
r+22jlY41gKyB2NS4xxMebzUh1CAAvRsdD1WlPrTOulZR4gV9IAaD/pdQMYUQCiw
j6eQxw3Yt59+LEsWZsmPNWfpmFUGyti8dMiUo7t3OLuqdJP37eG/xDKy5Q15nY4A
eT6XoueZXjlOnKCxdD9X6OGR+UmQQ/9D7d13N58MEJAF5521bop87wqxcF+tFmS7
nrb5k116JZUIF6b1U7qjkrXis5kLhQL/e0Yp5bW5UELTiLWXpYRL8lJDTyRSjo7J
r06kz+HglMfbh5U40e6PBhNE/HlsB4Kbwp6vnAZ8BL+kgLXTpphSSK4bThQ6UkpZ
WFtGzQwbnuOr5pcmgdW7+MuefNOJgDirnHrlU/a7jLcz7SGMei8lb9bhWpeS6XXn
ocoMamSKfUJ8D280jc6S2Bkce9gOPXXw/J5sQXkrdTsLdOe1+mdBrn1WYX/r0LoM
baHRKGI8ioWGzTzn3r0jBYYXKkjgwFNAzCZfHkWDvqrIgREoH2L5UIBIbEZ32y2s
EjiD6GSY0MEpmLHHQfEQqRr3s4uKH3xphepeXLR2mX3KkC5gPb6zTWSjN3McxBfa
1edQxldiZyrlM6yi3V7BS+uPS2JgkauKFVs8FmKvmPzhBaigWmMCXEtN3R1D3Npi
sWyPYkGaWPdaYCDc9raD6pVgXCCVupHF9z11UilHVmThQ3pg6pyrpcD2Yv3DuY0H
cPQ9rucSTONw182cpS6KEi2SZFX97+Qlpqjy8jlXaEFneZFor8Q90BtOGjg6RJxE
CkElucJinGTRXqdP/0T8WOu4pZKUVfXff4keed5zuiMO3vezt2SBXf9AFHEJ8975
k6lKIapFi5ugWqa+4tK8vbpW+dXkZDJTBLeGUqRfCh75oABY+gxh6/ESCRp5Gtb8
LlVsb5G5zmkyMeSR5rUX1gypxZ5nDGTwHI2a2h5IaH99+JjAvysB/pKEVlM/8at4
zKIjFGifp04B19V/FXEDnTAC/31QZ7/16HeHuUN5eXMlO2sCBM/2tPOHXngS82Iy
kg7VQMn1OuXOpyQHROiK8MoFZPJyRo1kEzBqT11YfNWZbrCOyNP/81qn7keL//vo
lG3Nytt847u2D4zb1ymk8I9Wx0JcRiZUbxbqKkY7cKxwhHqW+/CWfVi6LO3AeimK
sd2fRJX7ZPpgluklopH+wdYSt+9W0NDbyiXvsxpdQJ9GQKkCxeObgPlCEohTPqmO
GCjH5nBj8jO2S2eYbOncOqfMawMsd/PkcEFPHJr7wHy+jZhvdwhGOC4JYaDkOVHk
R32zNHFF0GRrVOFWU/Prg2iOkyH8MISFdQ4PaBP7j7w/Lcqub8RStL716j0KQZ8F
1bqiyo5t/5ALi4h/YiUvVZOENa50B77QmBNKv6Ms7OuN+oDdGIpAl/TV2FH3A93s
1WTbK7WT8NOqS7gCYeNB21jrUKEdhViSblLUnN/AcE1vCqbP6dl8kflknf9fYS/s
qnqw8G6ZxWHfKOf+sHk+QL/9c8uAB/mqikG1GNHE9EaWe65QpV+6zSZaQk+IFhRK
fq+ZeI+3qbYpHSHU4Dupu+6JG3oEOrxqsbHcnc95oYCafxZht/cLXlygfC7f2NOI
F/7S59wEI3PUIlZ6OVJPuIXdrFiO32o/BenBNLfJukbG2m0HfQzVE+Du4mBevZ9n
LsN+nNk3AOxfxMI00LMVLZtel+OS7BRyit2hNX9bsVMm99tiBtd4hKA9tF37Gn1g
9/MBut28FPLLas6hI2XoJsEFr4tdP7fedWgiQsgADEFCdwczKfmfS9q0cojb0iGl
aumMco+cbshu9+gldOLh+KW8+c90XoNHzMVbdNLFcwQA0qH7mikjTtO/e11WJZdS
7nL9aGY2oNrL4rIejGylQ4u166Q00Qa7qZDsv9d2tfoa6E8h1tgToTXp7f8mTcWP
EgeaBbh9viAWfWbAZiN+tG4ajwVbyT53SIkyOqzG2KOozkQCS1YoWKz6swh8Q1jp
VW1LKsdjvA32+GMDV2gbhbi6kNVcqF6Wx4RaKUvu5juCoVh2GBNU+ePGshg6CUti
U5eI2UkF1DBFEkMf6sAl/67RMNH68Ounat1D2zuPhRBfXbK6mTBcHweOnCpTCbIM
fzXzFaHxGI0a+I1a7bzGVMcHxK7RcV36D25VTetmCpRt3sNeCTzQT9oT5XBwALC8
FIPDekPYB0uO2iXIDwlJLwxMMnk7hSQhUcJzoBHLaW0UOJ4zlpV87JDHuQOAFCSr
C7Su9ZKkh6pMapIK0CXp4OptFRgs8JKM2fjw9lXHicRAAR1+wFcqvXJmpvyiWPYN
zdKUsqja0w/bAYvP44C8VPXoNNFQ/GDHcZNLp3MGCPSFrBA8FzzP78qNXugeyTWM
6lUbGr4NLLoYaaURPMVoIBZ2kvQm25RuHbGiUU4CKB8qIhhvbqfhFbVzLF8g2AK9
zff4CWRmpDBsJGmofcWVAGFIH1mN+9Ieu1ZYZg1DOeM5jdVzOZfDDy+tvhiY7SnY
dXxc5SjY6Q69bzPfwPLn2w4T60a1URkDg4/49u7+Y1KtfcMpOr7HvercyNyhffcq
4/opDP/7WZMl+OXDsUCOAazOY/D4FRF1PdTmFpS6AJUkEHmmLZycaAJZ/OkperO5
RdAwyAoM25drTV4PwrwjFpoES8tsMUwa/rcbM0vmPhfCAILZW/37KF+i6yQZ+dVf
uQfBecjYSGeenDCweGtJ0WR8h63Wa+E3MWRkXRjZXngCtMwWsUl66JSgjIzYvZY4
jqEt37+nhrHRi76xLKomctqsbvnWN4fgIR2aaJyGqI8cUlIap/QH5QylWmhFlKTS
XlBRvmK0NmoLUSy75Rx3X97UtSoJTniJ0nYp4RwJ9TvxMyF6ZWPIIrMymTWOZz9T
ZwtrV+ApKnel8oNOue8NQyZO8F67Bro9xmvPgVMiA4E1P3CKq/2DiFVKjsVocyee
0oLPJFBbauCeoONgXVJMCw7SA8kGYb2EeDHMj/EK5F/qYh6XRKThyEKLQP8qfdfR
9P/vtW4WMSDl0Ofeo67rg9Ax4U7K7CSmxMgE2ipdBxJV5+EqcoRH7A3ADwy+sxri
YyV2SXP1luiLcbgQDpW8D7ZAqnjHjsfyPuyUCo3qyAj3kUF9DQzBnxjpgkfnd2KU
3cWzz1PEbId+m9kyJrltnQtuzU18G9ZRYYBt6xHpwUOhk/8A5Z4AuVcg6DKc4bQ+
eNZg6NhS/8qQ8/3QJyJX44YfynPvvU14tADeoJE58NVJuLykxrjTAl6INcZV7nt9
xTHbVj77U3Bh6TJY56DZ3u/dSNvZo0gWYDrjg+VB2CuqTTESuDoT9QFFQK5weNvB
WfjU5GUhckf/36OBS0bWvgD1vTDH2BjGTLJoURflbtguKQWcfBnnYYmDuBNRIzfp
TiA5EX1zgDjT4xemcSHa1wzNwd/N77yTJc1POvzzvRpviCwlXpNCGKjvu2j/cftr
0dXU4peO8F3xsXz1k2CK+urT7scZC129mbfpFhnjWysAExBjYDrlAhJiWZO3zbR+
qEHRfScAJyefQl+cpbNnvjJF7HB+F3G7QxuZ3Ot8wSCp1b3SIEjbkClo7DWEz8ZS
H+gd4uFQW7qukmx9ix+EoQ7VtwxDBNp8M75/M6HonwgR+XIBsleHsk/48GZxSiF/
BpPEj6sYpZrlmZMnkPJly9R5SMUw6NxfXjOdf756E4Hnfr1Shw13wjZhewjsH5aX
P/3Tm+H3O7uLmov0d5eq6DO2Pt+E51U8nU+Ws4vXJrKS/8Pwvv8D+Ca/eNHvz3BO
54rpq1w9Z2bmkhOor0pYvIY+oNnfx3FvnvMH6xBKNcODcrGd6MJEnn8Td4ckai2D
UHCEJbj8LUu6jNDrkkEb6UPEZU8xLu5/eMvk7QKdnDBbs6OzbzSMdaBRZF8w3361
c3BQ6w3kAlKZXX6QJK19E6xkDMnvWBWNTG8+5RtQjTN9Pauw/PMpy91Mtj1lqqUr
oLDljOAjRIZM9kO8M+PpI7zxiFFGO80Vh1k3sVkeBM3JACh0HDfc8DU09mydrxp0
3pXveY3pPmbKBuUfnsdWUDInnzAM3XQ2/6CkPXf40IluQ31lA9PiUigpWhVFo+af
RAMl0H76lL6tJJC3YOIr9mZBhCtycge4z8mugT5S+z4Ti4lg/RT08cHTQDW0PGip
kI4xWrZKmlKV5GdOUsLz86DWN6rVg886zWZ8MXXg5x3Bc2LBrFns8Z1ddDlmVtKa
10wROEVzYYXrm5kIM0yVggO92F2OdzcinQwT9+mf1mrGxNFOqe1RWG9lnNfVUZNR
A75deOjAPFP5ydpkvbWtUY+tm+1/QvRSakRL/97qSj4AzrolRyVkWFqSQdTCfVpx
9YiBKBRN/tjkyZscJdG2yLbYE/oVDaqFjkmLwnhkucWdOJk+3RUGS2Y7hXOXfzdT
5B1XAncbqItM2rhCKSwb1MuaOEDCBl7P5v9f/s4GL2fPcuXS7eytXeanBnKA/r1Z
YpSYCYI67kdtko9i6ic3ya7BLiiEwOnnfJ9Q/ClqJNKcCPxBZnAZzk+BkKYtefq9
3nNnrxNUKjqTSit3sSG9g7mUiwUU2M3KH9IK+x8PTxZiU5jhKqyvdC2XiaulJDoC
awYmOaLoWqQ8OfGEmUGumTKM7RyuKd0lOmuXd/ztTmy+s5/+DOgxF14/cQMyS90i
bu64iGSsLpd0uAP5ps/X1TAUVkCsWyGLVymjp8mJggFswOsm682rkwFJwIjMS90L
ZRq2yYLW+aGS8W+GRVFp0vJUoaARVZ3QxKeJ5tzLVWwb5CVCyOpYhNxw6SbAjjPW
ImgRrLW5b/bTHSIV4s02LoxPOjRMqlRlixZV+xGpRGRVtOafFYTGyi+WnUASRnUE
9dJO7w1H3/qRXQ2yqxDQYxDe9bx9g9YHcA3futS6qu/dKG1p97R3HQEn9kFfIz76
Eq2qiDPPoTGX/XIAE3BXd6Oc68bfugChRdltEQzdlpWddg4qNiCBxGqplt6H0vzf
PEqH6UPHsBqWnkK9Z7Iyd1p3j1kVkHaNxudOK/3ehwDmlBHIvJxuSA4d9a/wr8ga
H7P8jfkHIQoTPLV3fZHz5v1vS+Dcn7kNs5HaGez3q1Q9kzhqzXV9wgXHJD4JAjld
UUdPVG3JT8hdsKj1i3Ah9vnJSW/upDgyvbuT8wCO5tJYprwz3vPeEln4XbnYjuck
aDJe9xeDHFvFqNliMl8MeRT80xENfaTUVa0oqDl8sHM09l/52VnDzqZFE8gy4+/l
i5ZokcDuUtdB7FnfR4fsCB1Mt2kmOQeulZyQEXvEO0irmuflHXM1zHAQHAlyhOv+
eLSmGfOCsBTUE8c88cARvq+IGIuSW1YAXuu23OOcPr9Xdb0GDi/q9vAmshZtDT91
vbmv3ytb+SJVYL7ZzdW2Xdo6IXRQgE+55HiZgCYxTx3e5JoVechGknUAmbLhQHqB
WFtGT/SEfyWAnrFKfgnBy0GYZ2bv+jJcchxbMu6fxMont50eOpRGtnhl/zGocmma
2osL0MKWO1bLGqn3lbSf8NhtRqts53+4PspsX0QHZXciC1jxLiZrIJrOijGwckbU
VaZkvb3R/jYqVQn7wAVkwr70InVJt26lk5Q8pX4TWWORHU3Pjb+mdFtelIAzwWRD
j4yCl4aA9e1Zrn1s6tNGKwJhOvQ7Hpjg3WLRAGELRdyy1iWlv38fDtGQYl7ZNCn1
dCeifnzNaWQShsiMxqlOUH2LIvWvngzl13chkW6H8q5usfXZUQe6rtDwKRTffbXu
fM+q+rJV+n07/l7+hIkR4pCwanOpA64kaJZ/2zPC8hgvNmTv8hnLuaF4+Qw0q23p
t33xkUgkOQ1HCo0Rhoiy40jDAV8ssvpAwpa/8sxIfR2WE/xJnjIfpUu/lbjcJInI
XK2pN9Hp2EQQgzx7a134yxZTMES9tjY3tOrjWwYxfu0opiRuVOXRQeyQDG+TbaV9
KteQMn+CQahStuG63e3nb9u7TaktdRyrBkbcLUvUnpzff1IcL4gfdKn46u7I+09p
xdCVSbwwZHAvYD60QbSgu3FtjvCS6VuXhdUlCCYg4SWJ7vkdMuCdpLRXeTXFcZKW
K+oN/uQRPtSkOcSi8iZ6uNhT0DQ8v1ikcp5VNqdH1Eq/B7nfhJTXsdjD0bHUbcNd
J7FhfsySSTscvaJgTsAK5l6qwTiJDJv0Ynk/LOJjDiA6/gMLXnosDaK4pM4Ukmsy
CFLbqu/ObX68IMIdyvI7gdgzE1PFFX6iWBscxPUSBfPS7d+arOPQnwv66zlaXmAx
iGIZoqbz0/1ii4t8x62FitwP+a81nrWUQxVmvSyRPwIJhXvWNbD8SN8K3dBywqcQ
21ETMV+PlxdVnaawcclMTyVIslTeP5+vxKTvjC0zqdMfLhdy16C+8EaZDG9q/X+8
NOKSfNFDKvLsCxljlTGsTXV6AgPIIGcz0aZrqluP9Mj/KQ3rKYzu21h9+QySJa57
erHBgXwlDFmSSd1lQ1I2uIK8SPnKZK74rm6u/Vt6WJeu2NVhh5cF1k3MIJDxirmP
cRhJmr87dEjVmCH9jiuakbGlxBozgthWUYOZ9boFtSWjNvtC/tiP4FpXrAl8iBYR
/fb78wtVD9M/IlJuzPe+w1iWERUZm9XZwpXW3u1ofn/AoVxaR2WTsz9gQGqgTcDY
Mh0WEvjcXBAvpi/vQ9sYmSd+EgyKig2ukpL0xJNK7A3spMDsMLmR13CF0UnXCesr
4yQTtcOahmz6OsZzG4PUP6mUQMNjxPKFf8Y5WGQkqaQE8bSWuL5Ysjjcwv4SIR22
iJzx0+4HyXl/pL20PXVsD0PLmFFwPRKIBf9quBlYa9hVjrc88/lPGF1d5J1NZhKu
wVivScVuv7EK8sGQR3rkv6bWKSZ9e8IeHTjNnbqtLM84FtArsCSI1qEugInRlvNO
6pYkn7mAPYk0dPHnjeeeu4Z5bxTeXOHGPA40B4iYqxAjeGG1toDP8dK6LWUs4Ezg
RjP1+QikkKH5fXgT5df+J+xPbaQ8fNZtChgbiK0lydXugzIkDYHyUbqMxXd57AlU
GfkIOGyakHQdnsYsqLxW0MDHsCgp1TioRa/Did4wj0f3cVAlZQWZOZ3+FwQum664
d9jI62OXuAjr/WjeSw6x+Es1kI4+IUsP/td6itKViTsUd+6YgJUKNxmJZ4oAn52d
pBoBW26wIw1qH13il+rNOS0pTj32MGWpKf09JxmfiXIvCb/jAh2n/TcD4rKJiNhA
56brzlGStH32pAmQbf1OP3Ty83aJI9wcTNvOw+BO6CIf+iUnSI9XqXsX4bLqa4fF
C9haE+PwpEwzpvu4slRqd5QvKNx0SYkEHePeECoHBzIzpBwUa0ecJQ40eCh+CY9o
avdOL8HnEMIgLqT1X3kVvD+2WSzPqxXYwYFROwiJICzutBO0tkTTOYqr9281NCN8
2wa7s14BwCyIsKfxIsidG4RRuV/TrF49YUatsSkkNabsvxBc4nV9zn5u+CYbAjVc
hlUaKy43CQywe5JVEnKRyDIK2eVcw/+MFOTsG0hN+j4qa6PfJLR5+VhbqrTQO1Pr
B+0c8c9i6sn+BD/6M+ZukfH452zVk1MRske3x6aoWvF7QMBYfqgtygp0pi3WFapG
vsnJ0Adi0FCfLZ0t7UHbYkjFqKbhla1LJFY9h0nQ68u0A6zQj8yY7YMPPU3fmgBW
ePcXSMBvqo3rNyp9fA3NP2Jgrk5P0DFJtCynR7vMvHauY6oc0olTuKjTjgtjP1r3
LJpr4ZkTDKglnfOXU5d/MbtAkBf85FiXTLxUrrxG2O3UmyxSzQpIoFrS4tjPeRBE
SAUX04w1VzeUxHAuliYSPvnmP/qGb6qkbcTo0MLKy6W08vJgNXe4YtVEd8INFYAz
R+Q7B2fdBIkzrrtu3VRc+iDLjmpka5kXy1puvRdhY8o9PBduD4HyizHAjr60xwCL
PME9OI2BltYrUt1iNwa54JxvLKv74c2/1VQudnVaMaH6p2a/6nucIeMluSfh1bWT
x3nKK978Sbo51z6h1ZCfBOt++Mggp9Fmn/tK4rfVP63qIR1385yoUYkU9SrkQ+W8
GpI+0C9TAP+TrJTlv7kXvAtigFAwwKcGvP3xI54ZRbN9m4YhiOe4SRq5vhwcYNkK
uHzCUwQugA/QubKzEC3cP8Xri03087XJ9efNcZfo2wi7XtesakUmMwygJmcK534M
qvMoNId9SWimqN1yOItnrDB7UMAHrTBhrBvWyln5PfQ7971VEpGEA4Y40l6dnJvg
0qNHmxR7VNMzmxAr/8oI/3mf1L4UwsIO9lLm8RFLLxOWgRJBeYojd3HrEFAdq3JO
/eyIB+yPtbTj3UR2WuEwAzFiytQ1YjcqMLQj8M6ScuO6wuDkFYqcoJAG6ffOLxHB
1iZ+fCbiAUeSu1XRCA/pYJCRkrFXE+JjIQ0MMLQmzu8J//5oxI9NFuZLIbufIyZY
HJjpHPdn9hgku49uYCAAFC+Q9apiaNFXfRnRF5jd0WDw/KyO29xcNYZ1KXoIcKdh
w/vbPx+C7SDfzXBk5IsrAmOJQDz9eUNerk2fKZVEkP4z5Hlz1HOz4U+mk6CVyX+1
97OfDtSUvw+g3aCGQuS0I/preJVfQHdaeYi+QhPkhjKXmNNdI+Pr8aI/luneXHgY
qJdX4WtoEmJ6CS4qYVePmeTlDBQ2RxWlSvle497jbtE+ixRrauukPwXqLWf4qjcl
pMTChec7K2+avmuip0WEn86NNzAGcHU0VmPlqDU0ifU44WCbKUSv2GrzvReasP4w
+Kd4Pk0c8SJWkFmKHfUnvxMfM8/31yj8WZC3/ZGzrWgbhmWNxqWqR89VVVrgB+U1
6FO9fOCZMfNqlhmGYA5iG4zfbMCjq9e2IZfPfTKjdV5CrtkYaWN9q7j2ohbUOlpI
tOQBayEd5UPMnJSQbDSoul4el3Q1U3OWH4KyHSHAOR3Sw5x9EVFJW7d7j83pK+fb
O6n0x7JA/35VRxz4adySPy3mOgtTg8d1gAvGsnKXI6jkkEA31PW2P6SCi9/3+vkL
Bf0ccjUHH0zG96RDuC7mfrFyJuC5TQJsO6fpqcHRglF1+qcFISu9vKugyo0ukIJf
xr1FDjaxs+qeRiME3X88CdDMz17B8yK6gTfLUVrgiCP+k10S7mTGv4n3G9TpwsZz
fekGNSPnTycm9eCKRZQ2ehNmXV8PEtKT2QP07KdyzEMSzWxaXRK9f5jcrjQsFTbx
KiK1lKHvTBP7PLx+K3BcacZVK6a7eMjU/751PDRfsA0wbbzKHXqblAB8XdKTSZUI
om0cEBUdpRs0B9nFPyMoBfN2spBboJUUtmCUw8co8gsUNUmgkcrc/SwN3EXNX3S+
mdch6HmuhHcLvBPoSkefmklFCSzsg5tzwX2WOqUIrjU74qrRpcfP3l2LU7L/saEw
RdRfYIoQobvchxcnXuX3XaAGQBxvz2aHXcka8m5GQONpKxl/t6OikMZdEzk8jJuB
caZhBywiO61O7P4dkd9p+0j9FGSituyslHi3o/gZszps77emcsLFqNxBAU4MDHdU
C7dGiSz9q/g/pmxXO0zPfJVhuQkgx2ICS2OS70/ceuQRs1XChj9q67qrd3Yk8bDA
3iXPXHTCfQP5cfIhkoQ5J+fOmwwhCsnVpmoRe+ICY9AL9UDyaGCzAoY54ZArJONN
kpRCDg+I059aMDQhr324D3uTU/+ZvQd5KAVkf4uT/So+FB1Noy+PIrCm4b+fLS73
YqLIwUrp9F77abJ0ddr8umXmCi3xfgr6YsLg484guwDDv99VzQBBXGUEA/4kC86u
Pj0bxTnAD0dM4HXqFdf6ATLK8WixrWq1qiiV+pRfoP5be625M0Kb0Snm76KyFOeq
j18KJV3+/Z1fZhOJdEt9Sh7spqqnSV0aFHgM40AUj+/E/ndVrpA2KpEKEWzB+WKh
ofxIitBbVaXB1SN3hy5tA0u69mnHJDY0i5WFqwrBh52VM6dYew8hf10ZAl0OtfNP
w3oCt5dPq640W6X3Biq8eJxRf4dunV77kBAzrFfFv7HPV8I4ZVwwNBoruLCYJmV1
9JWrCh2qqlkMLbhtEn70QCjQ/s0oAHzrcC7/elIKOyt1GpY+yEZFgdDb658tCGFG
68djYsCUfovxff5ioymYq09XXHAkBe2Pq34l9AwiGuzED7KlckaHycCst4jK/0F0
PQ9gdt1UyQFmUms39mlj2t1bILNE8xfBarpod22AVLW73T+tSSz+wHCPwCfGOE90
6CFbCOM+D32RE5sE00BEwX8XXADbGY7Bh2D2jOPXdATmic4dpFEEdllIe/4OKUql
25nzHIRiAJbX/JcRSdY1JZSgR7hhXtKSUx/mNF0sZwJ1IZ6NIA+glD/UifJpkJC2
MGiqGNCupHX9Cg4WKSSY7Bf+PJTb3tK5HLUP9maM5q1OsIZv+2PKP+DELfSJJegy
AtMMBflaJPiPMpo6lCqk8m5RVazbqaoGJD/80igwUPmF9EdKQ6fIjn8X52rrSx4L
ELv9JswhIhyYd6/ibq5DiefKoMg3/5NrtclmLYK1f4CxZSJKUSv4s5ywFO0BgtDg
6WHEyfMrUyRO8e7bHg3Pk6zbItaY9UzrkFLINHlCUy1l/miyMjfDiY3NLjayVPDo
QRsU4+h2i+YEQnlJfjV+swCAUPHevvvSpXdinRBUaXwmq9v/SUWtCAPOHkhOQRs8
m17P53gaWN+4yGB4TMiw2SlZXDDqzy6hhhRiDEtQPPHCMeqQJcKADeRro2I6KUrq
NADZ6M+joTmhi9yzHEU9CHp4G7UJWyNdPJXF2+ONTtXhsKCMKyTV8HjKVnnH3ob4
9v7vkwclZgn9iyWjqochekibyAuwH0FIXE4qGG8GxHIb2lKsZKI+VDXq+sp5fDR1
t/LSTQZKEjSM8N3b9Ih6c5P4tSp7vHK7AcJrzlvNtU8ofJO/AZmhqXMHU2e5gRpt
Ga0XEPeQp0r10Dc+ByGk9KErN62g+XeVdH6s1eeeTk/vGbx9FKAvSzQ9AWO8G42u
OWw2lDZfE1kYx0Xi1yts04C22V3PN3+ZkldxrX+/H378zeVGx8IBzemyze9ILdS4
mqz/X4gBT0BfBygyD++Wc+sYCFeSQSdNVKz62LpXw0J1Wwr0rZpOrT+/0hl0k8q5
GBU6qo8X3Ray1vFfW7vC8uggxwjf0QxRIHPaiz2T6UVmOzOazLPs41uh0kXEf2Fh
DLFcLGttZqjZWGaP0KJZZP5N2XkITFMbfenK4P/+Hqym473BX4o2O2q24zB2yV0N
UJJ5BnMjelTThNNWetPYuhJ3WjnuzpkQb4V9Zi8KnPWQ7uD9UnKgcGSIkAVf9izl
BpoSp3kWNMccai5H+vNo1u8UCRCXNpRRX02e87Ptu/YbUH8mooz5LJnSxALPSv6e
aRiMVKzX6LNT+b78pmsuwCQggorrt6TOh4MRxUAZgeKZfVfzXgwksKWw5Orz7Fbv
CLB94WuaQtqF19tfv6Jf1Tlh2YC21D9M75jod45LILopjALVo2WAv1wTEMci1NX6
mQxYWUT7BxZzUdosoyT0Eyo+Zwpd/lC1QT0wc9qVHvvStRTo//mdt1OfCX6IhLrJ
Vlkqa2ExQE+HnUWsegISj/6HeyPeARzKShBrqdkILDc4vgfryjbh4XSAK4iRGT3g
IYFnBGPk33fSi9hUPVQOP7+wy7a5xOb0tSSS/4604VKC5aE1mIKsvuKzez/JTUxp
ZQh8wXm7acZkqEh+9mQ2VdcZzmOXQCmbOoqPncPP3kNbIOgmGM/pKQSsElJWYhiA
2fd5AwaCLs3DbPghk7NI3wrgKs6LTWePwEYFhFiVAwDHa86H7+AsuT7lz65MtQJA
n9Vv+5OfV0HyK9yYmojdk0u118fIWY+YyBsRfDoP5gmxcSxhPD56nGyUuthzqg3p
ShZAQlpciV6nd6lQg63wx0PzQRXfdMFiYOQFWwdrdSN5DJ38TQ505JD6jodxVxlh
MFHX/PjufMQac4cSJanq1efQl9IP8d48KL9qox5PaXlxVkmBYenBSGjBrCdV3hVa
aAwDiToxKzDnmiBVTxWZl4Xamt47TnWv+qPr1hBExfR81IirLmNfoUlQi7eb+KfW
jQKIfT3X80v+5Y71BTLHYIqTrQA4Ib3RCzZyUBH+H7/8EHPmAZ1d+snIgoYsPGip
mCQn3x1AtWb+qVyikKxJrAioakxLCtpt/O4ayOJiX1ZZBfJ0FhjGb1brAnsCUtFz
ADyp783TUJn+/VMxjDiA832IUrx5jwey7nQ9gfzyIvKZ/8Ci5o9Wm42OgxxjsP8P
YSASWsAnU0VtOlh+Rzdyn/H41T/uQsuxbA1O8ZNiyFB2UQ2LaTdGzhn57VL7oP+2
XigBmOb5c20WK72U36yONuayxXhdL66VrKVoxpd+AoOtEuTuzzglpnBppAWHSSnR
k/XCre8s0y0igMOAubrbqoFQ8ivOPQXYZMKZDhsw+DslZoIAqRRjcXQQQQjVPbPA
x7UVZ3JUwjgV6fP2Y58il/8CY0dB4egJLjQ5fe+ml3A8y3ewknpd3uJb0O9ecX/1
MTsC6p+iPcFLnvJT15PJPCQbpb5ULlmKexmW3jeY1kIZ+gPquYf1vl2Uo3DM1yo3
JReUICQbtrE86Ky1EUcMdt9VOR6kAEWISygT91T4hcpn7JrLyfpoT5IzxF/ez3hl
rjKY5oai+GyarOd4GZirrumamjmDqiLOHRbQ80pVI3CgoYUmMmqP/LIUwZnNFlyd
CmS1zJpjtG178TY/IQ+NIK7rtysTCvZOgAZfjA5V8Hv7vmW8b03onJXMNZZbLEWQ
fQHevFmbhR5/JQ6f6bQgSi0/KcTtukDsvUfzgM2ARTBUaAbHvjI1bNIjKBA+83sj
wpITwZWLFvaux9Jmm/6XMViB+cIXLHftALPbSdGH2exnp+EnU7or2dRb1r5BkSOM
z9pJRq1vFb72Y4rePYfH2jU9KcbSJhKMAEpSWt5kJIX4t9Qmqf40rOGIOObjGKz0
U73Po8OjUWYtlNipRkNa6QqMlBEO48CPopWuFrv4h3vfoyBqn/eVGXtkYx+ux3YY
FzDiny1NuUHIXr5UPux2YYhq+TkGtUGxW/odjt+J+HvFT3d4j2nMN7PDe5hmYc2/
SCPLGcNO+7sslX7QD3dcqSA6RxrBkFp0KmqVPyPNkeYn8JUKG4XRE+wMQtAy6/pl
ovhwCOekhhsUo7lT+6hGRAZxyfxW1spvCEkNZLul41z+GEwoVK3LDijvxLxw5z4x
nRSrHFgCo87DjAsEq8306FC01+ChprOMbnw9GFQB8HK9Xwj3oTyQWA53FGav5M3c
RBOTlMPbPtZfSz1jBnyACQCQ+bkUt2abMVspTkyuL6dXJKRfBCeJ50lE6w0q0mgq
Qd1SBSD5mMyc0MLiaU++hPK9nmV47l6mfy8piMej8ggKli/Ia8+0hXIIMGMv3jaZ
pst3/ut9BnUnc9lnWpAJfPrw+bROqnwIzudLDU6+RoDP2C2KH4Y1P3hqVnt6Cvbo
tX+C1SEHfzy15Ee/ZstbW3tdRs4LQjx9nGGzEYrUwXBaHbE72R+x01iDgN12s4Mv
q48nNXwOdmQ8mVwyVGt++ym0aHLQoAWPN1dPpEUCWec2YPP+5e5IV0dBeV4tPHjs
yv0NC7qckLAN8DTFn8T8atmMRIF2srQNM2eVCjWsPRnMtvsNHF/blxaQhCMkAhR5
gOMjQPxNKZ4Khz/GMjn2dN61f6DmhTevCR35HPDm56+6xTFjBFZBKSrY4lMDFiOr
+JXgECpb9ucGaBwwDDx1Q+hsJSkX/u1HHNrPvHby6mhTRV624WQH5ry6i0XL52VV
G6rV1UXBYJJYKqzC4TTwqSIg/CHsN6tjHAzWsx49JExDQZevc1we5bEC9gO/E/PR
6Gg1kK2amKLzU7TJdb2+ZDal9VxAsNbV56LToZ3pTuqOyzvAbFNvnMmc2daTvNkQ
fHrdRt99e6XzE2wbse3hoLnB7E2JR65NYOXuFBWK5bNE42xnRC6/aKZMvo1dL2fF
PuBBtLzE42Te6C9Ty+2LmJEgjpwmm+ZyV1JPDIKypk9vyyRywtaZimZj2dpFjqE8
AlL/KqldTX0qdqlhgNQCGm1Qs8Moamao4iKD61rpiNGeqYBu1pjGjf6ymLvK/nx/
LSAuIc+1afUmENDgNiA5ggpysmT2U3bgxIB7PH9NqpNNXijJj/rEFVAiMw17D7tH
1xuDtVzfnJ03su1JlQf7WoY8Luz9T2KeMZUTHZguVT7IBXf5Z0MSysXxqMDuFhNq
hPziqhoUB+Si8fdYqZ/QI9Mt1Lv3t8ZLICVxSLmlbzjNk7DjZKZZp8QW90KmHL/X
fgQQmq53g4aE+KJlxZhA0HNlPcnv+zFGv6wDjhsZugY54ZG3+zzskAHY6bmSEadY
f8swMBBs56WKwjmb2LgKKpSYzWO7YYa2xacQ3XA5+XfuNf/9kojTqNOzL1NBuuAi
LDm1GaapPXUoU6dpbvBdhjs6yoAkXuF/njqPht1AXoKmQrNoku/Df5NStm8K9yog
QnRDecMafHntyvxkK5jkxzS9/I+PleBUCBtY0+K/JN9kc4/pQ3pAE3w+h6nlWuQ3
KpHl2lC3p55+me191MZRA+gEkzMv5Zcp7UmTQGAOQ/BqBLlVEccCt7fFa3Tl0OID
8dNFsEMSv563lJjOH9OmpswPbEanRD+yAAu5hTQ3GzKOIxF5UqnPu+/eehWKtrma
6tnNi4d1XpVVohHagIfTFchyaRQWX+V3CUo1Xnv706qmVWpqNpAaH5bVDjoskMUb
iJC2BGoBM/G6Al8NwQaRGV3Y4gKckmwP4M8M/wDa3GWAXpEfvMyZE/z04uJNf49E
qDyyzUM/TpWsCmjIrtrB3jJqEZiNROvms5VRUCRGx4EZHdj/K83W72wr8hxeFmYo
60OzgNwp3b7n8CoWttVVPDVJnqcHaUq59GWbMJcWG7jTQEjhkz4qz+BycECWpZt7
Z7CiDdRRF7I5I2BFG5HC4REUOjhQCgnquwRUIyJhwiWsHh9knrnfPxROPB03KNm1
8xBhhh3DZzEIvLN/OuUXdUrPIVpKuDDm5C/P9WJ5anCHstE8mCJ6t5ktGz57dBpS
ndAlJkBVrIA9ybvVNXB6lSWJWNhWwpFz01cYxoJeyOLzIIJzvgQfCdC9dgrJRG5A
vEB3EfcqmcsEBNXL3ar1kR3WBNXYkQP/EA8N/1RZOiiJzc2SfRXrfAc0O3HytJWB
IRbx/G49qN1xyszukiQ2/FFq/Z9/9kcchFnLMfoy2CAUiXjhyr3IbJ+LGo2nkIXo
V33yAr4mofdVKQ0L+GDed4ji3g3VJANy1MD9GEirbkniDjHa8AlfeaLRbcZT45JZ
roNOM4pLdoRwWb3rJQgGSMPE/Ce0HOk3fzckUqPdCPeXeWJFk7t73Ks+BMpBGlkH
q34TXxGBb2/2Xm7yEU0riJtoWUq8716pk0m5eGhWCPMDESKgtKuwDMAPKoAC4ikb
3FdTsPgwJ8KB6MtvGSDx8aLihYn8kBCCVNe0FfpVWeJ/GxVWE6QfFbsa5eAoY0YY
wyOJOQxqERwt3eX3vv8I+6RYRlE2TdCEBE1YR8cUuDwM1MgLovBWguL6QjsAi733
N+xc92RB/nYrob1TWzI4+rwqmInDknTdBFclF6jLyplWpxrgMiKF0Ot1GGvGYC0o
O4YLubryN0CiRP1FeVnpagDXn4tln2SsRb1BqXQGkujcg3h6SMk5nMntKCPS2uKZ
BhvdX+CWFTKMs99W0wmLHi8Kz3t/yyagS6DduQdSKkgRfM3OS/99Z8VlHAn6u+bE
DNxNs3Ugna2bWUBXMHSCrzylAm6ovpHazZ26+3gKzLzYbXIQGaYl8oTIjCJNRWvK
7XmH8Ryn+k1ab4T8mOfvD+7Wx7L/Ef+NyaEYnWEXWvewxjthrR/pfmzT7MuaXEPl
DwYzLaFVV6p1UWfdhG2s/IcTFkrnfTsmmSGWKUc3j1TV7NgcnzuUSqg9h1izmOb0
LCDU+6Pf3xW6IZNSzIw9L9XWmuHcAyJWhvRJI2ZM2Gmqg0957cnDPoRBmJrQ/1ZO
q4IdRK1BF1ks4iiFHtosI+YNjLfBtFuYoKt2BP3nKgkymRPxGri8ckL+dKr4evX9
JxKS/St7r1FD8PA7DF2QiGjnw3N1pN/rcqh+MTo38dfxqLWBhT0wtifWg2Mfz0Ar
l0Dq0Mm7YEr3Xf+YBACeI6tRgAmpWXDiZKFSCQ1tBB1pMUhK8HUJ77PGWh6/zVWN
lMst/nHJDtjwrNYWnwFe2aBiIG6LbvGibSblcdmKTPpHgmA94J5GXgh2mB6zQfs9
Xbs38y0qzO918t5CkINwX7sBv37zwBII5+woxzLujHyV/29PzFiluZrQZbI4DYYf
oa5cKxpxq4l1IN3R0SAQi+pohrU8+t+O7OFLWRqChu08ImarMDlcR/CWAoEiyNnD
AeyqfvFCwGoA2VeD2B7Q+AfKf3LIrlrFH7W1qGPTT4nCfMFJ63UmhA6VCUJgyy5V
PRmqMTudUmZ3OEBTiW3NuDpnprzUJOvkVduUrQnnczkQfVV80A6HYqA6TRcymJpg
PsnmGGEH0R7fAVl0WW2S2eSjRIduJTnti2Mjr9SU8DKqq1iarY0Lk36Dj3+ocSqI
LTjk7MeVmms+gcp332QO3quzynnx4xqd9NESbcp14ztNhnUn3gxBUBQdTaGKg8Zb
VN+sNWH/sD/W5onKsk4iCiIkfzeSDJJLkF2OG7VO+EuBOFPakJeo00IQzJkGrPmO
4F9BZ2ENM1n4hxAgBd4JMRUMn9Q2/jGdOfiVOXLpx1LXNQ8X16aAN9abls/pgQrB
xaiW0jwyvvNtJ55LkqNRlaVqJuGFlQdfHWuOx6dNLkCWOmUnKMoDx7ioTV4ZuMD2
xevIpdlt1makLUjRBKVXz4kMS9K7fNxf5fr9ybQkg0VZwgbqyouhGK3QG7LQaGl6
3iLyplZiOkBJPu88TWy7QVLv7U1Ihp2j1gHuQtcBBuUoCA8eRixews5hzMrKkbw6
BUCjyYzjNjA2iHDSs+xu3n2eQuhvOLkV/qZYQ+AmlblO54cY00XQ6uljFh64/jFo
sGnCziEEYygh+QpThUMMPBZ/pw0IxlIQ3GhIAlVogWIXh9F5v+qt6idMtgoaT23P
otfGBxP1l+vorWd8tTvmChCXWZYOBxIGJ88hFcQ6MVxFRHj5nJ8EbIURzLWf0d5D
7QcREk/64rXG9fOF0dx42439jobxMToDBbsZTd8gpbO+fjMU79wi6KYZO8z+A3Vd
s/JA5w/mtXGdYzRK5OBa45ntAfBQ8QSHoy0Wl5xUrdnxVgeMmsl8mwhFcMXInEHB
iij3dG082ZDlThW748TMe6Tzpqjts8vd0/Xf2zzXug+UoLZic52RujrbRDzSy3HL
T44uEs8GTVahCfwPek5TV9Pjuet2xMINflvbmR6PxC9G86RhrONdCBNx0A+BnVgD
LlF5S9gz8Z2p/mU5iqtADx2UikeadXK/TmQ46HCe6Whc0yEnGq1uvpKNI3kX9UuO
C0IWPGLanGYBp8L2vo6clI3hdKQeD6p4Y21Nbo2P3yI7WPPiL+U5i/nxCCIZADWq
sRmNmsOPhYCX8xx8SzWSi7YGizwvbBo8VmLdxc3RpgHt1o2Q0tr5+cj8oJXl7dh8
mX/58hsiPGEyjDp6pdunIFaTQd9a3ZFoqF5tO7Rs+zoCXc3BT9sBCfwOtRi7OY6O
hGhZdp0U/k65sBpOT/cLypMESVCoOCL3xZRReFikIdzf13nyn6ePUjp7V5hZg1/w
GzYmNezXxYmJALrqcdUN/3aNya5Xvn3L0+KKi5NgAmz9lCk6TBWMJYMaoyWzEAbu
n1z+zfvYkIwAhAMVaBehswmb7bY22AE9Bwl82XnlIqlGmRIRTTfUEydY2a6uY70n
1k8p9LYgXkoKlWeON9oFsm0c9Jz++D40nJ790liBcWFzTVGmMOKvTIySQQgMuFod
1yx3U7bONRjrXCIHlXLsPsdxwI++qOMw417MkGCgVLSSYk3TEbnTc7vPF/L4Vu3I
yG0oA5roC6zwnET7Llfygh12ky0Tcgvjb0g1jstckFSPU0dNtyhjM1GsjtBKGhHo
8BsK+QFBeGTJo07Aer7RK2aqN7/ksBsLdo/x7Bd+okECWnHHIFuxvPHY5/CiueVA
4E4OEArVR9+WThQi5eXPNASBcGDQ5rVMrv0OXAlrugX4ZHCjXn1EdvuKGlSw2vE8
fskZ0M5O7vbvz/SHV9Auq0M6EMx9ra/BaoGeBvLvIrWogDof6hdN42FSq5ApErwn
ix31b9aCzMJ1pQl0ofYHSIAH6mToxSx/Pne2+Q+F2EhsaAAfE/P7f9gwuAe8hvGQ
WV+vSf+RKsNJ0t1+N09kVkLk2FfTn8F1d7GKd1ZVtRAKXzmkp0ZxWA4CrweshPRq
f8mi5HvYwsk7XedMGuWZszRReHWvaqMfAMyxnzmDDdOA7qSsJ106GoRQ1bMfTmj7
ufjkoYYk7yyYUKcLlaN+OWIA0nf5hRJMiS5FAaFDVl3SThK8WYiSCnbFQp/M3Ijk
i1jQyaMObj0EOhq80QB9jIoCqJST2yS00b0W+hbvQ0uCJWbi+fGWS9wJEp+jLgdI
/kqvcAsy6yeKEE5uddoz7nSeIYIVeWh4TvQFLBemvVJGT6y9YAyJiJWpEL8dbjJy
Imq9cs+Gd7dwOkoJQpTgUAlBitIpnJT0UnfO8fq+N6Ekff+83eNW7hICabJWY8cN
hYLmQfvJZ5OIK/PykAgVdxHlp7AXVWZcloikk4ZWeOaGMx8OpVAcXM165wkO4xFx
cXbR+hXFg0/ZAT38B3XpPOTV/H4MW0/DueIHB59V/5XSaXLXxAIVUE44IBriLasz
r6RqXDO8Ergo6HphYIIJVcxdy6mRIq7foMBFGzMONLTSkg/m+t/hNWO0i+IhImjo
f1CfZL+AJZb2W93qHAEJZ3LD93VWrc0d8OojNCGcsQ5Fk5lEWdHN9QPiMjkaMS2H
H83LR5K9SUP+5p8zNX/3wcZvQ08ueKQBWbtFSPUW5ff3A+YqjD13ZcoTbXa1+1eW
iEPRibwB4ROu1W7JFA2yBm5RRNs/EsmmQBlU2+9oV7gSxT+nYPkrZjdhdwAMs82C
r3d85NjRISDy+WbM+xSF0YdKg0Vd6jP2StbYiw+jSO6RVJ16ckCS/ZMR2YPTNvrO
6YyjH6T7wg99y9WpUXvZZ6PBDAWmHrnmeBr+MQ8Y/qON688rcBpaM5nx9f4peDgR
/B+gFr5TdsRbeyf+t0DWvFneAOsfuDIoFp/lFK2tbd0kZe6pSK+aFT8XInYPqhnW
a/h8Zhha99KqOBkdlgYiiXggG7OHiSeo6qRlGstkCErJElVeHrVR9XWnqKChul6P
caNoA+HK8iAurhtY5TQkIx5FxUW37Li+2mGfBCh5XVMEOwNJn7BdYnylfXE5mgL6
XS0hwdQ/yImz6EciFJ/y57A3ht7SGq4ifBgCw9CAS8NXzchHOSU/F7IZJIjGSxIs
zwBY8rbnYgiU9iEDwfD4NccbzOMbYu3BqBu73TCNZpkWfUN0mdPtkVQ3IChFMuQ3
KCA+5UnURV5GAcJYPsF1mpBHjAgj6SGHdN1Bwa60SuBOgJkrbZ6gF39eRcYsx5uc
oOw9WwDh8rNHswL56PV++FAf6Z9OkHFHTpCBtEZoM5Oz+L2phCsKlJAZ+REZHrft
tkvCR1TwTB5w1HRB/bP6vH4hougmgKyv4DjNJj9eEdm3lbRPNM7JySL3MQdYFA7Z
ZQ/bxWeqehXB9Wn5uv38S6FKOiUyzzXewvmjY/83QX884a3wsh37AjHK8FTP00oJ
ZwcmlCBmF3nTvNtg4VjDYGNKTKrAG1uMF/PH0VlvfhNJLF94J1N6HCgHc5Ik20tZ
eP3OhVX0E9u1DuzcrlGR2ba/vNvJmfH2CdFVazOg+f3wQlM7Y4R3CwWFaOAxEhDb
J9GpLQEtFsoWvC68vvVMkDz8836+olz+oNkiXUim9lWycSxDUp7eXVHlpzJgnBvy
DhWxzupukCXHzPtYPNYD0w/c0x3yQPGEnCghHAaQ45etonqL0tzxgQ3/QQmyuE+q
tQ9P+i47vaV6FC1+keIjiLMLSlcPr4mqomzmLeuL55ok4VpOXohHADRcqPRBL7/T
ci1a4YYeOi2+ZUPoKCFO2op41fI1oPWDBJYioVms3hja7uZCPUhVMtabGLSWGExv
Y5WCxXcJ76zynCL3A6VkyxvYJW217v5XCSKxGr5OeXNZk7WatXjvKI8H8CKy08UY
ljFFfVezvQ2yP0J+k40ytO34zu5xPUgaVlGa5ADyjGBuIuAo6k56tir30jAx9+bk
+j0Z6PRnNuswcCUJNh3kxZYd3a99+QeZZLkuWz9RWKl2WiQnQPZS2QOhKQzxGzp9
G8yez+ASNCPudvQaxs4cewz6FTWZeKShwDRj8+0pNLa2vwp2F6YoP7Q/+gQnWqAS
ciaeHuT1mxnLfQv0cdSgrLndO9/pIMa3jinRbmU9d30NFtNgoehRgPjGwQnDZ2hD
tZlT+mZ2Xj6jZvmprQlZJY74LDDGueiKcgF8CZG8jQSPvSwBFXMCyieb90S1KXnw
Pqchhp7okoyiYj2i4r1PZiotpK/UGA/2JeQ8T8tm8eFfwVTMVceVVxMydfBNFWQU
mpSs2cq/FzKfvibZQVfxNhgci+uzHitGY8UHk+R66sEB1gb8ElbEZ7YQyPsN8JSI
BDgyXGTbza9shnk91pkfrSkO07qYdAMt0N/ZUFjHCBnGzkQQwpJrburfqwFpd5wL
r36talKf1ai4m29m/OR0UJdpkN1sTqmGce6EVdEoygz2GolhwRfxvLzQ6bME6IyJ
eAa7vOgV6rQH2MVHqtqcgwuW4iPAy9vsILJ/6CfEIy7OmxMI/QrhMEumCGf4cR1w
s2W9QMrlycko+mOGM/AkRLowqWMbofYWZimswDUM+L9dLA+meUqSt6kwkBFgM4cb
aAsi5kijQ9zXhaz5laoBCzf8d0DeWI9jqpCLmNAPA8b6LKjvZmhcZpI+2GEw7Xdj
DqBJvghWGczr5W2AOQArUgTwtMBdGXFi9gfkLRumcq7Cz+GjjcuHSvymlPwO/1fH
27mDBSMTd+t5YHYZji7+5QWfKBWa7KyJJQGAjfFvmU77GBrKdjJH3aBQGvy7xxLy
7OPRyFRsws3BPO+BBQA6Gv0K4TCXmjrTlsfmxS1N9WO+e8fsY0OjlJ2+0kA2RUW7
5soXUQ0y5yq/B9omR4gNksHLxAEzu9iI486e+3ohcr5+W2DBKinA8pQ3C0j8RIuo
jCZ+H8OMPIyMI3OiUXsj7d14xGcmjmuWb7gnBnBqoir0ZDzWDjbdJLxbEvwm7/6k
CXIqOebBdTgW8tF1sWd5R9YnuQI3xQmOYxOh3fysb7NCMIS42m+Q4QZ94Byin6vM
VBBHkitCUcjRN9VA3WbS3YktRRvu6zt0MuLF6kQhOGRnFhDzW9gmoGicvclOp1mm
5vYpuDmPMu8q290/IcatLzrl1vixkHg7mtLXsdNSY0spTY1YDnbdHwN3LoCjteMs
Jhgm13EBTCREdOgkiCi5Mcc7rYpWq7GH+zo+BPcT1UA2km1p13I4Q77svUWoNQqc
Ges6n6nTPKymibwCXIvPByA0aykZH/Gc3uEJysV0lAt0Mi4489G6KrMM8Sy0aAXK
xGGRTAsy00270f28AxWsNIRrbZ9+Uta3ScFdHHzglCJ2DjfXiuOisinRXbSc2bMn
O3mx6qVvVxKiz8vDOuNb0rOfcOGZ7rPYcEspt83dTfYM2wkYOMWJNN6liueO1TSV
LGoVFjT8gaxVg7xVpXjgZDE7dn19IuIe2sfEB9goijizyOqbJDGnPAWhLV49wTpd
Hv0fbRzN9KYj2lZXiUnfF85+BM232mvhZOhODuueqznNJgTUWnJY+2fNpybxgJd4
JD/WKIQ/DRW9A867MX7WqNOcX9zCBPaDEkR9a7nbiKvN2mW/QRtKg0PjNXYL2AAs
Uz3egW9llp3nCJxn6wLKlqzPtSEIk9j84nXb/7p0MZi98Kw3+88NaG8oOCUmDR3K
+0Q4QO030jZsmUblsuaGz1Wt0RWv5Eq9VzFBzHdsShQ/W6YM4wa9qApFBeHiYnjI
Ff5XsPHGwR61LP48f5m4R3UoriNaWUDPLhsGbAoAjE741LIDiqKbYGPbvCOH2Zjh
Rlub7XdTNwujuBWCoMmHpEh9vYwJd8dS7cR6LbtoYalniFmSVqXCKpgnHjbbFoOy
6YK5GVN79fiuzJavQP81tNTLrFpfqU35iY0cskmgLSFXkt99fzm0r+ofo+hoeum+
71Lby9URV6n+Wfn9FQ8te1a8alGIyTnxzoEY7duxfKhKJbVy0OAR90PiPeJ8Ius7
FplO1fDBMy1ZaK0sO87irUFpvMgeqxi+XiCw1lyVnsnRnNdbbvY+i7bgMrCY/S2R
dIogEjh25LCXokMFHxgC19gUSB9HvZkUb2BTC3p5KcOGO63ZUmMCQMmSTMD59+1h
7fszBXx71MJ1BRi0eENENTYhkczOFUHi9Fhk3YIuSaqClYapQbQesVelmrmnd0MZ
R9tiR9TOW1c3ufRmX11A0xeHcuEWSRxeHYhS9zBs0cec+Rw4O/dj9AcytyLXhHXH
Lfx39ttQN7zgRhiGd6krEFaSzc0vCVFhkhbj3x2vXRLxnWft2zMmBs0uoDAKdS/k
zguJ4mbDd5NIjmB/4x28g2WGNVjrENvT9EyT43Vvl78GDe1ypwZqIQcd+0jbOvVo
zukOFxJPsK6Tyf0zYJHWBzIkaMoweDyIZAAaDjWtTaEohBinUm/IuSCQcneEH7I+
fVJO5I4zqJw7Bs9ewIKlTUj+FeSduWKbiaE/bCz3TMcPYOXKgpvkd31l7+rS3gqr
hiJ9rZHyfPBqagf7jI1jqZckZC8BvAk2OJP5d2c4UfCjpxqBLvqLh2+LygZefgIi
9xKF8hpl4aSL5EtHhXMRQAKkyWxly8tsQmeyXHEkbcam5jWOig5ETJbc+/uNMgaC
9yXZ6z0VpPVZpnZpcc3F4VNZwXG8S6NyqXl9pmDWkGX3atWPLxmRC1Y8WnOrOVxj
gGJ0/e4CmWe0QzDzgeGBHJZd3GHzqLQnac89Pa9DbOeetUZicfRfH6AgOHcXeXQB
koUiMox/Epc6Cwxt9hHlbDAyhi9jzFrrKr4XGG0jM9uZEM6QENJAZc9S/5VOqNX0
bd63+3WNx4i+7KvWeic1U5F7HMCYqFoxfWoWtJ6qyxh2qq0bY1VGdLZz1qMGOyBx
jFEouE461sv1HMOCbQrjduPsX2G1oRm9fGNf3ba7CDkOdWPWhYx0EZktuI2WdmXD
9+TTWrjzSRXbx+b4ICrS9MztjeqZzhJ+XLF337WgRWE3jyh7uqu0z7l4t/RyUvaW
VCf/OolEjSwdgkNIV4eXTX0Z+L6U3yZ8F96XrfKO9bRKee5zzlriCBlntnHiS/s0
UdFY2wU3bvXbo6MOLNRjc8xCLmKAawxc45bdWdnePpis+nVcD6fFe9lQ6ZYlpsvg
733UCKmBWYAU3RG8PLn3s+Agyb+47nvmiKhTIs5m+pKGenXhFQ4Ce6+CUTnqxNmX
XC4SkaI/rxqHrJYto0oZBVj64dnPppTrYybrH7w0s36+p8BeHsoBPQfZxCfsH5kC
ZeCGfaoeA3OPhNB+TBCTuMIciqYsKg/yH5O5f4PcWTgr+uKO+mj7kDCHnuNTfCqx
5efd+EkQ/DzDPVYbaroIPOofvzN/3ox3KeK8fPE/lv+IcPNbBdfsTl54v1dneSTU
sJLQ73r3iiV/6yKuM8wRlsYAj9t5tZ9BxyohIaFrbGoI5IrhlkDmxTUaT0NSZFmq
y1+u6Gd0w4m+HYRF0xJYfcWXDy7tCxTrGYMPmkR+2cSRVWpe3ifbSKjCfXKNPlY/
YOfj4O3/TuJ3F/kMb0hqblfJ8uyhMTZIa/jzDdKZqQZFRFLyuyoe9bLObEaQuQoQ
Ur+xEV3UGwjSNLHNuH+F4e3kDaVU5glP3IypiSsJQZPU+WQKs0zxmLRudRiGB24Q
9H4Pt3DShAiCmmaM0CZhv1kIrgdn5HxMbvGw/ZH5LcpgRNeTiz97ExOMRo04/jui
4r1/sDy3YuvNOzd5X/I5igolB8DMTISZ9XBKaJ0tlMMxqvmwkMt4FtOfETTwn5aI
v1MNf7bgjbruk6ZEy1nEjMOjj4xsp3/ZCwa3TeC8yTJ4GwDhmGcUvaWsAWJe1ZBe
pADCxfOeNjHTD5SlTtPydy8Que24gCY3k7LfiHVFJHVQhpuuoGFAf4UK6XbiepKG
zV6u56pzmNd1EpbFw6eDLQFWBdXjeWs/jq4vIPU0Egju8KgVj1cktOtK6N9U9KHt
nuv0dQwWcWJukPGh8DVPtgd4kg7Zdt71c1tzxflR4rCJOKdhwHaZSbBxJGysRlZl
ePypSznBjQ2FbAZpDKwTs9mwyZWb3RI6Xj8vrRAO9nQq6JAFzEfKiKQN0JqSYNGq
yLmONKYFkgAFmN1fVT+34z2HiUnQQwKBBzW/vV1S2CbDc06+ilWMY+DNb1WTpEqt
G/UZHhHp2qhvqt6Pu700Rqg2RNoC/VjLUrXZ1vBTsPFwyqEIysNuscQkuIux4DHw
6dLQYkL8FiAi/PU5WRPWssKl4EiQ/f5W1590DZpLXE1PwO2skF5KQaY/mtCp3vl9
RJQPtK5TF470SYFC6Ui2g+T+hGkq3ukwrpRposQodFzZ/ja5ywtjRSLqprYks6zg
tEsQh/p1rPhah/2Branme36mBUvMzshZ8kiAXMXonNzgqh9m8jiZpw/2hXqNySVZ
K3Zx8tWoyu+nD1XPi7XAMlkuBnUER8YXa6MW+Xpx+2Ck3/L4MwzyA9KTFlgBBHxX
KjLqRSvzBkAh/5FZ/bpyoZ4nEJcPskjgzTGFN6GIJgOcG8q8cgJMIjYfBsrDOqKd
ATiKynEe89qZK1v6rk+Yipwuli8yhHPthSn2OO0RO2gKn9Jy0FMgRnfTqLuw2Yix
GgoDrhYpPRc+BS1LOrnfwNJfaqCggAj32qiorB2Sk+AQ7r4JIoQ1wc4cRu8v5lYB
GaHM8ogn8KwfK8h6soGnP3HU/pwGnKPSb7PHk2hW0ZS7pPCxBleDrH0lX3SCTm+L
czgjY+fW7BnrrsjYYhajlh4zrpn1bKQwO1aFNm0LSgNfQZ1AHTTPevGS9FEhWOAD
UcWrC8JvjWFqWqscyXiJMWb53zGBDrasdDyGhjoxpw2/qOpKIcJUmFj0SOzWCBkB
XQlK0xmDx53ML2RXSRwuy4w0ZHsL5FIeNW7lpBw0Zp0Q7iHVUoaq4/bSJEH9tsT+
s//ZncA6lukdCa5S1zKDsHIDyJQfmLI3Z9rFP5VAdPdkO0yOVVOaU0Ub3uAwTT2U
kBPkK/1OgKB09837cgXvpqoVmsUbOtFmYydXyKplR5XXdg+CCeQYqqlnjVj6eneb
AP9BxGb4Ix1ohxQUNhkvi+PTc8omeLu1rJ527moCeDwEiuL8csRNGSaLcR9Zx8TT
b1CKUrnmvo9hTKyfWSQz+Uf8qbKP5Ufd72FXwmTAtvW6w8oflynv2Hp2CfDkmxoY
1zm+ZZgXO9hjNugGTZfqEktXcEVuR7nCzB/dkeFJ7pzr8ZSNpvG5KFTAjaYgfO0c
Dql47wKyHkdJuOanB6gA5mUiu/bZPIntoxMlhwaHKkUkaoWCfAk576W3SuVqMTWp
BvvWw7pNb6E4chmE/XXfU8c/I3v4CnQ5+FZGNb6ZDqWzU5UL80iGRQIqfK+0TCaE
aU/vfEIVWRL3CQ8gMgZe/WgLGwj0bVp4bTxCKKhd5Bhi4NBQOi9lm2YyO4T6Qin/
29iENeR4Z/HvlqT6TIAIgPXMvJq2Bdd1ZmDAvDNPewX6E+OuMwhst8NKhame9Arj
2PKySZlEiCxLIKAsne72uG/8zXJvZXGqQlC1lEKUsrSjmuLqzm7jrXprKDlE8Y5g
ScfeK+dqVROrYgwywIpEkURzIH/OWdBgKoaI7Ei5K1qcFlnXDIsz4xIgnA3lfa52
0ZeSguR/uGv9lUKIT2/Ba8yhw4ydcOgKAQDUPfmhmYYVKhG2n8BbZaIz9ezPJE4S
QjApZTwKckqaHN4byqBygDv+Z5lChN+Sco346FPwqEYZDN5QGQxWf7PSh+JBbubt
WnquegDGy7gtJg2mX7UGBFjKUcxCkG5A5l8Zk+B4SjcN4HpQsrRdnKZLJOy10tbT
TdLf0Tl78vi+frFejQ6dS4570EI2ecDYacXwRPnyK+hMLAm+uDGT1C/zSiJjpD9r
K3u7kcwSk6P4nZcMQUSbSW2SBWivFbjwLr2xsSQ7su+PzgTUjYoy8V7O6RwVOLGa
CSkflGbn+W+DC0XApe71HD9ZQwPRH0vbF8PtBj74kenayAYs7N33PdpHvmBBLbV+
AuE2wWOGUsSi3Jq0MIZK+CD31WlmqYpIwKBrggSEVA1n3VohPdYmnBU6rcW0HX1o
UvFtB82/RFEU3QuxeojweCAvJtRD9AYpvSCBkKKv7WnnTDvqt5LxrtXHvTBInlNh
jmzHOl/gsWWkmjpC/tM8F1uUPYyYO4FEblqyFnA4rAGt7TlV4M3NrQb1Z41BwSbt
ABz9kAXjDylaVkq5k/7e2sQJpAeMRmzom3BzblGgdVEVrhNspv7e1LzrhwNtNyik
g4R9G+pxsYVKYvdWyQEMXNN4oM0DNB5xvNrMPAnzjuMI9SIdJoutboernoNQ1Hjd
cRRS1V8soz9D/N8JhJv5+WQeaysdQHmUurzY0EM4JNJ0nf0+4N4vK+xlCNjA9wUc
lJzPoR/h6Pnd2KuFDwbI7k2txko9pKt2kvsSsRTdcNKOnIF0LEbVU00lm7wLaPrY
qmEXBc03EcAqOkLbt9pdaqKXomeJrN26s2/NYvpNkn+osnmSjiHhWRl/dqFVEfCh
PyzRMtb3PfB8mo+S9QZvyP/snJs93MExEnfCweRHxUFoOmR0uZ2XekqhvexyOOtf
rT9jaOGM6gILZ4Jk+yzf7lkIkOUVOnAI/of2p4UY9czICigs6eqJu0aq5NOAWujz
xFjGqXs+DD8PIzFrAXS0xwO5oxoo7ZEYEw8ckhM+b5yVP/lFKq+zjc77OS1Jru3L
R6O7aQPrVAqFW+snbggcSPIngclcGrPtSFOg1atXhCNB85YucZuL+jujQKxpkIfy
FiUHbvGCIG+2zt4ZD8iNkzYce9Vrvztta2I+UlKCadXNTtJa6uYSCaUOt55KVImM
fcSCKgcnrYHH3mVIHOqC+5xmwG5/WSHu6uuNgepD3f7kqMe5oBXQ8QstGSIl8aZl
vxSKxUVPG+u32bxODjM8EzqmMRQaEKd/ZABPzjkbJsbHjuG4evdbMmZCM6PtbfcE
wdUpaoElqBO6pshAY+xam4LCo3XoeOhcp69X/SXmBueU4Dr0GvgMTuSQqSf56l68
oo8fvyQXr3Rn/HXxx+vB4GtH3jixtroUAN5yP9FHYJAulraLyyJuexLnblUDO4gN
NqOeiy+REOQWXwH5VTOja8mCdY8IvcpmW9JxFu/85fvvOcD7LlmyJEG8kd13GhVd
gqlTFwgBM6GZc2wmOZBrCZzHGZeDGnc4e1dhfEuUdY73jN05XeFzGgvJkCF0KfFW
2av2Cw2qUksHNKcr98RZNsqYaOXkhbBN6zo8+UwdJ9IqsnbUF+XxewNmngsd+GW4
kytjWzcHhmEX+17H4caZ1uhPaDq4JLn10XBXMKiyfYMzhWQaRhXkwUM3+Zn3CRkF
3l5GQY5tNkDZeTBZS3Up1g34Tp8Jis7Y8rExxwSKrVQaePiQ0AzQ7tkAvpUFli0g
0XruBO992eN/y0bA3bRshn+dOoq+q9fl2UFjs07IvWsk/lmfFyyMa6TO++Al92at
iJrtBklVcRopWvvcNu1KFqfjsaZIEAW3TYpMz8eEom/CNrK9AqqyHl2KvucUrBAb
1STwBw8x3ZttI5B9kT4wbAd36wPr2/68sZOgFzadSSk3HCzcXkgPNPZNrN1w65UO
KRbFnnwBGxqxJ11ejZwfT6cfoJyQT1J3GD5G3LYsgcFMRHm5pN8AqKKWa2Pv0c6v
GT/VURHj/RVKw0j+Xd8ld/X/MC5ojAg3gwv2dR1e1hFaYAqFdByBii8myy/q/RCR
De9EMQBQIlL8TKDIl/9xU3VCYD9qru/pKhtbLONvCYOk8CSMq3QAmswn7Qsu7cQ6
nYNGfDmyRiWmgYr7A+l5dyZ9W2bsrAc9hIXj09njxBHfqx9LKWcygDonD99HbTMx
pXRZ2rmORWY23mSa/aPByZldO9bc8e0ZOqAXfOUTkv977xFptjxrmpTCF925rsy0
ZqYhAKAjKSlssL5PGQtmUS5R3VPnBzcNFVHBCllYFmPWcp46MsF/N37n5ladVy53
OxN66j6wboNFh2r2LSCRSYGuxQD5d73TZMt83PeLRyCYL10sVNaQLvGdc6KdQJsg
BjGOAyfNCke9nZzKESqx094abSkEJ+gj9hCdnslV6UGk5kuYC4azoPM4WjJ+7IYb
bEmkRVSzMgMOxBG7CuRAXL4IJ0+H8XDXMiOvsPdAMTSB04yjuiSduppwjUp4KN2Y
3jORB7mrYVhD9Z4WmKT/vsGj0QK0VY8B0zoGsbis1gHA4h/H09kHvoIb0ebVMX+g
Vwc53BHVr9RMRWf2arzvT8Os4450y6y3Q3Mn695cKwD2C+QeTtLzlAtYoEF/b6Og
a0nFZ9DnP4vBnt1zOmPy1kIMBu7p8lJgfoGSus15oJPlMn66CEMun+OBtdPR8BmZ
pcNGo5e8ZBopOPwCDwc7Uqvp2HVX4z+Ah5owzwyAaja//WSYYWZL33vbH4ifNIuW
OPik0fYg9PWQyPRxLBeRVF3KatIkPw6+KSiVw0X7Bl1+KXwVFRzIiQBMltE0TGym
x7yNXs+OCkaajHcjqDqlopSwJpxHbdM42o52H4OUFnNg6edLnddKHYexwPvsq5PH
MsAOSjnVmEgJjCOCuMyRHeQWQbymEVNbue24rM1aHhXPEOSldZm1e8LEtV+UapJh
v9iF5YAM1Vh+x7dU7Tlg0qz+4VR8JtqENyR49+AG2stvyWGNhJF9W8UUJwt1A0nI
5KVY/hk3a6JoKbtmNG89RzOadqJ8QWAvkVmsd+F2e1phVDLAkMx4/8ke1DXze81K
ehzrGbZkRPcSgq1IrF2hv6/MGPtj7jns00fn34tS1MFEXtD6qpDF6OXp1qF8/tiL
+A0I9tcQG/X5YwKKJzs/JaqtQclVoVxIbXPDGiEye9Yrk+IGn2crcoyHHdklZ54y
KdslJDFnPa5QaW8h1/W8RoTq/fU6ivN98eiOlwTmE8Cz6qlnP4F7HGiJPQoo8m/i
baftp7g5oyZixusnPXT0sXWow7QN30y7FWoRQCBkAYOqwIDyGxlCJMousTW0Ma14
Ig09hs8nO/jhnhKIlV8s6TntAqjquF8FgKIXZxSgu6vMEI1qlMbJxplLo+ob+jhw
Zx6TPIrWZ8MWbCd9xT36xlLDJAlwTFpdfEiDLyAJD8XTbsVXP0kVopTcbU+yzslm
8D2aRQdZBYRbLv6uEH+Nwf+2pbGj4Q4nCfoKlBN5RN3lQs7Z8bEYgi7i/aXxyn97
MVb5OQj3vrUkMjQtfcb8a8Z6e8zsNqquAOKestz79xLY3cQD26DYqXKN7yzzkWCm
h5zkVRQUct8T+SPaE/+SOGRzgZRY1FJ6FZpB2if3LEAJqfJxIXG0ommN9/mZZCno
/byNz8vM1LDBzQouDqC5M2OiKHD//u3Mm3F4Km0ENpoV2XTMuJ8yoMcb8liGVIl/
x266KmfDlPoXP06ZbZP8o1xj5fBf9pIQVxXvKKdbgDdSYcP2qF+ijrUn9n7BeFed
cFMzORyq4qkhRVov5CKsFQxOuR9O/NTu8FgQ+dnNvEkV98VvDG8yBJGrgKxT3aWW
Kg0Mm0JcqGxeyipLygSn775UUjAqkLvsoIlXxf6phsHXlbp644Svgsl/zGrDgNnk
9K/VexquE9FpITUbDrrnCkbkdf61fIb9LA8AIgnFlPRzikKGXL/Ha/Z5jJfLU7U1
sSJpYMx++uLJCYThPqP2Rv1OXbhF11SG/ICi+wGhuKKlVJSX/TuaWhdGZ+3JOrlr
c7k5BGHjFLAvMro+rxlj4XMc/5ZOQF1z6ipGP7iHbPkFeHA8zBKjEldXQf/1GvW7
CtJDPKp19UmARaReqPFumheYOvfvjdxD5sLIMVHGKHL69Vh9jC9V2o3nvjpm5piC
dnnkTrystwehIGVIGn4d74dkaNzgucwFYo3aTWGLPr0fff8CtLctjDfYv16lnanC
SpPxP0YdW/OTsJq3SKNt11IkBRqTWoADB1FB6mC8wzHhuf2WL65J0mqn2gepDQSN
SC/J/mbAAliu+7loQ6AGGJn9IJGMXHYaB7Jsj8t1zz2JQ/V8pjbHtelTkOHXsh5e
W3KWdrl5fOXl141Cxwyyu9uD3RCBmzJxhyGp8UkdA3tO+Nv+/SwjKRlrkc3NNVny
vnttap18+rSC1XF+oRvmpmSWSHYIHY5vqqnHy/DgFhpZ0WJ9QjtJJNGEaIrWU2mZ
j2ohvU3vysgc45N6mfdkpKaMxDM1Tt80ULU6N/eVQ04am0hLQGyyZt9NiRRSI8g9
I64MTyXAss2bsyb4K2kcIaSxtEjAMenIDQ+3nYPfS1aoZunXk6Xs/xL3V1yK0QOV
aYtLZbYs6VXeZm7SKqcIa+GhXFIEKwdqpm42rcJSxc16ZKI3UvnTZcNYUnLYhsD/
0xlqZv38h2afixJFRDMQ/7+NGG/skqgnV3O8kbRjHz4gFZAa0J8/5mK2NayzyVVK
/FeWqLbJVvX87NT5IVB3aIuQ1fSRZvQvXW4EGXjnrP8M7DFFos8wKrtqdTPyopJR
W+SDoLv5xPHHfTbAfp4c/iXdOsjInmyf1rXIEGcuWtRZIpFXguXJP4RwK47JZG9B
TgnFcOY799HMQC7cRnPNbQ6oQHajWavpSmpMh5XOxKcE/wkHlXnhix3U8zXHrQ//
n2/d2fSRUHgUSTQTu2+/jjYA9L/zIgJzoOq4EC3ydFY5lRpSG6pp+KgfRnNONwxm
gt2Cbwb54NKbnz7PEl5xNv0E+lXg4ShEtcBv7TYYn8Tq3GodWytzDSXfgjqj4Dve
vUvIn5V3WSvZ6rAemWW1UdYGiTBQxY8k08UC4gRD57DlFvz5hp+9atK/sppgU6rb
6KOqQH1VzOMy4UqKBDtFWiSE5aRK0srQxNpvt9HxLEcsShhTczyEUE/Ct+Lkc2wD
d7GMzFDgOptCVoML2eTArA7Xs7F1H7/NbkEKThKX6jHqjBampCNh47dSFq1UYmia
T6S0zVh1XxmVVNBBeHJDOwVEeLdtSxSmRXh3UXHcbjBL7N6W0B61+LZz3o8vc4iT
u+7AuPYSbQy48glD6jsL14l70hZY0Pm8l7TfT1ISf05aXJ7VlvjCaACmPjNgPtKD
YXB0LrnRuCi5maBDSgSxT0qXCcf+MW0dYLa3LJZvwf1L4vXCHZSepchbIZn0eXJX
s8MymTsRrGczQLKnyZE12u6iz7X5qoVqMKGl8Xi58oBkzDPTHZbcRhp3RTpI4l0y
J/OnFJ3GnXOncb0+69G5yPSNA9OClgumD2j2IcsjyehLDSbDdv13D1Not7lg+5ga
cuMIqkfSeilzTnP8Z8vbOfj4rPYPTdQOpZsw/2G99ttvIRxh8UPYMHZV+N+dmKHH
4FaB4V7YaSs22UrrmmVJ5/tq1MktUq+EnWdY7CegtIyLyL+BO+ZrJAMDZ2mpjpwG
7vMLSxQ1DLYHjHDbsNJu/yoy5UNwcJcPbgcmLbICma95kN3ypuM4lJpB8k1yIXOV
1+najCHzMswJ19PfWQNVw8swGbq6ft7/b5h1FeHA82MMEEeb7j5zBAqtD/29GmVV
RAaXfOvKewkr1XYlqdwMaDUrpVfO7jjWYFmXW3Myj3UAY7FkgDtptLlA35tUy7E3
kCOzA2nYEq26ckgSDGNOpfSvEq5YnIqVI97EJz9LBL0/N2yygWUcoHh5vCsfc8iL
kfgtTMr/5/D27z/S12XfN3meV66iRq9UE/H6M7d5392Fz2xx4SYFIYI5XiudPEEy
wtdK7L2W0C5HsXV9Z8I5GYYDHaB8rz7nK+vu64XEyKztekBGLTO7UaaQUNuRSFlw
Xt8aYvaz5ZvteSzMoe8PRMTABWmGz5Gb9EvSv7RjYGtV7yialUGX8V59pJwo+x4J
hHwCYLc2iBaDhAHcDA4BqGHdRSXoR8rkqKipg6PuB5pJ96MrJ51Wo4b4WdPfEg0e
oYGcvKvgiCgmnbRfgJFB3kyWuFZS8rCQo1LnN2GRLq2LEfiw8eMj79btC2+Wrd1J
KTUZTpO6jzg0vnr/Z6TJA8qFY0nIzzTtdEcwc1GXUS2NkiiblRM3hAsCTFe6r18q
SafU9FOMga2IAzcRUphQoz6owbQPUhlYiM5ayclmOYWMSP32H1pzegwiM3/PP9h/
86qk/s2dfyKMIWhjognOl+cAPCJ/JSCO6IqBFs0xmTiMLbdEIEWV7vnJbhhLONLx
wJ3DSgRkiqrwFvZ+qFYJzWDjRym1jpN6zpK5zUxTnHgOs66zSNxR/gPEEN5ENhBb
yDwqDzjJ+XVS4RfueLCB/0GSYceAIux3Yh+RS8+iG/thUqi4B/DMnaePS8gAToiR
X7NubR3nWxmSy4JuJKEbYCi5bT+V/ZlRWxHIXNuXoBZ838VwYo7m5Wve9RpounmT
XAcc2p+r4ME8NNCa6Bskfj7XZVjE156MgZYGdOONFr2oPGhAwPBYonLpoVFhfKNx
SpZqWYpxLCNQVnz4pMzL0AjpGmQ+e/MRsSvYpXcmP5rAEjz4rE/fnwVVrnBqSVnX
ZfqN/jV1/7z4qch+XO95OjS++PAy/WUlUwrtgCmf0EOOg4DzZPJKXWDk7aUt0QOL
acsn+kthgc7HuRo2Sn5PJi2YVbY/Db0oelo6RTVi8wbwTpijI6gdLoEqDBzf3hRc
RXluQnfND70Q5vu+G0v10hB/YoKTt7mg8ttr9hENzKjKmicfwI4MzbF9ZZHADWWD
7gx026ZPHdOIr4IWm5wGX3inbR3orczF7nUfxL/a7iXAxfg0tM7g98OAd0fgxHHD
o0ow5z5fghtASDgFFUd0Kz6oa6ObwqDwqLItncfzDNZ3z/OnZDKsY94hWDWjaaTB
hZC2Ulv/Hlw8TUuhrnL3YR5kPpxUj7jMWBmSLDwnhM6FYV8YQdwzTTHKNHYoFS+t
EtjubBhnzgixeCehQZ8Ad5msPBFroFvN9j/21m8Mbj3wTLQWyH8DsvHtidFtTVZo
greG3rGD94/wxCfpfP+DpDGaNGZ/PppySFiXXgiI/w55lMCHsmy8+t67STiKfa2r
5WbOUZWhqloxVwGRa5x2wNpUxbdgap/ewno/OwMX79LYTAu8+lVt0fk/wJomR2xj
KFvfKer/Fnbkuuz2OCS5AGRPWagMNXCSPTxS1aXKDZkEy8k9n3e3JzBszyUscdUl
u6Z7PCL9FAXUoRzbwSBGPHZqYYArWJlGzzx+I/f3xQdr3WxK2/h9lyEoeR97OG0S
/V+C+izHcTWQ/bKxFUS7vbfGPfVj+vUqQUX8f1u81Nyh3PCtB9pkIe/kMa+TlsRO
HXveLQY+oOhFIQd54FyXpO8r2H59m2g7coej4zFeBmNVDg1OG/8SK4V6qqmxOj1X
o4KGt8wNFLzulfIkbgDpJ4zqr+B//DfdOFHIo7owNmngdJeDsSmNT3hFSJuKSf6Z
D8dyGYFGRYjEw068HTmVVnHiy3AbO/1TFXkPLGOqhIkwqpZSWlkFqQAszb3jFasH
nNp0BBaW9js7XltX3Kb79xRLBftc4AJOFFDPMkhGIz9ScNwkLzJEwzGQxAqytSIA
dZubqBtNffAXY/UgZez6iofjEYWe3d3lukInewBcQ7F0TPGOxe8hK+QymdUSUkXr
WmLUEQNMnH8yCvrTjQ4VBGiZ8YWDyXU1B5Svl7zQMQOc/Vf4r+BDMtOOUu2SCxEj
xcwfzlkgc3hKmsH1UMGnEo23KjZK3TWBD/gJkBjTy7lamiwzVoLyBygCHkTJYgmp
Hvq1BUGyuk4tAhmJjkMemWmVjqwh08v/TyIojwATAILKJhHI9OMLJaCX9wkDjkhI
y2SJXZ7WqXZIqyLNm/FTXzwu4q179mE0gLAARfxqpYIxrpKBac77jVmMIcTIxftK
uMpI9VmJLI6LMt/HcZN9aDgKuyjtSTTvzLbyzrxr12gSc3Yozk63jcA6ZIjhs7hN
ND9szu/KqAsqLACQcMw+iSr1QOzWnUUPVfRYVJql9Vw7cChirO/nglNhSPdzuo/f
4r8BLAmV/lqqv9ACWnRElFj9GQxH3KHgNtU8VSR2zlD3bYfcnB3Rip+BTxCVcFVk
yAEHj89lRNOL106I9b/vJsrv6FSR/OXG1l9kItCeo3LE72DneXtveEP8BhabEUTT
0tt/9zkHkiGvySMamLGQj/4InEvn4ZWTGxskE6idgK8rjYH8ilORSCZVcru2BG08
qGPEkuvyningQ2kl96XW+Cyi3qy0kYokmezI76F+kUo3fSc0xwk0Ou7Dm7LM9FDh
7wG4AfMBvK+hfRjSoj7U0GkfgvNTiYNplz/gwMRx3BMy1EhVPPkSDDYkS8IYIl+L
DWLrKZFiHBPj4GTfkVTzMZgswbXY/kasMSbkFKTK3hyX6TblOq8XzcncZJY43aV1
Eo7MGtogL5twNluNRLs3dYWeutqr3SyrJF2mLIhqSayDmhF1fTep8QpZee1kgln9
2n+wMjJTN/t0B/oV3hgPJb4+G2AhNNgF5HV4cKKrxHle3GrIXWCDRukcs//GzxQ0
KwpPHL2C9lP/e1misxNaQXCehhvEGVBSute7Fw2twJpnL05iBxpWxewmQ3qx7wiY
Leiap3Hle3WrqouGBhPsqEtCnqGmI+Z7VHO9hfI9Etp+NMvEV9w4Sj1L63OkwZj+
nFqj04rff42G+MO2rM16Z4mQX4dUW1O3D/HypDCTNwf+zPOxKLIqSFZRFiE0h4xs
I7bG1zwyxRtQZ3w6e8qNIbsM9gauHcQKw4XqbFeBTnDMxnMku7PBQmHY74dsJON3
C9CV9Xe/3HXphKJbjEQgH89KAZhVL1eJkDeCsOy6TQbYPyMUWbAR/ZS4jdlq0SPK
rvE7Y3ge06Op/aTLnbudUFw/P2UKLA+fAucL8a6viZ1WduCdXkFH5me/moO9eHU5
JKIrOTZ0OrxaO/Am/reyUqvWsgmVfkGLF9pFGLEkxnRH6T+carIoeRuSUkKy3mDk
+mGBqEc1NUj9iMt7cH7XFTJWXER6R1JF8hVMd3v26/XK2Ldyip0OxgIVhgOuYS6U
+nrBBZGneSruGXNt7QJ8NJYB71awPkQiVds9yVNKcY98cUr+QYS8RB5oNnvYgC7l
HF3InfhSCn31RZuzVSNaMJw7skv2C/CNBBDMnfpaILcLMLSwnLiqUiYovaRgioxW
4UNWIer/qpodPt88P86X3e26K1YxAfJ8YRra+WkWORYwqcy3+4TTmVEbvC3CHi9p
w3U6LWIO/CADCqvWK9FNvBWqwT7atoej43FYuoxUSs9Jaoih3J6CsQqWsL6eb4TB
4viAqd/O7u3aFljTNsysHxtsZk1ct+WxgnTtH4gcmTJD5iqUFY1RwO49XqkzOnpp
pxzQ9zK3b9BYc/M1ueaMYgGOfx8eTARMbViZKrMjYAO0LpqJcs+ookHu1EIZu0Oi
fnxX9jyErI/jWWvpuwfTrCol0oGgh5rb4qAr8T1kDmhNPPLHrELKjQH/zpLSMcJT
1HOAlALyExWL2vW3s9Xbm1Dg9BOTqR5/dftAu09vH32sJRj+2WNcZLtVa5Vuwqv5
qXO0zQyHnBEFFCUtiEOn2tuof3h5TKP389urH+fEro43aoZNOQURjUoPtSkcN69C
GSWYH/SOwowUGDPOEhqE2bI0p+POr0M5wIGb8bMp5adHa3Hd8BdVOrUR8mPOcyek
/gYVDacJGF5PKy+bPCAzw/gnF7/5KjvVqc33nU8JvUTDlxDqOqNQh+PvsaEvcvc5
f9t13aSxMhi2iRLy7MQnkALcsryGHRDmJcUOIzkehVuot/kDe6r7mOgbiC2cwNPy
odYEiNVTmOimcQwfr9k2PdSCpqxmxX1+pNU2qBxvQuyQTkENL4IdgFjBHVgbgRDG
b50jkJ25uJTbt+EAAeCrK9FS3BpiV4GEx97CD9kLzwKbPDEXD9pGhDrHeYxKlDyP
7IfEmlzFQWzZTVMCbJpqd8Fs/mRPS5nUchRxutntB/WJoMWIKCg2TDpo4MhM3T6w
R8kalKwRtXbfSMMmBXBPB5uVM2mIUyG4ZVAnYF5VliLOX5/OzElTX6w5QGxj0uAP
ScyuAWNdz8fIWoSb/hSzyaqRLwop3GXi1F7Fv8t56Fv0d+bbQrRNq4lGxam+WKWC
GgiFNQkyzDUzLzz6cevGDXc3niJGB2fHREG0dFzy9cbblAUR/ac56kf6rXtJfS5/
jlrju6jijCYK3eKU8Agm4t6Cap+nvqg8L14UqjzJ/FjtmZyJUCcY+KQscXz45zdI
XcSOyycru7loMNhDQhK2HVHDQGYKFo7C4gitKN3mIIvmuCVVxvw4+nTJuPxoR2Tf
F0Dg+VboK7+byMVt0bqMRjXf60VicHLf57Tu9Tg7sc3sn9C+3ANfD0B76PWIEQTW
0ixvnBNYOkkaMYcc5hao/jSXa6PmJmCEPQ7u5J91hhbB6Cy/DWUVq/KVlAgEFEru
A3z8xC/+uqrS4GfOA3BNqPWwVnJLNdbkmlnlOhKP3W8yJUFi5NODvs0XhJFEFVH8
HQctXrA9tNwYNwAXP/QptcNDKSCS4HLfkxZBoPHnQSTr0D2GeBOQkq9t60HJcHog
V+eDt/gRTa1Jo8KCil64Ml90TvrGrkB2rk7DWVXxXMeyhvZz9hTEQjN6MGMcQEi0
eKujCxA5m4dY9v58uldXrxcXvqpnqiywOwb1al+hFPuZfe5hzaXi4bYtDfDOyHqe
4aMggWcPIifQ5dc9rxg1/OYoda16zwZ1gE4Pf9M98fxy4Ww52eJWdPDf7yU3jy1T
yrbrcgcXDhY5Z6OOlkh8gADDHuZF0EBXXXozXyAxN5dZ/vh4xm6iTHaUAOk9jS/i
zCEddiCeAFlNd8e4+ZFYRs7eR9WgVPIgucLduXzLVo+UOypPGddMhjAZRMXrFD2V
ctyI5MsEdMd85HwzM2buSXHupuqCXiiqmH3zunHS62EdXR8VxaxJyJDBgC5bzfN+
ZdQbhJw5/kioPh870Y9hdVQZKcL85vuko1Ixcul8r3ftMgpuzqmtDwnU8typcTHU
Y3m04gsf+3yBBfKVbH0TATxwqYI6HXOM1KzLszeDC1hJkvwiDtv2jGjL2kcw6Zaw
zAKtNuDUmvDh/zB/6duMqlp2KDFZrRGvOh6ItEorKgGwNH0L4Y9sqBs3x2pmO8Vf
xKatOC0cqisTcPaNmdIOaBCQiX0T6x0imV8GUCwv2FpttTaU3HSr8cLZcLJGo2mT
9aqt4OOz4oHUKDKoPstUpnTgpf2bobmn74Mpkmxg1qk2HII+kXpBoks8l9hKQHO4
+xpvNR0lpRfkVO8vQH4aLUJI7IPNi4ZnLiUFO6H31uY5oE2rnM/rimqhYvmHzEa8
+FqIHd3dJ0HY7Gm7+bxv7IdlXR7OE0f+Pc29/1QblFxF8C9BwFJAQoOT+Wzl5it7
3G2CEZCbh4gsWbSFaqguvwvSbJsq4rCZgsPwkyeGlKtOl+eT8wJtRjiDv2SSJh89
3FKIY/I1uXgm/VatMCDq7ivLl/RH0oC/kZZvC7E1xRk+ubS/RLXbtS+rIYQVmgis
0nJSNjr0URZaOsWhJ+JRKGPT/oX4XicPendtagTMG1hvf3mKHb5hZGaBKapnKlvF
k0rblzVtzjQflU0HR7Jzo9IGQpAU53mn5nY4bnos5mTbmqWQnwR9xflB2Gda5YuK
0qedSWoSfyx5wIsv/BjBy3Qul1IIW7lX2u95ZOlxW8TzNacMUA+2+1/st1zcxGe/
IUPHWDD2xNUOI+o91wRiXejhSa8diDzQGUNMsGFg7C7OoxM7//EzWhFzHW5WtXkp
FUwQ3qE7yYP+gV2jbScEiRosekq3nRbte5vZFBT6LLzPgZjw3+A/hj56zMF4ozzV
Y375pOUA6xO0iOEQ5PKeZKAc02l4D0wYvacwdODE/BVaC3d6kZsYxp7BiYWi9wYj
/dJF7rl99R6vOSFDpNy2eTfoRY1FFvjWzareqXJu/yC8kJAIiOJsdsid8b2nX20A
v7gSKlvvR4JhvYUFQ/9tk/HDIrvtA7PuDuvZNacBduKyV/uIP2hM1BYU/jUPVnd7
1k0k2P+HxJRa/m692TIyTk7U61eeQKimKsZaBaD5+Tk4hFuwgfiQ/W9q7zszp2uU
so21QaTMgebFjGMn45ZBhw13XWRTO2t7ioC5FE4G8mOLxzjpIo19ZFSTMuXfB3zp
+rXIF2wzXGQzBCis6/f78AT678nhs9uDlU1ZBbe8diEkRyXopNwgkpEPxHvWGd8v
RecaUjiKSDtztXeRWzzc7K/zHoohsvUszmdJsviIirAHKDgyHqx9Oq83lTm6qnP/
cbPNFRYWXq0OfUmb7fN7QNEnstV14KJl1LsJvkNVJ+AjeTZ+GUu222TFwGH24nYF
Bi6Oejt0LoLi9PKYa2OgDT/9KpzSF2DuO4CIrLf5lCnCbUPtE/VzD/QD4PDZRldG
4ck8CPtIzUOBNOKKam7PS8Y6Y7RV7l3MPIgJMm9r8pyJA6gMylRe2RkonXWhpLAQ
FzX+iBHTTvvrK256WI1mei/H1Hygn2sWfzWIc1jGbE2t0VWbDCaFgWZaQoqGt1Vw
posmfZPT8zW9GBUZjlEaFeyvd66Aea3osoxDJMh5fdx/9i2EwdYqDARzJC+33HZ8
QEluHQDxiT8+Jxf3085pFRVf/8XE4fP69baQgArS+E4eDY9SevYHhcMVz2V6HLKU
/WPzwtfhHS4CUG8B83dCV/lGbZvOPkI9iqkfU5Ytz4n65F+c5yBky/MygZv4FLSx
xmf7s7F58ll0Nvj6asJRkZvUOjWkqqIYLqFwsUom7mrzAkBm3YdZptzscNlPPhwZ
VTjco6/5iNcN5r2dpDutooOZFz3YSXSybu5CwWQot6HPgSrY1s46YrJY377SCr1S
oCDg0d38gwngEgwBheBwhQdVz650Re9BmJeUaEHLhccR9wS3k/p0tdSz5lnQnCqe
86PkWZY+e/veQHBlaRSRybd/YPAuLmJ5cQ9LsyUCpXBNpd5vBgLUamlJdR6N/9Ro
7ACdT/+QcE7H2Q9c1xnMJ3EWPoUwO0VM7oZQVjflO7bhfFYbTJWWIPGHMjXerWG0
utdBUrz+6Q82caIb/SpY1bOas8RuO4CBZqv6+ww1K9eErDtJkrIpXX1OqNy20btU
c2CYZYt7NwjeDjtZShgiC6zZAWxf8SV+GAf/kIld0DwJ2dkRhg4qbiJWNH2X1n+7
UrqZUb6Cv+/rLZSSGoiOHBatM26HjHlI6CpEtSOgRk3wDE5ha6Ujh1Ohknqb4T7n
LcbNL6OwJqEDQx51aRGajzWb4IPBTm+jCHZHzokHPE/4duhXGTb1QJxicR+11sP2
Hsml6rzDRrzYaB+mM1UzCP25DP8VZVW4pGOF8wWtKVjpyboNlcEAAIWVkP9ZrjHv
xppFW3iR17Q1WLNRwpEfErLh+ge+heh5gzV92m7+I789NSzcgPfrR0UTRSYe+yEc
5bPFi36BvSn45qnYnHhTDtSgKSCT9kKHyC0ZS0bcqfIZq67zUcXl0EkUOYu4e9v3
f29iBxsr8JHdInzsj1BP9sM8P0vpYWR9T4NySsdUszqOHJxj6inKnCrX1t+RAI9N
fxTDqMjBVVnpQSsYJeKW0AqKKqF+Vk36vAFnC4PqQSpHofnHcfXnAhOqoPWZWC0D
iZGaV2+9jdkkayxbRnTpFjuRX2BqS9ZPv2t3Xk4IRYhfvfbfQGugmRG8XotIPTDt
j5Ciao4rTJMKWegiZWIuO0jJAyEa3526IjC/4FohbAxeLgu/w3OUaxh+MG0Kcgqk
JAkPZKlJ96VcuHjsp2YIaYL64DEx+Hk5Ib5+g8G9Q00g3zTLxCoFRzBeTsn3hlU2
lylFAKCbmNwcRy0V0eZam5ZkxEzHZPJLNEhi3m2MyNEstHMYDfbQ+ZI/K65aMMsX
JU5EHNChlzA061v1gIx/b7sKYJ2z5HHLRZoIEahQRurMOnZOvzrJ7qZ1DagFlKNl
YOPCkrXwTG/7NAmYzkEXGvsxU+L49q1Gq4qSrh//uJqdV+SxRI8C+Yzbs0PaoI5P
xcyya8vBfJprQi4wSCzyfZmuemLz5jP3eY5Q2jD/uwn3TyXahX7FbilhY5rUKpRA
gstdRe/TXDEfmv4ftzLoVNIDjgcv/nfRY7mdmf1LMdc0BMX2Dkybfye9CT2OEPEk
LAm9Wz+cHpQrKkywfGhiXcH+e6o5nMus5qPKvvUbl0/sXxZfg9c77x/JQMoFmFp6
teYmHIVX9OwQDZVZscx5NgL0rqd/kTfWUYrUBiooBt984/NpvO1gNKxEYazoMbOX
gadW0fpssmNuqpkS3emckvLSDPZNcMEMwDAvDN6HgBikdh6jGxvE8ski5/mGJhhv
Ls68nbn82kb+Xh3ziSMk/JklN/u6hJ7mYjE9QeKx0dk4kWcdLegWcXNAMuXpShSG
3KVfTeVUlE5g3DJ3e81LCW8ifGVBrJVYGL17v7zB+riSSWI0jImWrWobx7FSnnyG
9FaxP6mvWqLGoGVUGHWdrL9YOrpayRmYJpfl5n8STLESVmw1/0cne7P+JFS2+eL3
jBQFwNAaLYTDkjIvLJY2mWwhKeiHrNpxIfJWxMYEAcguK9drKVpX+3l5fiFRTog7
Y5vkkuJk5lc0/RF7hz+1TAOwyYNFOxFWILHayeUhIBlnMyy9jQuPb7MNia7SxUI/
IZK9JI+ofdaSPuO3HrN0xj+nCVbyBv7JrtjjRN/d0vbLwTld7pMCskzuOkYe1poU
p3F9zaR5viNATYIS8QHcII9u/p3nmg/2sttJMVJ5xGxa54KOdgPMukehQCmxKloH
aYeiCcZrZ8u7lMG03XNy9nm5DGC3RRb8WlIwBuo8DETzZ/HvfmDL7GJh2h97GDUD
6ayh7CgodQ2DqnTZ7ip7JofU41onJRValLmGnF4y1+p5UBAGOtCIvFu/YblvMjgR
7A7Ekgr/Y04WoGYxBHzvOBDpLgr7ImWZJOEMYlWI322sIIoxJRmXEfFRy/1WJEs9
HJutAc0mbT5cEzyzSOLL2TB4hNriUTnPK/QdZNvyldHE7GX1DCJaszdadcKsPrPi
gOEiwNKl0bKka2kw03uWoKpubVFNoZp/fGhvzJzlhMoAKl2p8eigLHRsLWSYva8c
6Qw6tBc2LIEPb186msDqT5X0D9ZtEn8qdgFNSO6PHSa3b1izJ8PGFHaJbOSBiJTq
6GnuDF2qoVrm0/18WkJEP49fwOLIVu4RJlyLuOTIGRrNXDB0kXGMxrvZ4fbmc6el
bE9Eatb0/QTytaQ8B8e2iYva7SzmQyhP5E60HhmmW6L3cTeGLtXl5y7P40HYpS3D
QYQj0/xEMOlIvtHlzOD3fJ1WrMh5G3v0/LA94IjECA4eisBmAPo5kDI4Y1zRRpV/
ZCo309/3xLidXEIvOz/QxtwlEPiHkxt+FkPCdvVnkr9pKl6zKTo+BfvHq9NASekq
0Ljeso1vjkXHioQIyT2yTiMJSXf7qSLgZQWeVosTHMx4wXs0tAah2SomLrk0pEmb
Qdh/se6vnRJRB0Jj2ZfGRNyVqopXoC3L5ObyP1ROGFsEGoBt/kfbgyIHCN02nd8z
8+//TKjxSVE08f4aEAkhsiqesdf1Q+QE93eRrldc6mC1czKXzH2EoFXKiCjN/vxh
wsgm98IYPYr7H6MX0QZKBzYVLG1VdMzFM5I4tvSIKZv5bOKxJQtR02xMMr/YbU8a
YunO8k4BiM8Z1U/rRb0F34qHcyVS6Pbqrrt4xeA/9/BVZzssEGgtF2209yT7ljgb
Ck5ddAfApRbwUBVFa4r3TjmzQb/mdm4QNVnla6d2bFHH3BMDovIdqjlIFneSJ28x
tlVqSH9zhy1HpFx1K940hom0hLl3kz3IoxEGv8mNaDOnMIjWxhc+6hio+WOl+MZI
lzXmU7l6krW1a8oPZ5tr/kV4TBuDiSt9cts9Jbbecd+KtbT2pUQgRV6sDtLpCcUd
ICAfhDdEgKGrREHq/NmaiU3cy27owosioDwNWR8XRVyJestMgRB24DyjCPu7IZYe
kAzezBJxYeujXbhEa8jMEF9ysR0aqqx5/6zwBwn6C5p+n5pjfBP/LgEGNLUy8wKI
Eq7YKRBgPMC9Mz3qg7dZ7C1e0HWswJPaHAxJcN3rfobDqF72jI8CxuVlvzc46FYt
g6rRmCTZhtPG5ATjPIpOlWsUlDc6QRaUt9PRbssDtTic3Iov4ezYXotstrYspjdZ
/o0ynoWbq0/gQUIRURhebNzRl+AuXW5JCwRv3j1gp6UKzlRQe1hDj21T7CujVyXX
1FMmQSS87QekFKkhVhhfCSUSIUJrDBPk1ToYC9h0aEnV/+rDeI6X7bde6RjnmVa8
v6OjFMkos8R34XaeBMrGQZ0LALDji3tkXn41NXz1+6BUZkbMKdKNzQxttcq9FJ03
svJsaRyHKk3dgsasYvpfOOxIVSBjdHrNIsDLa4kzzs74Ynn0Ykv53/U2Wb5hwpMb
P2KkeZSzFBIz1VHritVsP1fNR5z424aPOkwrzpyRIEK4fAvCx3hatKhyriZRJ7B4
k8bYp10by6F7RyVD9b68NxZaZjb5nOz+GpQJOHnLJSR2EncIGMm21Tnifl8oztBY
rTOQ/QT3pnucgQFSGrORcIQ3BDb1QMGquRGz9Zzt1g60ETiT0XOf4ywifMl0oPYL
o2scc87eFYI3OE1NJ/mCAnEbMGOfMhGPj4TjxfvM4WDWoLXKjKZnoAv/7gB1XSUs
yBVHgJIJg0Fomqd8sV5MAZxxiG3KrKqv0OohTG3e9s0Y5bnEZGZQawK0uDl/Vd1l
+8JkfH09lFz2OXC6e4V58s0NFbs3+B0qpZoVWc9UfI0WsbZGkilhLJfhfkQD+dHL
RMFBYxU5XOC3xj+JYP+fmfy4sgmr+8TAwLpDNNfI9yGawNXpJofgYsrj4Mq/pFh1
7LHNWo9ENvWI0FmzxHLLtWjzGdVd7XFcRUOKDS0I4tZ23KOmoNV6gxqIDmcuTZlM
h6eU+LSL0bXY4r7Lz7ThJW7vcWyZ/snZNA2rMjq//GmjXAS8QHQy5be/g0jiJdty
st1IGVcf0ovsXh5Hg6Wt8M8a4SOpF76ve5BRnVPw88ZifheAQUxIRuFohIpU8ivL
dM9QKoTKxrS1TnRDsJ0LTYBTlTptwh64dtBtaljoN+/w675AIZdsE/YlX70m3+Pw
R0ifN9rWoZfV4I/6SS9E8U7GEg4OM18P8LajRwBHAl2hN9PEv8UlZdYwUailcL1D
OaiWBZcP+sEuoMNJj3X4obJU1uEspdrP48izaWipQ2tPVYQmxMseLmtwIZHY3ecO
EJmziTnG2S6d/yPmR36pXJMaXf4803ad78caZwfRSjgw/LqPHetpDu9i5qGYNirU
s5eI76RqoYGveQq4gV8GR3l0wiHPrfwI9Q2at55/GnaWnEG68k+pxnjAc/vOSQV+
CIS51vx5zE9phpdFg7rjePt5KEJqkpvsUD7ccecXsjwLOiL5j2RNxtsxiJfgLBAJ
VgmXZPtXySrepHlC2XQ03As+ZKnW5hY/IkBOx9NuZ95HNupcYElPsXALEBNI51q+
vCRLRejFuEM/LlJrGFb+c77l23eGnvDY5WO4sPXoLwtfV42ZR+HQDEZQKb/5pkU7
1DhfFvsHB8pcOmPbtzN7ovKLNyjoAUIPXGcf/4Uat16pK1vTfeNFcArWi5cL/3kb
vDvrAeR1TU9mbbl9ratQdYY9Cgal3xMy4W0PdB8QJyPZRNdwrLl1ULspTHLzZp54
tVRMrbfQMC5D3SwlLfKPc8xcOin4jXgPd4m9XSiz6Clpk4Uuo/ysnZO+D7/Xd251
oEpAyuukndQ0QvPBWKUm41kGVg5H8vcL0ssDmUOTaKI1/ctBLYf0wajyu0rho/Tk
N3yLWTRkb3/bbGW0/8bIjBuEvKVlXAB1fw4y5EWM5hy3MYAnUgtCc44i2K+3Tyrs
04s4Uo0Tf2gQ4awVY7xqWj1wNHNETmb4hbyWpnCw6J11x4CrGdv3TaMc7WK3Soh2
VJVFy8F5fF4kArHRa3+MkPm233lEYFaywS6VIzitnYAvWTLpTq+P4XxKipoT9ujs
/DwlHRRD7do1xxRXdIC/U1UtD54deb8ktkjNvOeiS9dBkk8WWoqDzG07sboxNc0e
ByCmiiaNUbOOCk90FkMSSPVbGXa7wTdPZrWuAOBI7yFInbuPuyQQoM+FFIWGbicR
sReyZSb4Ypnuqp2NHvqCCle0AYmckihGBANpkKhbBnaMtuMtNJvIknEOwT98HnDv
6fISOjfwXW/tPE9lAXJV2l9AEuM2XgEpUG0ECaNvBIhivkWXCsJUXvswhUuBBPLR
8Qj12/JSpj0nlCF9kCL52UH53v1Tfjd0B1Ppnoy4Edla+V56foXJi+YySh/UwQP3
ozKtyK4JjbqlRA+XmyuYqkEfcTqiMmIbWSe2+IdEVXAUCL+CT7+7KnIyImp0aBNk
sdmJhon9wHjn28tPSU/IO82Sw7WnVvT520JS7TjgwvSiL5lXAeEmRVLKZfVgufNc
nBxM0uaeHaU3SfXhrqhPtC5G4Q7x/dXfygHMhSEP1lZ82DmWDhudvprh+wCuHlV7
1lCoDn+skMzz9po22CtquW6HMXrF2vuBUqNW5pp/Y+nh6Zm8pfe3MXRcfYMjSJFo
rcFSIxhUT/VF82xGV9+HX+GZH8m4zRPbc6LZ+L0UMD4PdUPXrIPSRWLMhFclkQVc
FWozxM4TKXDecidEttaN+MqfOpmxXtGJDHmKA0ujD8ovYtaLoqrcP8p5tfyPePWI
HQTP1ceVE5y+htzxaA4+FqkFpuzdbJyGMm2szYxhiuU59EqaTeGcAqTAwDzG3e0X
SAmdWbNrjw5YK6dS+ejq7iFu/2r6PJjstA2yHOqrcByI1147g8+6n3Z0wMx2+Dbv
29VWJuWBqoSXT9vXL9ATLwmZu47bsh50owjzT4RImHhXXLn0uNrXvK4VtTL0CLgT
6SkDqGgDpyCE379XQvJrn0dPnDbZnwYrigd+BYWZFGrY/iHOuA4DRk0DRmRWXrJ8
XA/YolkaJlo0oi2zHFgxLFZWfKu/r4VawU4v5PVbxoUscJ4sfzcLrhAysrD6FSuo
diiZ7qk6Qdfm5s/Bg4ODvVqz/6u43+N03i0PNw70+XIV6umqcMD+T3qnddfbn1S3
WJCiz11celHlgewUapZuPPODPu0axI1R+HIJ1MhJlJ/1OCI8i7FTzmZ2jdyp1IG0
Nnh7RSg7t3PyMDlD6p1IEiPUYp6JGmzZQThVJVtTMsMnDN7mKUME8+hauPTLOlTs
aqLDU98wdRX52cfiZBVzps0jr9/5hKKYaq3i7K+2H1D6hrSaWGIhKOTM1D534uQh
QBSs0x7Ga+GcIrLiuq35jpgH9o4DXu7MjLhldnr1EasTN0mZqdffALF59EWJX1IA
CFYbQKvqfgkEATd45o9GOIMwSGSLXLDujPbkLMnbBeR8zu4C2EsuSRuS+0u+EY//
kiDxQNXekbJ43+8ng8XX7/K5XFN+hdVtSNiXXtgcdYLXDtzC+x3DrK7oRG2iYuiy
zHyjS7mC36KA1EXAbeLL7cE1tb4/WDqKOBwECsmNrTGg2cPJhD9gB/f4p2H+XoHW
2aCkJElRpgBWWsx7KHPNLwnyuiVn3N2QRxBB89F0wn90q9A9gKHs4LeTEW4CS9+k
jOc9VbGGOl7TH1e34gIg9mnIyBVlGE6/yjMUqw8svuFr1eml9Eac294l/VcTdag5
UalLrI4wzlqVjqKmndaYgmRgBAarpZq993pA8WRE/klubS6cH+PWWuucVuk/QLaI
Ma5Nmg40oK33HqncFGx1fzP3xzvhtOzCsmQVZKXdukHWyMn4SYanHG42aEsgf/is
W2FeheUZ4kUJCr668G6yx4RH28E7KeAq7Zum4Qsk0gQ2SXjstQE/saICaVG4xoUZ
NKHETq6hPOHIWrVkWB57QT9q/W78cz4npF0lm+hoEm/zg4Lb1EwZDZ+oUKdpKpzt
j22Afus65WTf+I5hd1YugSgpnZrOcHGAaR5Mg670pjFiGzv8ApVTzXN+T43reL/j
xnta1foQJxQiZSsOOjY8crSdbMPngIs2yUw1Ho+Sm9WLlVRFuaxs/AUfbq05xlbi
F1VbPL547Xz4I2k1XzNALEsMZYBnRpUGNm7lZfLKPoGCIXkMOxzqj+mS9uhi1zKe
h57XAzotMgZ4yBfkSepMuAtUZGuG5M3p39r317XNN0YkKpfV5ASFzF8YpEwDbGpK
tYBnVB7YtJqD3paqWtrIpWCfCeUADEQ+qJkxzcCwRQlUo7dxBrsqv/j4cMW4asKj
h/PAYXirHZy/l7UxA/JR1duf8YRQ5Y5JYg/qr1LxwWIh039rTEaPhRXkeJWdiE++
tWLcxd/qe5RAQLVv42A1Qy3eZ9s7DW2ENFiAhDlkU09Ud82xa2cbm6422PYJDciB
OPtRXFPmMXu8bstB0ITbGM6dMFjWfpE2BA72yVX6/UeK0Xxx2rYv64NhOGZB91zW
vtTQkCWlKlq50XbkaVA/Zv28PgueIjzwgA88zEXIlLWuYsnmHL21yrXla5jZtEpe
+M4RonAV+QEuWXRuwUT1DiVYZdblI3Hiyhwrb/K1vv63jGFqvTjg6eZhO9ws3hkW
z+D+CFfY3BHS26iSfaGE+TrgvR/wunzoBR0wExHJF0riDC0U5V/5uszMTqiG9Ohr
SZwxJbaUEX9nEnDnWg3hJTivUgmLBIpGC5n/jsINlppoCXBaHsk1hvzqUj96uYPy
WUI7Rxavv3dnKjYwtqE/EOeXjJGhhVUk+Fzc/81k1+QkqyR1IACfg4WjFeZaqnaz
bHdibsrtoSCc/BqMZ67M31viyLKuJJCUgtuyilTfWbGXm6j6OR9PuwHg4crsvndA
sqLLOfNHrpoplwylDn3lNYb751u6HS+vWra+gC73jzLGaXw7/IxAQCc+wapxVlR6
T7F+aXlIbNBov9+LC3idIFgT3R3tE42cEHB4/m2LPIcjLRDl8I0y5BIWbmPiuSK9
MlP67dUnIqAEOvmFTfYPrba6eRkjmxF2WvTM3NPx7Z39pbnJUdRXtwIfNt2LJ0wi
9vHh/5CSFymtZM/XVTbBw/t0S2GnuCVwffrzGcnc6RL1jiTvsBfw2qZqD+94p/hU
fkhpzZL236cQQuJD4JnMlZWM8mG7RGWIt8HGXL6tiqbVQXYWphKzmMr6QMvEHJOj
+Wz95V2C3gTWoOLtnPoJWJHkLjxWIkFJivM6JFwPgdxgsStQmjNYMBGwTo2lVmho
fIXx/95JHmyjduLsx4c4vynH5taL4COZBxJJfDmxNLptprVjIfy7JQRvVA45Tw2u
0BcdRDYd+B1OGgfIdoQipk7ro4xDMNYkzNAOcaF1ISCft5KWi9hq1Vfpjhm5wQQG
Cou6dEgDt0gn/T1h2gcIg/bWTOpnInOCrN0l78CBtdFPk1h4yj2ydT4Mq2budNw1
pPrNb1j2Iz57YKQzh1i9S/DeriHEV6bObv19JGiVU021wnSIZEalXlRNAurke1xX
X+ziLyXbxXybtFupn0rYtMZS3KrEpBouDT3FViwmhBuAEzeH4CA03p1KTeLed9AF
yPFM1gTg2LNKfN6Prh/VI9h/9xqG4uvuasFD4zEH4hASbpemgzPAaLeA/FlocHLw
KvwxehH1QYKuCn+AkqLZmQ1Rwq+AuRaSPkkRkv9ErIIBydR+HZNm9GkGXjXX91/y
8Mu3OGPcBouS5tpDOSbtEm3yswxERJ1gxyHFASYprCCqkbsStpTqIi0ICN2A/Mxu
5UG4mb2tk7gxELNnJ9BYpp6EScZDvvNuxNj8/0HcE/qt4FbTJ4PJjTbMLID3yEMx
5hWr9rhjEQhkyzltS3op7VKi6CC+pYWfk1Mg33rp7/ccmWmd20y/hM9z9WqtXfiB
pOhXSdpT24p/0D5ywkINy5Awh+/OPdRzcpqa9v4rA9sGOe5ltRyFUwSNDigC+y7W
zjbIWCcKSbpH44DTcNLU5ER8OG9b3I/WH+IR89v4Qfn3lxiRKR6yaUZLlmJsep2i
Abc3N5SJrSdWjO0kOZycgm5krKw8y3jQCnsWZ0Py1YdTPP4x96cvjnbFRoJHRfnJ
o2S5RaMctT8goPHJEP+ifB9RTJWr6GHO5M8fe+RCdtZwfD+SkQdPC8GR626Zlidi
DixbKUEwjg+Bf5L192zVtih6uQ9jRiGAxKs4xdFCdJC9RstmuYewm8MVXcTT19JF
1qlw8abGrHhkjRRKqJK0pNpepWi5p8ICjtpxwc6MvswMyNSdElyOhqqpXFGmznTY
HU9j7NLJHbIL8sFVrDsHntnafWv0KIz3uFuWDiNArClCRu56Ik56VRasxLpcGE5d
q7vrq+MEf3BnZOEr1FWqV2iASZfK5C0B9CuBuZqgB4EXXrH0V4aEObhrNrtUrgoj
5qTk07QRplPJCVaNDanuIOYLhVXdDq0SguH93wkwAmBZff6uz9sd9h9zl60+0xEE
CL8W3/ugZnBi6tV6UTtNDsJzPQH/j+gauwG1XWgtG19/G63RDCgaK9c08hvRZbWa
JHXJas4A7Qag9EXnkmdubMz243M94ZANsVh72brfapiECgRBeMW1OOKAjMYMxJTu
bgNETIzHnjxPd9oGOTLXffmQo4S7Jbgk8qKpG7l6v5A445XyiU93ZzIewcdUhysf
UnFsA2eVnAeD71Bs/O90/dJVMlXQ8uKzxGHHboqNO/+CBZ7mvF3qS3GbKId0RgNF
k+uUF8iQClRkApt8Qd/N+5tT9pd5toa8is7ZaPeOB9/ii598PdusV7Lg5lS6+S14
DEAkWWgPzDwPmVcnstIzqsfQ05XPsgqRIEG/sN2kSi9MMIjtEjtfFTN3OiQjXTUo
/YtcYBWvjIGQLb6QvhjfEJBjzhWKsJ9BctZspB6O6NYGwr/R5DSF9cbj36clQL6l
KsL9diOVfMyqVD4hMtYXCvBaRq22Ny7zj1dnVQWNlO30H0x01fQqya/ttKD2UwxG
qOTZfILJaeNi2IiYsKg/rqaHEZVUEYWxJXvwA1mLOzemLDV4GBAuSKzHrxrf4R+F
slD3JuGspSorC1Z36ahp1nT1ckNTRumXHRGJcTwmUCKnhc2L41YeIk04XwtxJYFc
jNZGgqoOKkV65abvQQ74bJA94WBJhud+TCR8VAXAe9ZYOLuFhLkg7Mef1JDHb298
5nvuomrS3qr4cupNvyujgnSAAO6VmLq/2fcBMmEA1L4U+pPzAD4uIuMhU7AjyXF3
n3/GhfovToH+rwqwxi5lftrk47g87uF1hdp3bcWog+d0Cv18Mr8dj0GS5KSil4wz
o9FxD4JsjUAyAGRbp+wzKEcpGBOzhgKVzPEkKtjXmcXp8FbRPWLrFFPFlSLbYOqu
Ir/6NUTxxHM6HWAstpEeeFWk+cjuNxoQtAieqfVOEKMx2bTjjp3rq2hzjDxid8PL
E1iZgNI3cBhrLDbjaQCgPLQDBTqsjyNAZU1zxfdG5Knl4YHWH9BCEibRDwSk4xb8
L5inQIp2ZymfjceoI9TARWLm0Lry89YXfv1JwROoWSGFr1jMqsw38L/MiDI8UtaK
uP62EJwajAvETsWUtNNrs811lCio5LKNqhHXau0WwyrFmwC9xzA4jGVI6VjNMQQ6
ADJ3XaUk3bb43HD58V8DYZy5QgEXwfVwQ1W4vvp64AReeFrZzQpcBQa36NVFyDc6
C/Fi0+2rG8ltaTfUeZqG1Yzzue1wdEKzdRYA602pmOaJDkZrbNYfEJ3NVQD1m6Q3
QODmUn9fGJPPg/S2o91hSV0IPg0aiNElA5mQAN8qb8gFq1NKKbxT5S70+iG++l6k
rjo4cwi19OPsJnTTAAWlD7IQmCFU+h8rlNJaqSb4aSACN31nojbnwjHdLl4PR3uM
3kkxVI4Ti3uKbole4hNcjUQ1//qHLIXWujMTH7Yf5Ydl0IZ7ylyKibbry4ENdUDX
0RQ4IyHKyodWjO21wpfwkGdyYg64k0jLGfRSg8WyWTNPR1WgoQtTz2GIuINXCXBe
B0HqoxWwtDPT9Hz8zUWxu3nzOaQ+DFHLBh/6nCamr3jjVS9n4wDHEV4qa8TDpyuA
HIBI9Ey6iJhYWzPz7IQhOMGG6LWhj/dwpAJRTN3mjOIDxyFBqs/4f/v8cjofzONz
usfvY9z72W7hi72VNoR5sq6o7SyGaUHeT3xdvemGvd/NWZX4Y5YPPrvwhzZZLDms
h6qapx86MTfL6b1/Q2jsR1i8wyR286Rlnzui4E965Od5w3LWJR6h0+JkyqqpOFFh
pQcQqydDFyo+JoPeHk47LWlAT4a1G8wThFay4CclGaBblIyjw4mtawQlrdd1jubi
/LLCBd5wlIREmu/iX8bu4EYPvzD1XQCIiDJGwDhxs8wgIAYFqY3Z+1XkbGk23T4J
PghZIiJnWurnA6pBDDjFYhQaNm3yefL1T7iV44+Y2W4vuD8hXKzlXbkQEAfRHw64
AEIvO690yyBnsyVDbGqR8vXweCT+T4CZLU4HhX1oq+wwdaHkpxadnR5isemmSBoA
RxiLhYolMmK4kSIghCX1h02NttvXj2jAbRtT0zKoQp8nx/bTL6s3qVfn+JCkMbfy
nh/Oln6wYPFZiVXR+22mDn5U+A6LTpowMDdTvTxbHelk2uZRWjeQC01PT9Dm/AKW
IM0OKleSbykl8RqHNyDqgNIaH5udwh6QqJzcADzi3byLj2JPEd7neFrBtQ6qS+Se
JKrcSJBb9yyDCo/PxkkN0REn9l9kB1IzzIPU78N7iNcVv7P3bwErJbs4fyTIRi/B
rcHlyw/orqRiKeNMUfTHxGFLdnS69/B+/b3AXv+F4Y8WwNGa73JNbhKzuJXe1xa3
wpdJIaCBFw/32IR9zrugPMD/leawNOkjcHk1rEwFH76/oxz1q+ldO2q5GyWJKlIh
Pk9tWTQPucqLbpeOCWSnrhsNlfCS83eoTJeK/2urCLhR+KSU6S+LK3jJb9X+ZWqI
lDULGTaS8ED1P4W5MJXjqamPJxaKi+4wtp0Rzoppx1+27laPipTeFcvmnGevY66V
FWyB5dcrB7Aa7/G9w9b0bYStRO3ObNPpYi9010vAXX7x+ZoOf/nE92AYJE1RK9UG
lpFByiVjAJFJ0OdnBlTbGyTlwD0TB0aFzS8f7260ez54PitzSzzPwyE1h+8/hz4C
RD/3nBWyM1SXO7t8s8/sjZCTijhvdCerekAciJMNGZhgVCPZvYM9539NTwl3VUC8
ediMHpqvILG20USKfD8YNmtwK87KaU5b5Qw3phObarErhl4faQ/Wje5lZoEC7Xz0
R0GKK6QZfffALnRbcCJyAKzaxGm1Brt9DrInIzzbn2XsajKqgHiYx554/X6I/12q
QU+bmWgWOld9Fk08l1DTygoWo1aqhcIs0zZDPHnXP35sZ+Z3SFsnbT+uz2MQiodK
Mjp2/llJI14YlwBiPxYJEQfHBX8Xe5GLuUNvXgXBy1iJzEA127ZYgzqswu46a8XX
GNw6ibLdAjTljNn1XXfB4PZ52b5EcTyz2Thuv/2/xjT930mp9XDkQN0FGzpzwqwX
N24FjTiWBWMrgrVZeRFeXzgcdDSlXEvZpCrYWItbBmH2GmUOUeGnbOXHlj4UlEg5
nL8a9hkmeXlZlohQ3JuKCvfzDrwkS2GFA0/mhKJD2poPIX7SILwCduRhXFD9+75m
TKLvar+tlO4RB4X+e++X7gR6RgYQoH3sfA7wjiZ2dpJg67KBO2W9gZdf+s2YsgLF
XdXTYDiJUPaY+LstC2B7bATPrZikQPxMMHUKXs/F/rtT5wHpe6v/WeA918CpK4VX
JoMkcyate+cy9vq8q4SzVAbqGqVguuk0gpGOnHuTixJbOVRR11Mp9L4eAPr74EMG
+iRozby+hbzJyyj8KRwBKsF/rwQPXwgC9NGGUPeO20EfN+p6X6w7f5c3g3+Dc3f6
iOaBTHtSuJ2vbwZA72St02LAlUHZFIVUP06/08bDdIEb5GWBIiJq/Ji4lwnTD1t+
nK4SWtqCCIhL8vyMMvDUuMuhHYr5MK7+fxo85kyQs6pWdYzsnOWf8+gi1xnt4PSO
Yp1/c0undTYdivN9vssjYiHQ59iydz8FRm0yZGxBwWmxlMrJEgt9QRYLjarPCJpE
xlv8TsQg9OzaUc/KFMCOZ0e7v6qW/C3sF3Na9tuKhOvnyonknZgaMuhThOgEzGS/
YCJm3wePOy7YTBFwF9Uan03StRWzwh1sOGVEUvVQCb0JaDxRb4G9WEkJLfZ7l2jm
yuf9FWzW1/lin+QR6gVCzhBtgehtWzMZWkRgTs6ZvZCMv3DSwQVV3ppXxyFm3XKt
EB2171qyjMAnUN7veBFPXOza73sF7DqfTADpMN9pxUZpS2SF3mFd1vP/0McX43xC
amB9XNHVgNKVTlh5TOolOTWuFizWXYywLqzrlU8VDCrIneS9aK+LFIT0R6h0c2Sy
p+7kmSGf0iZoyP59ipOvQpad3JPvz9E+g1M08FEgIt0PA9mG8Rr+mfGQpbd2+yqB
AIVOFNNKnz9MZ7/mXLcHF+lRfBW16VFDvAiXbqu7XmQI8QDtW6/u3LFm8aQkzgty
LzvAmBeVvExu9rIZ3McStNK9CM9euHEZ8ELhwXUBkt/ZfcJppLuU//c6fp+iJneq
Qtifi0X7rFThuDZiBLWtF4UipZ515F/cGo/bueUA8vLNVSU65ZW+XJLIp7HLKEMs
y6pW+DDYisgNlemDJXosXpIpxpMbOtpwn/ZIPHHFSEdTu8U2PeVY8pg3AWC0v8b2
uZ9XdFaH2lj4kPZza5uzVjR83xAg1K7zj0KC6KkJ03CY7EFTu4vf0QjFtZX5BYJb
/zjqnNeM0v7ZrEhuK28wnbxVcJ6soYChBfqC2HjZifQ4JgFt+lXNffl4RMUbkYak
en2gz6sabZcftTVUit/iFu4CqPq5YX28JxN7r0J1Jhdl8ZkHwBxWqIOCSG8M8crK
VTf+byyJrCLzcEBx+fIkgTX6k3LbheCLTw4aaZRrAtfXjlPP9dzw/y+vhZfG1rN+
kR0Ej5ZwRynFI4jEIdUVyTG+3s6ze2FbDTea1RH3DUGsC5kmUkK7YDef/jXWGc8E
qxsRIERJg9FKHhIIgCg/fYjpkK1pIGzlqj7xyMjxsfAkfnTwC6n9HtoWqcDZxVPI
9UJbsAV9OEDIrxZUowta55xPq+48/k3ok4YRIeKkrED0yAnDacj7Ea6jHKyNliIh
EBYn8WPHgM8wEIFu0ZG+WUrLSLRCrcoAPqKTedTO28XtBM51ecu4XcoKdITk+qvl
cru7Unc0TaCbdezpt4+D2G29a573pohEW2hay8c+tzKIHSrxmbO/xBxcPKXGtbnt
/D5WdxY60QeN8zOaNIbyX3dlqerbXLMsO9yqMllyy8Iz6tIIJ8tYUz0W3l2mu/CJ
lwdvKGNv0ghBWtAOx5+GGHSo5kLO+BFI/UedoRmzZpAqCnU/YhW9dtfHIdcrHaWG
JW1b3fjUUFsxr3CrCd+sizK7s06MWAJC3ifEl+9E7SxnODVvC8WayBUvCx4XFIur
YPTr7Esii58LcxN6/u8+fW0V/oMz7j/5Ofkrh+PdYY6zuBoQLMOLq1GtvFTmJwUr
ZDj6f+1dTctdGAYB1UL4xt2tByVj8mPQOYmAtJM1ow+yJceb6RgyOcgC9JbbM6/K
+Y5lJihUa1JyvLAXn9MCPv/7zpvCegcqkvWHd61+BYn9+p1vSqLNhGcDhgPx8kh4
ugRNAYOMyIblFdB9eJEiMfHI1fcda/bv30x0vNtJhkC9wdlnfBKqt+Isub6LzBfI
6I3g+H7Ac35IvMm/GVRuBtGlqr+4czDzFqrmnbi0ChLRRA9k/XMeW7Dt8cg4l7ft
RjSQxFUV6LsklXyMqAK5eiOGd0vOq5y4pRA6FMsU14Y/U8efSHEnpDXpRBEX2Tr0
TK/VDNjQhdtccM5KiuaQf1Wwh2Vf/4UOCUiqV4FJwg3dh3OxKA7Ndcq1QC64Ud4Z
/R6ueE13zS/bSMqbhZWyR7dvVj+Gnqcq7WJ7o+WtYctYOLqDxNBaJfFyW3XFs7fp
dRTDCQjG8JeTGohl1T2DiqHRtB//+rdAS+MdGeTwEX4aZH24avy2u/EfW5arAfQI
LpnlnnO6OHOEQA7GhoAmlkdVH/ySKaEIV9JsHcLaC52oVpF88LcGnC4tiPRd/ekf
ONHiTHQXaJFd5gSnu1GdWBOy1oLKpqD1L0QtpiRQORvlZc8F3WxXl99l0+LZo6ce
2a8aIMN86RZaWCIrd/sq+PNxihC9E6YSmnN4R73nZpHw8km/PvYWdFJ7PC4c/Zkd
1BjSjavbuGSNpKsI2z7akgOkWo6J6/QjLm1D9R16IERLXnAmeD9mKoxSH54VGpAB
ZPpP1Whuv1j9hjE2otlTsRa93Xz/tXhF0izLMeRluvCLYN4sgxIbcjLatgjpb4pH
jt+F0sUNc2v8Akj8e4Oc79kAzw4RjUinHJ1g3N0gsOaZyxdGl8OT1ecJM1+TYU1S
3T+OkKbxbz2relSBIe8WpY7U+D9KkIclwjOdUPtCnJKQ+hVDhLoO3svN6WHEHecW
lMWM43thTTHd48/fix8qjgsX8vi01K9BLvYEwRJJQTdt7YADm+LuRrkzpisi5NDN
8vvmAKW+RB0owcr+kHoGwUuRPyYv5r1SmKPaunpUzBCVkcbeh1mHQxwFEL5hcCfz
EtYWAcpD7K9Hvdi4SZZ71iN9JbbCfDmwYuGKtxqbTCq127wEgaOsKK8lraGN8TMX
ktuvqNcPGm/43Usg+c3npC0IBLRg6mR8GE8wCXcbudSIXW3y8CzKj33AvX607ww0
gsmeO5VC9xLhSPIqvj0Q1V5RQ6iWPCOPgLePJVffAhlzghoSMToWLeRq4vl6/FJL
t2VPz73isD2xkZt0bZPsFUqWV84ovDrjK28a1sI0g5WA+V0kuti5jQ2RgN1ttVnW
1ry//VryNNoLwbc/1a4ifRWRk4xzSz9/tR1tA7rrlcAIWINMyqClgd+WfHUXqWgX
X33ob7Jpmet6SN3HeoWMNekutmz9kuTw/QA2BC99dv2y9A8S8C1T3gaTzZsEUWm+
RM5hLKwRhacCpWfV2Q2s55EkMdiNi+QKsHhYdMr7dWXUroUYOF6oBmRf90SUyIrx
OZHO4uerhEntDMGvbNJlNmE6Jcnp7nIDnqrtYPa5+51g8AubQ4P39wV4krjyi7EQ
C+WJ4B9gYYS+EiHyBhOxeSLREd4p6TBY9hRYBIkc55BHGU8EU2MBA9irN8Sbfazl
y2MnidRDsZICR7UWTo+FSV5xiOkXCus5pfQ/gQJrGBK1nbP/egGgVzeNJzCE8TnY
mcr42H1WzafUDy3HYKbQqK5HRZPJjy/pJszgqR3O1c2Bi7P4Csq5qAsc9Tp9ZJZD
9wmKfS2Dw1wpOYW+WGOmSoqlsOVP4DDiwmdW66Ph5ShdKWIiMtyMTv8kxYTBrYGr
Oa/xn8cKb2TBs7pNG9aj9p867WLc15dE1KSSHTavzsOgKFXV2ClHbs0sd0v2ygCG
XTbBfmyngqF9vVstf7xDE4fVfBWxR1toVhgK4GOV/boT9GV15ftCBt8UBYY8tB+r
5ZEEjGX044r/xOdGMx9MdOk4tDXOCBTDtSvCJFzJKmD0lB64a/fSv8QhEi/8rLK2
ghkOrXAwiJR9dh60v0sg/9pfpDI4ZW+fGvtk+nbUVPFFeWqXyTCKW+e/B5jm5oAt
byMdNrI/ugTxvp0N7vkz4iWgbT97JZSRh3MtzdVJ4TRm+4lJgHwhLG/gTUwhTsmB
mmYzAKKBoMoIFtvUyZPhHQU2/0aqr/lmriaeN/NMaezsEZFbV7MrEAWE1MFfIVmw
my9MGI/68DRgclZ+hbW1BMLl26e9uvFtomPst2nymZXIMRWYDSzNpkrQImaA/4Ai
M38y7X5fYtQlzbMjXgTst0prjFxXk9FxJC1lnxZfYITrNBTJ7c2wLwe0nqsJAw88
jzKvSX1KvppqI2QwyiMZk8hO1QyQwUCj4siiQreTTJ27vnP7AXD/Dx/a5Z+vO+Zx
i7EWTTMRuz5wkooqDyZOECzFDwMT2lKNagECyfm7yIealjA1RPtQCGOb5kEkSXtd
qdP67ro8+NdmMHw87TafYrfbIKicd5+DNzFL11n1iml3UjYA0csMsjQQdafZtw55
NH/T1zc4jATiVNg+M4C8fEGv28YNopyC9134CuBtzQn9KEz3ZCMZ7RFklPxKPo8Z
uU+yi6KApF7hOlO0Y1PYz+vOaXiXLTSxD38n5DWwdtSkDdy1WhsoYY8OSgA3HUfH
fX6GINQCdibJyx5zAZ/BXwav9Udn+qODJVY8lwqq9qVr9c7hT9plmDAtWKY/3E/E
Yg+dhYM3nls3uPj0OELrhSq0zPzGn78uFXtQCS20KZpJiuR1bdTxYVbzAFvRluN9
BM4rLcxKcQlXIGyfvz5etaccvqYUG6w6lVMR+ZQVloHOgFoVepNd3DiRy6aJXJB0
qcz06T/KDY1BcGBYJOqJR/jyD0ymTrP6lOF9zzzqLVG88FVYvJYVaAMbu3Ijgtzj
bIDnyWMyxExZsIbDKUK+/k36s4MgeA/sh8o6ENIGkICN/n2Vg+o1o+qyTqBrwRXb
uQe+aEJQlhgayO+FMPxDYj4VkbF7tfrnF0amQPY3iIOSDu5gZvS+Mr/7ABC1bO+R
nO3uaz9DNPjTthxXo/h5aZWs0eH8X/Q42D7sRfhNo0hMt/ZoLwHWoidWBQfxdYfv
LR2igPPQgT5DYjzD2RZaC/Csny91BoT3D3nu9aGy4lMZ/IC+GSaXoX/FjiL7WwAS
tTl8eCS2cWK6u/1x4Q4pm/b6NBUhF2tdwEPSVb3zWuMOHtdFCEjE6GG++n4fSZK2
hR5cknpsdWxsz1iNZohpGOKLyYdvmd1jpzcLKw69aQiafAF+vrnwdwIfG8+lfuwU
jNvn0DzcGuQr17t2OFu/fQRhvjnpyb8OGqCbuNBlWdlPdARP0pTgr26CmE3hFwJ+
who3zmMvi8oA22BAjbePS8gMrNFNYmXmNnOihpwtaOZG1d6of36yVDoFxDApe3Bh
gWrjY7CpaWJ7HXrXBiH1HLJpOXKsr5D9APGgG8nxE2RG9uagThrVbhqqi1OrE92H
JXIQP6bFrscKB5Q5ND0YW1on2X4EGOLGiwVUc68bsev6sid4eOPaATIPL0gw4sQE
UGULeX7oaSMjbDy6cKbeQX4M0r1VANqGZUbd8RBR3aIm33ggF4ou4d41l1GEU2At
1oz+0ELeulXnOlHVp0G509hM0KUy/7ScaT1NL5F0Dc74wQ5IwsxWwhASq+h7YEII
XZoO1xXSXTovhAEy5O5qP5PF7x709M9ftl6JcxRO3B/IdGH4BHsKUd2usPmQYHvQ
fDqin+uZOR5FWZ+VrgrS/Y+MxbOk51ecU1ZKiN293YILD0JXgs/1w4zJHofwM/nE
A1CopQlINAKOo//RgWLKQq6zyk/8IByzuHi9SYXT7TKbX7Gdu58ADQV/8Aog2G45
dGAK2eDJQO7Tj2FlSu3xVN/nAbVseUXNbkRPhAVtrkPQzBnx7EFic1LNpkF3hdir
7LiG/JB2R9MJSy19Nb6VW2QdUbIiKaOtJuADrdD4eebjQyo06/MecuKqahqAuvMw
DYwJlI34A03cnGfydnQqAFa34i7kmMgfF+f31CteouaBbxxFcoZRUoQG1EXnGbbC
GKjSl1wjtpXAA3IQIc6KmO5xzk34K2SFoMYiQtY13oWa/uWQxZ1yOnhfa+NbkWRK
jLIqYi8vRkaLSzhIPsQqOOLUyt9CCQ/EquCOudU+i8DFDMOK0Ra1MajIm8933PrG
ZUWiHqY0WtcPo6f8IlAeht/9mXsam39BUJB0ze/p9fyjHvLBuar+ZFwhHfXWm+4J
iHS1e8G1fA74oCWv0bZPofRSMPUhWWUGmgFNA5yX05Tl06cOO3uNFRcOFg4x/m9T
1aCZ13nZ8qiBY6yDr9HJCBji+qUdPczaD3BFHj9XT6sh2zt6+iaaldZbLImsDRuw
33oNawT9Hgt3gOVM4JFfyQ8fOs994k499Sg1hVrDmfpmDgUqNkn3IpnlfAXwy2eN
c75rwTUoENfjCgxzdQLkOc9x7Xl43F7x2RA91mcX3yPJ3Gty3+WoNJSGD0FW5KXw
gKB2+HNY40qyXhV40z0l7W9+2c9WLyAUtAHJubrajUEGpPEKQjxhc42MrnyhLYvq
qgUzzwVsv+HXFdYnjNXR0JBDtHMzHfsKtsSIzW7QT9vycpRBwjZYAyth/u/trdTj
o1I+NJKP6fgYiX9dPrLhsbf2MKIwup0UbA5Yg9UsaCsgifJ5CqB39Ffb2BFoTST7
hIBiDUHBaET/YDuKsMvU3MDzq+cPyriRlWJ12veUkU0CxJX8B1KxS2va/vdkmXBi
uL+PmkPakChVopYCkqpux7vfv/3zJiq/UgwWeoXqJX8j8aIaCq5b9+laNxYmT7+7
EY2+r1bhoiGoRo22R87WY2vUe3j+PMblewPW/YKhr6PZtajZGy4/G+fQ9V9h4p/R
u+8LDuSZzBqz31Wy9ef3qa2KFaVM4MbpaXlyGGn4X0I3vTFh03majTnf0EBHksbZ
a9yDFiVPGvf8W29lrC7N4iFtetZP+Y69N9J3P3n2CYBJUo1bdd3KzXytEA/kH1dA
OXBeKtfA8HYdayLqGOOaiOcYmw26iboiei+YIeoE7DxDFzUFTaShr75FUUbLfSSC
ecgKUAE9VIrYDO1h6FV4LX+IEzDIBiNfr0Wgx56XIOAx3hRYSTxwvd/QjR5qxz9c
jBUTrVZCNYqrpem8h0bO60fcLnlx09/9fxNMB7D4bJgK2PmFCNT0KdvQd8nO9WMm
hdRWWS1jGkR6LxgzcO5UwVODN30h2p39sECMWADSGjf5kGYdGcFSgIP3N5W1+V9s
RcjK4sdysGGJDEwIXJd6L8g7u9ai0dwEAHqlCH6LeGK3EPsofUizS4pDBdjDFolv
6lukLkwzTatoq5kaMR4yIDakXpLYPxVGHx49oZDIZoTxgvlBWlPVngbB22U3axhc
Yp4O5UfkzX4YKcGGO3tAslPIIFXD2CjmAcNQ8GkeVVrvWDF714ztGqgG9I8MFb7x
OEhMBda3IsNhhOXpuZwgiRp/ZcliZ+HVpb8qEWHGGaxMN1bUnBLbjdw/iv7aWbrE
bNnh4ErrVX6r24v4Ut4xaa7gCHdfSl4dl83GsYrDBjfnCFBm8KuYKAyHovVEBMHH
oKaB7ZVxiH6Jnllsx2f1wWhLZamgKjMUUpdOGEkPefN4fi0nkiojFQISyYExqg8N
t5MfHBnLweKu2RRv+xIP7fOxE1mkuQsraOQJrjiBrYgGZQxOoYLrQ1znELQXyGjM
dAdF304xUiTmgycYfe/U1shnp8RxdKqZcUTbxCfCt3eIqJz10sRtYg/iqpDDbsUD
JoGbt0uNWpDBa67/HQWX6EdTdsWmPOb+7A3KjqOYZ1NimP27EWNQcSzrJsP2/xxr
buPEOZdPA3YMshRzDoIGNCrzqrDDeybrjVE2fyIrHZvVq4cjtxT3tK8lbwsbHDSB
WNTE1ymjtuB/Ajv82q030u2PYN2/o4RUbISsPS0tHxHMZQ3KGqkVZJIinC5wn4w0
RwCXzSVWfYKiuyq62hJz5O1/hN0AI2QcBsqwt6IKzr+f+nMcaMlFK8vNSlTwQ1GD
SebIuSBf8UwXJY+iCA/bTbLjqhj0ByM322VubtO5V57H3NkoVnkAjDLgIz7Audet
9xUrblpe8gkiPJhm4FKO25xan4G7M/27gQSgTh4CT1/dyZ+JkNhj6DyW3f11xAd9
VmVvUcKvN8hkj9cXOU71p9MM9Hk89ebRQWDnHq53tk3k6rXdz4g0mquzGSml3Y4k
BJpE8h3V4XFGMg1PEDInmpERfBDjKz50ozLlF2SP366LDUyODSmZeXMabbX5ugwd
KA0ebJDrFKd1wnmTT+1ZITZRWOHubtSSx4FU3qwS0q+Gm+DuYYVBQBlOOl2Uc6SE
xywcw6oudikkt8g6S6a2GOph27hmcU5VyGIKoUeIBjukuF6mui2c1/5ALaoMmj4T
MuCSSYOxm+30IlmuouJgJZDWdKHfP8WBDH3QU7wS/gTo/W0zGE00Hp2+Jd/GelIH
O3nj7nVH2IAAx1J9ZS0KKy8j8GPP7l0vkj2w6ED+BFyXIGceBgFGAKW09b0P3hM/
GGo5JtP333tx/ALBSDRaVP432F5a47XPWV8uCObZCpWdjEYhukcNZLWcDSkyNJoj
qJB8zXDP2deOhecS+GZvNPWbS3VmIAib/2W3OR2teEz8KuUy3mvpvTM6moV9xcAa
uuzn9mMB8THPIPq5u6KodWllMoLjjixVpkMVg9B0RRW1CR1iIBZsRfNL4Ek70Rrd
cjnLQOm1+JejstXtbYzCH0KHpFRL3TOtyJbe4a8mPhRSSlkSbEBnx4o2DN6B3w3y
UsWgm6O3XzcRG5lE1XVWDz8Qq4mn19NK4cc2+r1M/ieHcH2sF0TyvKgSQChfUb8v
hxIsi5JtVC/SInmTxS4O7s+tf09FbU7vozw/y2yQpABCQelFOok9aEeSWN5IjZns
pOmuEtEmDgmjifnkxgrxAb16JwROVGUg8rr4WBQjxNOP9pM//TppL04Dk5yPOyhN
20vhDYgNA2Dbo8RXTr95+6vWdOUnklpn1wBZNfgegraYUD2r0cjgGrzBSD4pncM0
WYGrAqxLSz/FSBfJF7Ee9XSC+2m/uUdjxPscSJ6KGHmw+conrfuEFINMcp+YaPDU
558rI5UCV/QRTifpKf1FX49C5WDQtpdzkgXdTszEUoDhyo8ItrQP+IEwupthJcUd
woW3S+gyujZ4vGTsL+hDMEGBN4CTGn0Nu+kBSg1xhBW4T+r+UNcomCltyZpyIzw4
VzJZpm4oCANxPXm0MAHVWx1vBAW97C7WrBdI9nQvDlxndRdUPXQO3H8dbEuMuj6m
7M3s4eZTDvSmx/frKjs3nBhhTQLNYxka0ZKF/exJK3unHB0fPvRP+zBuVqE0p/K2
ZxbDIasbrJAv0f8ywL90T+3AFALIwu1zwpZJU+DAaQ2GLO8bxpaIczoYf9kQ6YyT
Otg7Zul5Uc4h9W8guwNvAo2tU28quIzlMWJh1ENIL0gGQOsNktS/WvBkIH4dOscL
l6YwK6roUqWSFoTwU25b+uaNNP7lX8vwMEx4kwg/+AjHirDKCIoZWK97s5IXYQTP
6rgG85TY61OWLkFTbIBaHbhLvVvJGcVIAsyiR3+PZOC8QfaI2Jd5jKcppJn5K+BP
UFwKD5ZZ1Ox+Zvv6B79Zj5QtYM/3MhtiMMlLRm1P2aN1Y9fE1+FPO+S3NXGKdSqG
vzliayUqVE9zaygYecTTrbhh/Scjn79yYcA1txHmCTq9I1CPAI4ujjeiL12InZKK
3U8kSOKrTXlMmj7ubBeZ2AP8Lig14qTBHUXOxdouYtthhmbp6vKvv9iReFg1Q61s
sOnKpC7LQw1X9TZakwph+7VDy7xYIUqCx98GTErhumiT0Yh+Tmjh4PcEtd4UCiep
C6S22Ytpuf4c6I8Am1PINRCNMiDRC/pSvkbocUhoNuYngaeDhgSQurf5rStaJXKa
Z2YTpIjWcc+51uaYIBGeF2UWzSjlpTIYFLZmhb6BC93FRnDHzu1Mo3HrxxHer5Tv
RjWoKFAEVIyGfz7lEMrU293033e33rM02u0dbsM1C3taXTlMfCmcgAs2Ji1/sfuc
D04Xhj8PAxRAVQjEjWGFzpIFoJzSMx9rl6cvrTY8yOQtstW5na50iKL3JouXnXcM
Ss8UED4zqMHq132KrzDVruTvqsgfYm/ROGFShEq6m17B+nMPgjIhU8ez0ShGBWZE
nQfAQTAuDGCXAX4mISJjLbM7/DXP5Dx/82l0RqVbwiXBtgpLzj8cBLwSQGE/4Np3
1VX1DRhYpnb7v5ElpavqbJ+fymyTwHGr/Svn1GXAYcCSR+pPOetKOfI0vyyk8Fzv
IFs4mHvwx1fB5qlunLgj02jN6COs6+jAHlo+yk2nsKi/1c7y7m/7dY4Y+zVASJ1W
ril1AO0q9oaDVo0A4eW0GrG8ZbL+31NShqlIn6Yk+56uhyFgU/Rk0qUAwuwMFAPc
KX9/1/5DU99O1MCS1CuFY9mhX6HXD1+RXS9XA6Sx0ukAiFebRnDxHCLH7biqqmCR
VmDKUSA+P/yGUESx9gCuy+zUOxJGhKHvSz2bQLvnEPVOt7iC+NubWHKQFTloUOEF
wrR04x4YGmhISPMiU2N2fKaSD0McL74U0RBEXFCe1EFwDaxTGOcyhLWy/36XnPBI
FQ30pFEyTUQ1d65w0d8bzgw0O+DT+b4zNX7uQvmmNTJx5CPvEzGsdY8lnMTfaWq/
yM/15dRwjDDYjmOLEQcRM9M/D3KGUPx/SDwBZHFx7g4coIx7wntpYTb2/pkfeg2l
LE1iQ/2z/ZGKbR7vbCcHOSdo/9VyEpCkmBMP1YlnLTxY2aUp4pfPUmuyht03A0d0
NjjQAVrD2kLl7pxArwAXAH5Zftx+jMWs5/HWwo1VHYhd7pfqOarH1hE6F9S8w2nS
CqEs8W9FCPNHGVfSCQc+w0Znrvub9Vt4t3sdjitb47mz1G1o6jo3SvaCuuc352FS
8n2mEPoUS58FWXsmPYhBbbq7dEFjRKUORd1mPkCkqvJMdgyRIwt7H9ZPpyZwrWIi
G/iCrFpYhp4u46jctu+5wBA2jfQgRK8RJTVWxSyurjRXM28S/9lZ/zWplOhJK8ou
TWgqk8jKWlwACfMta95VUDmNrQ/xEJSpri9xwif3x+v1sDqw4fdDvTui9AqCbfKt
gqmRsXjpLU9MDvXlCA14WsrGiJ7gr/7YYdYaKCSZmH3gK4ymDIlwzhIsP2KKgvq/
Pvk3M7ftPqA7baUP8zxJHK1Mu2s4gZf8K1YttXAYK+5J28Y+WgH5OjKkqb4/wWKN
dnvsbLh+IFfjKL5XkYItD1WK4mnwTirDSVQ2bH8KGr7ufPYGY+wJGqC7Ek3RLFRD
xx/wD3QwqnVMpSN0EUIDudQVqAV2Z9fOYpSkfLHix1EF5p90H7gwiq0eDTN4Byeq
Y5f3eFfcsIGS1B9PDoNKld6h4DkrhtToxf1Djeb+TozCFzjlrLfMpWL+jjV3WQBj
thtKKO5W43SPgpd5KJC+L4jPEDF7qf/i158GK8zbCTVPrHDSUcu8293FuVchh1AC
ZpC/7ityONGI8qCp5+Y8wwhKF2wT/ZyQWs67jf+25VEwvtY81gT3Hzji8qNPt53+
9gSe6OBERXe66Kf/8c6ENclgl5wFONEQii52s3EanGCuxLQI0Yeq3VmLvTFnQEBd
X6la+5o6/FmIIhjEaUjsWVAzk/flatt+D7rIiXGQosQuyYd+0wx5Is/qMUQbbeI0
n+wsIIDrgeuTHlVCK6DySYEi9+NaEhaxIhN3rQSjzgop1KUGyWHBaBk7M1GmJCFl
WiUz3zQXg6OVQMYZhFn4RU306tSM9ifyId4Q4zUZMFdCifEmNvUn4mgB7PbLHrr2
XKfjGXn/zXObQh9aH3uaATQE9DCwcDoxrWnDgOSX5gJguLg0fPHJ1bXhiNRgs0ll
e1Tl3pKCXsy9E+hTgWlukp49/EMOIcUa+dpxg3TLO6uHIodlUJ1o3Nx/+3ZG5pC5
pvISWR9RRR0TnqnrzOUI9neNVE8DuDVJIxTsIeMK+0gH6fVcRr86HX3CcyaUvNi7
1nPdRIDXixUDhgNagcEKc2cqg0yFXSRb0san1s6IxtvhyPSs2cGVSBOMtHasHV/1
/G/J3JH7ClvgMN3NHM1GXL/eOrdGCwV/Dvah7IJpD0jcWK9M4Y/+9M092zanSjEc
eQS8ZJSk35kYYlzGAZHYHrQl69XtHas7oCIeZF9yvLouaOtMoOokwBonTs8/X3Xh
eL9EL/lI3F5viL65ti1Cl5wgOkdERwbJgHmCy7+wboe116E8K5y833Sv/zuPaFg2
2sqXkvVvLtPqFY/IfNH9HD7WcYhhBA2TVgm74Tcbx2vkEmdh3sEYjBCbDC3WYHGr
766vN7yUhbHZ4kBvyyUhGkcT4rTXyp5DHpDlBFpZzD7dv8p5lP8mdmcAGGeAOBjh
LJXmLAdVxPER069gQ2Hut/r+bZNdAL8PMOD8hknx4qWv99BTYnjMSJUMa5ZVLSWp
CduKc/JAnZ506b2u1xZFZg5WPCX2vigLtjHflttfzMVfZ+FaVtQpgCBOhOmN7ZC9
S/Pji7taVqccnjxJok5JTJ/xxObedPGTkyjqWe74ODHQnvsEUnuxlTeemY64y9ia
7bIDg+H0pWmIKuicEm/H/WPLdZLVn1ikB0gqPB91NiM4ItMSlMrma/TkEqrd0lgw
4LI0zHGkFET+MCDlO1mgZmIRSIjKl7jj4n6d+ZYySr/8IRFdpcvTX5Lrz6ZxnZgr
umEBM9gKyIV2IiseDHcX6fQiQAFihdSp1d4qQm8nxiiwf+RcgRxm6raJ88gRtFAe
Mf9cER2QkidWGs5iA1wkxwxsF1MBbE0kJCJ90TRbvj8NgFRkB8VxYVb2+ZkU36m9
zZLc1xp2PXZsOO7k5M+EI9ZwJrsAaM7zottPYA9CeAgLCHL68MMeILvlsrF61GYG
oL0FeUjPByLpd+KTEo2LVW3pgPCfhlVv67idVeE+N62mfGc+sU3uiWlPjnpzdL5y
akaIKzFGTG3NpbCVR5irgBd0qjkGpLYgmWFokVDeY0DTF5qGvZ0g24bd10A3aR3N
CupzfmSXBkdGre6oqfStx2MxsWxASic1dapbCas4GWp1VhMs86s4tXmPPO1GJowr
T0iorv7u2Gd70t6uJxkkHqysoeWSs1tjrEmrHLdDTh1jSCIUxaOiclfpWBBn8Zc8
inMbxqPFDld23ynS3x4NK9aNQjKvLGFE0rSTdYr2nu+IWP6FJqD3xqDd6JEKqNq0
Gy5IIYf0kXUPziE9EluW0ky1RuCwdP+yD+0G3URhvGZ3OjtpRimUYX316I3wRUnh
CZ6Q/AZt7XChcy5g7Gpt9XswkkiRN0S0g2oW0nOkqnZknFV9XE6uuPnwEarawFIx
fsIdVZT6LVD9DulTedBGNvZ6LTdMHqpxbB4J2SbjzNYHUI6h34Vx1ZH2+fujM/Uz
XroCOiFh6EqqP2jmMA0agwpVP+BlRVjy+1sLDDYcc4alxtSVtUFu4DgkFN9v3m41
kZvnT7k1ZvaoaE2YWXZ03okuGAWaatC/8LrkAT5hxatyG8MjFX6il81vLIh72Q2o
vXi6tdwTSAsdw8v6cZ3N9rb2OzZ5JwlvCz5g1zcAIzj5llOrIAiyAuw5fS/Ty71J
NiZZmoOutMxveIhfP91kO8SRLgRVgLiqtW698+6qB4JNn+VWUpBZ8+VF43/j41lC
QmfHXw8UP9J/Gb7aSTDk3Sy8FkH1hxnhHMIVNnkYrxJ+3+7lMN0UsbKrj9gWxKsX
zOS0YkH9Nz6e23U5hW+fuYCVsFijU9eKl7NzaXAsIPxVHs4TLn3qUgLrXPNMcSJS
wPnlvj2mjOBJS5qgjmVJ9A7jIA06fz4x3HffU7MhOKc7ahWfvWXq58iHyMhf2h82
d2d82frKaUulJQSuey8YzegAORenCJ3jYG9nFsMIPGXPdYLhjbeLnKhLW6nGv6wF
osrrp6mAJJ00cdHrs3CJ4nx/Rih0RMwxt4q0JdIws3f3GQrSxIF++Cq7azyFqaS5
65lX6ojkjxJkK3ohGoK9HaVkO7PBqCfp9pQYzxxf/MY6KiFoAF2i/+LQ0aoSk4Qr
Nu6Haq/sQ91vqA2nJMYynDBIca2siiWqDXAEfpB3pFd0X+K6VAnpxNlgO0lUJ5dL
TRfYGPvuMHCCmGy89BYFUIxjKyC+mMgGvdRxIbAO8MVcqBvhVbGPkgUVTtbElQmf
ucE2rX1Jlr7GBkh7ZMsYY57ti1d5PWeLTDbpNwjeyE+a3t1u2vwFMU17fEOPhuOf
KqZqgY5tPiwcieio6X2CwflcePHZlNCorYgafw3HY1U6RkczzG4VBBzEpB1cT1Pp
K8n1H06wacz/wuMgD0mHoHDkzNUF0etDB9A+kb3JlaCOzDtezuws0jJP2RdQOgfp
f3oBgsTCJ/bwgRSMEwJ2g9wIaI9zwuqoKWVtCUn3p5U2jzehxb8JXsbBtA3GSXZ9
FyIV1uJ3jcsFuhtSOLVWycYaE/jWrhhdHhCJCWpwSwBigV7blGGF/wfcISKwimmT
Fu47aUsI7j44ChJvGIpjZDpDy1FADncph2NdGkegJApc1IN7ctWSt1oh7Fzk6s7u
sePyeZEepPdRiJZSQVfTDi+QS7Bjk5BzpVfvMVfzRXuzajv/M2iyqFAS/XgQN0l5
JZEbsW43jg2GR0dOZPDTbDTGbL848ofK18sFrbKd98RV0RmUJLZGNIlfgPCFYMc+
mb9YEeqxG6ZqcsFbYTZAD6n+FOwlgI+TrcDornTaQVAKxXvvE1kP2p/hkmyKoz5f
du+GIxdUEwGA5jefWL2ErcByfOkFdXLS0nJk3iYOevxLFfAZ02bSjNqb4hjSVh6d
y/s6gbbxIYhU3KvgwOWxBS7nqoNnpm1JMTpxSoI+RmIVd0J86RSGZqHiUf0coaKX
L0nidH5LgHNXkYJiSEOJE9cgDB/4QsNzjVRUHXjEcvuxUzEpuYmvz2rn07iWgBC/
GJ38k0xlhS/iuYVXgzZPks9Jz/s3JM2Hg3CFfhbCBynqPmBcMXH3cXjWEwjhM5Cm
eCNgTj12ZdBt8R0Ak2VdjEiMSJe2kfKHROkx790r8fEfaykib1D6MeZERLNgvI7m
OZqLfgO+FtyyEn7qBortrIiJv35Pk9XEMNgFwBqrO/WuKaDBeO1c/IK3r90yBNtk
39pX/zK1kDK3X2p2qVvBvHsFPpVMqa65XWwvA6+D/lW3mNa21/DTQ/FRP7BQD20z
4JbtwAlrSQr57o5T2GYR+174YOgnE/Gdvj6ttX1HP5SqtkfJ7WDtqOD8m6yDYuSv
gXuWIYXolz5fM+0pWjLCNzq47UXPPd4LJndCbHuvv3oqXdKaBBjx7//r9//9kr2p
YRczASao7nIwU93/dxCygUwIVXIdW/Mo6VOaLeukcTW45mlqrMfBe5CNOGFHNonf
w+Fu5kR+sQ9GYFQCiDlySC9brRFiyr/wF9lzSrrUccxXP3FLzRNNfCG3z3ISXgz4
oJG33LpUez60fD892t4viNDa0vneZN28LvQ+0MhUqsXCufMfMWbkkDrUtV2rVmXP
fG5na/Nq6c40sB8txrWcp14yXioAw7wJDMK+jMXi33CRgrHcEwASvO9yuXuzQ/P2
jdno2rbc3whP/XqBdTHVbumeYWfRNvwNYbY/q/oCFsdKCiwFyFuok1ugzWZbDzuC
OQryLGx+2mMMWmaiXmLRZ6kgTm5HNMI58FyldD3epirR7Uyk6W+4fh9N2XlPGZLJ
k22xX7BGmdhG9ZoRn44HeMbFcQSIATHM8u+F2Z0tZQPFCMfOJ5xWnoen4nkxyQsS
yMZcq/r7Fs3V4pOx+L6jfKupRhW6vSlvellrnJsCXtwY2sM9OiY8xONAlKkqu8+n
z0BPS8/8q6mOTAo0svYixZUzq4plgQ37k1uZ0+UDO97rLAemW610vnSd7W2Pzaso
g8LyPdbQWgbG/87YI9qtkf2y/+MWCo3nGPdkkWgz1zcH+/D0AKWxOx3SCUPG/24t
2e4MqvhJlk75CNSfQoUCIyGP8qiVJi1c6J97jiF9qfk+GAbAPxnsaxUUhdv5M3AM
JvsR56rmpApUkigDWPRYnIE0cLwD8OMTzI+OyFCvF52jKkVAYRg0Z/kYjGMtjjK5
BBeQzDFhNCBV4CNxvrB1r8sUiPPVv+wSXhpzTkf3WRAYsQfXEqJAysfqI58Rw/FK
u1MvrASCooC29Nk7uqqseeRjvi+uEqd7Nln1GvdxWtQL/JvPFjwfmMlDdp419eDz
bqLQFdnfECCQ76N74MDJK9LoCYjQxGcoZambLJJYi/OLgzi1iwF+E1wG3zkwNu01
dQGbtbDLqNs/xTW+MJyGKLvj5d5xv3NilFMb3jVceQFY88cv/Sresfh6k2IluBC4
4INE0h+EWUYioeMEDMXpWwFnp0wuI43yLND2L4q2eTYrgxtIbnWG3yItglb3tugf
BmhuPCCN0QrYqjzTWw6bDnMmZxAwBP116FUoeVr6o+PwMDtb44VhmrpheHxXFtNz
vMP5i1C+mMzLx6q4ZZ5fW5ADiadrT0a8ELGH8lV3QCxdGLxzkTA7jSXqinUte5xt
ZD4SKM8HcMKitPXedccXj7K4jvf2S10/V4AHtvDZ0PLBg1rgcxpVcCFLksVKi2Cu
k2bt1m3WSL6QJQqA5/NMPn1Jos6PJ0kg2CtO93JlsQZL+DTeu3EJXXTKvPVMq6Yv
zF8YoaZIv2WypELcsy/VAwB3BH0HOcLaXVIdQA9LgqagZR88lao98YEcQnJVbXfx
bhW6B7lfLfznRssN+uld1zJ/gAFZmgCowMqWGpfctS5SqHxL+M39nYZKxxVyjudl
NfEoEqIQA+OIzt6Fwkz8U+zfLLS8ivicrqUX5QNbhPwsyvkfvUU//4flsnVPoAxS
cjnh1t79PobtJJAnvpRQAbWGNEuwYX66fLuMuIKz+8dwbvNj24VsMfpHFpg5ypN9
N1+Ac5DcETnDg2BKEcx6ROJhhmJsFxIUAbrvlFZ0NtoOPSJlK5U6X7BwQ0K4Jsry
7zpbS256jwjvsw2K54sTHRe07MwLMUIjTyUor+pH70uYqy12bcFx+MsoCBgwoKld
Me0ohzVaefCy/eKGQE0XSddqI/VD9PknjRWjRG3DmrQ5sP6lmiTg6J9sNMza+fP7
7GlgpIePN4EiaAIYYERFRHEUFrIRldSuiGxGi5Tojh9k1ZITkSkL8Eeod3Qtfltx
88prbkaXgJCfqXTIiQb3UsPVMo6HjeJvsdpU5rouFE148yGFc++ppAN/fkzzfcZ1
079pufI+9Hzh0bUySdM2mAefG5G2iIQgZF25jFRvMWtXClrx2WAxESvJ0iW0zVfi
rtoATmoTzKWuB6HKlePbfD5u/FDXQWb90vJcrNXT81hIp7/FO0fLa0VsKut0OURd
yKFGWuNxiBaja77zlvMZeX4FfliPdYz6UV6P492yDsJCB3DduzZTVX/fx0TVtBmV
/GbOtHS2Bf7zPzjD288UuYUlvSjPS9PqA5fTa2v80pwEKLt9lhRb6w/XLbwRTT37
myYzV0xZHniXNZcjg/XSCqMf5aB0YxCQT252vay+I8AMhGW+S6zWAAFnQDX5mrA3
mh0mDiiW4ZIM2+NssdhvYSk4zJdeEpQTHXa9t2R1xIniauPrgNn5ePLRm+P1+bw7
OK2JHo08Ix0ZbMUywjTx+QspRDRLCRgusAxA/CeRKLXr2KFZ6bNr5/WuwcIqaNMB
L6IHN44/8GG1WTPjA/Ri/ZiiF1F/w0o6d79/8ZmkDFbccjOZxREsOReYQ1NK5UxE
Lbu6YizL3YBC+aRTjF8a5o+tGLAnUOHdT/bWuVhoOzjhXQAq6OvK/A1Yl7rT0wGr
65sOFgLqIUaKL4H3LbLZBsD6j6cx2ObReB3PseMR7VKwW/LQ65EBAcqL5dQj0HHg
eeK5aZk3QLxNmnjT88RHSHL6HZpE5gJw4/pJaW8e4gZnAioWEoxKp3+YkpduH7yD
odIR2iHm1Grn86xIV18xpPhsAD66hmbWglVPJp69uLSS6YMXNylmU/iaPKyEPS0U
QmukpDo963HQHZD0BdtLcGADOTj5KK6hQsGos23gNQuRTAb+95GJ+KqOTUXxmm7X
l0MvfZx2HEGMV+L2vc6XvD6oeVMtCado09YO9XNFdgIk42s5n2VgAks4IKcBptka
VCInO+j/9rvhjqkpT9K0++uLyt7kRtxH2M/RkmGK0LdNge/YJ26P0Qq9Smcdnyig
elPakYM9FJUzcOqJm3aLYlZ+YSHnUZhsu1MmYnePolZxSAcBzcl/ISVtQpAnOrgK
8AqEsAL2Xx8ZIbYpokkfTV2mg+PIGieEtr4SZUItyNYsKuR2SJDd8J7H3wh7K3ct
Al6yFMrq/nnBZE9Q/mmIUw3C6VzrJtKtk9sOWStmc4BY1AZdWyhi+5OqBFwqwLJi
FXgcf2N/4kO2Yr7FZv+/7DShtUCTzjhws3Ut97t018lScOLjKYmA/HzldDz/Mzcx
Wi2WkaSmO5xFemm1NyMjNXTpSZuxmxYL4B2qp60UQ6vSJoP/kQPTnCdB45Ap1hGB
SafFBjDj3hLDQfHpgmEP9fXYePpqUOXWlMACQzGOk2BD3uVVKYWFuAHuIqE9Club
RuofoeVUAdSs+cHMZuUJREJzunExRqS9cSXee3VSLMMRJEgSz5uCGlFGRE7iQen5
huSfRtx09ZMvephjPLqISVVnACPntvybaB/pGyXaaclySwxQV57O4e1L5qxTuuZ8
SYKh/oBxX52sSiRBC1IwXfh1fKMOVXDCAFv0ZLAGmFjLWTahg3qNsnwVMnUzSgRA
2jezTnRQ8jRjK5jH+ZbondLXClyYyLzPDEXIrec975yWr1cqiMhmstKxXi44KnZ1
syEKRHAbzocHQIyKRWA38uoi/WR5Lo8xqYebIVAU+LxaR522SDze64vo1zzSvZRu
TnO+14xASRJ/AL/lUXxKksb+bpQU4+dQ5ZmHLqiifL5HE+duRz3jvhK1JqBS9UvC
kiowdD2Dk3twtq0IKhz9zkJzH9xdKVS3SSSpFaiq4l2yBkbVPa/yrsl7+v5sk/MB
uJ6De5CwxTEpJ1yTGLXC9utmZkaCJJdji9kdo02YdMfSqInKnBll9L3wryxPWX/g
Log3ZrvQgwXTLgtc59Ih3pby4OosPh2+NrZhWzGhBBjE40qvkLUeil4NZsWMHw3K
q57cQ15/4Ja5waB3OSwC057UvQZ8KwdDAazQmNnWt+itWhVqFyzslN7l5F4XFyEH
MYoFkYeDbYfjyd00zvvrwFy65DkbpuFNxkVpjJkQmgc9rLobCY1Hy/wY7WoruPTr
bS+75w+ew70BqhB0akazuHuP5L9MNB+0ZCIytyZd+4pvj6TJ2QnZWWf5Nj/PIw6g
gsCcmc4Bh/+zyDKoqAYu5/HRsyIMUwvfwSjxio+7LPiwNyRLPm82bKwtuKDxkeyO
S1Hvg9keiepflykFCbXeI/KG1Y0sfrxkR2ZGjCb9eWoEcLqp8jjdHw3fT7mqHJMG
p234xsN6nLnt3pMTJqCgmw80Lc3xRoe1NTLHy7HsenBN3sFxYgx3mSeEgcTM4QuZ
SnF9d4DXOUOhvttqDu1AT5BuHSSXpU7JuJhWQBC21p8RrMQeB2ZmBOW/AknT4l36
wNLHDPemAN3k6L8JxnghDlMHGeQRmksqEW7Koqjr1NJe/ANLxUAmlacuD1az1gtJ
HwYsOjwwg6Tb6P8hEKiswoLCyXCY/DYXPU+K6hKkDD8tHu9NQ76+28P6sicFPQZZ
MmDIwI1DmXexdoAszpMvA04WOLgWm7lpaDcUEBKyb20We2TX7ogmwp+HdlyjFxSw
L15roSpoFoZvedj4J2ag8lRqxCv7H4lrl1BJt9sxGK/9h/9bI7vXATaqywiI5ain
jc9945kN7yLp/vmAH4CLUy067lCw2iWSTs0OMtNLIgkeCjp1VpIPGtEVVPjs789/
fCE0Wfror9CcQuQ3PXQaIH33k6FMFbtifJ3BcXq+XxYtEb88vRonG/3Yxcm4xifh
ZH2Eso6wXJX4dLwQApcDGqG6fScobfVrx2NwPPqEyeUMau2tL4k4D6znl4EdQflg
brr0EtH1ayjnxnGPIrwfA5f1pAalKTslxQa/AOETe4t31+jDGQYm3p9e5qQ0ltSs
4m7bcuyMuxh2AbHmZDDtg++BDUpdey0k3i0fxWQSVxv1s224l/AjAUt/OyjEWZGB
rnsTzP5PRdmOyyGcjMSbMgso4Fe4oZPPIdJ1sd3kq/xBfO59LZNL8UhL/s5wZflj
avG+uzGi7w8L4VN9OF349tvS3I4vb63JAgmtKkpsTPP05AZ4Tju+cdRgr/ks8NQ6
OEOYe0qw44F0+2yQrGsamsYGG5GxBFXrWL/ywPX/yrxLb5Vkx8ALLXeYu7tfCpvh
L8+HRrifW9bbjIGQFCQr+9Ja1aEfs4spgb1GNuJqz+yHGLsPb/4u8v+9wcjSZAMI
g/pjf8ubhw7xDoeZkqWljiLfczfMevv8sDSjBeHtq3GJb8qC1FlIO3m81WvpDhI0
eZm7jLE97bWapM1Qugx126JS2dw/giSzxWCQ5mKGh+54njJMQwz3MNva0rUT6qDO
YEjzQOES9XqIJWTOybes8ETEZ/dU3mXwWeqwIT49RMC5Fb0vAKjD1WZXt1J5XHsI
KbtOg4c/5ke2BSN3pJK9UueZeJ597ijzNaoyG39ZEaiN9EVbVK6Q9NPsVS8t98DF
ZZKq4F7ena0Ppr0d0olHc3U+bsnWbQrhXQFjIr8J645Uy5Seg9Tz1LyLSKPqmaM2
b154W//5079140eXXrXiTzvLptxD+JciUvWdc+nJgRiDAmrdk72VPvh1m2wYaerq
/OXs1/anfZS500e2EHkPA5TVUbv9WMu2NeTAekhAOJcyGq+J8brc5nnBvstjiOCd
AuWXL6y0ShP7uzZ/KQDWXafH7z4VYmUVkqI/YV76mS+sf/GOFsfGQGX1spWepqv8
Kq/8P4CrdvZ9kphsB4oB8Wfsa6Dt/Y09XHXA4NASU6CNKJ+UerSTQEGWfd2zE+a0
sE2CsqqW9Ot/r+7YeMEUPQIy2mmBYtfcvS2bUgVdsKW4n+sBJWxv/iV/lwIvJ3nH
0izbFAZtkOcOefcQsvK7HaNwbNA/JzpBzoRIdLvcro1xukxZPOnrSKZM8ld1Ykov
ghAaBKnkkLY1/qgSf4TCpVoWcQK2bqXjS7PFcv8uybxu2TouN+9Zd+R64GftLbVt
g/pGtF2QXS7eudfHUKG66Sb/tazf34cMaXKpr2llwJJ9Qo7oVVylpAW0S1jE/wdo
+rY7tjsFvKEVVFQ3CpcXUIm0DdJmynjVN8cmbbbJL2/RpxpYbbaR/1GuUGY8Svsa
nGjJuCPayvlUib2gycbIl/yHC/cNh4cUy2Rh4pdGxJrXog4Fmo7ON+an4qBFzPZC
1h7L9ghL+dk1CyCWNPAg0x3r/4nxLp2S7yGNaIl7QrbX1Wf2zORCMea3RfO0ottA
vqmHmlBheauDFfqSXHbC2kRkMfhXRcV5IKM+MrqwaD1aOUjwuCdEMuNTTAHVTwYn
teNtqpiUH5k95BGTQAmHMKiTt3WC/3s6Ze4xK3ZWh/c+GpTmfscuNptDDGn9L6qe
CrwJIYzluBhuX5bdpWvJ/P/bXADcoa1ZL4ameslMOHSH6TaJdHAOfBgrhVBUgKU9
gMJ+L9v5zSI7ccXQFfrTzF/tOdsquuRNMjiNejW+jz6j6vI5EwcxxpWZkgrQMpBt
qUvhOwcryudSAIuhBlHwaA5nzJHIgvLjUUXATU8rhNsNREBZnNlJGQq0QyPaD9Nt
sDYZ/d5TbVJuORVIA20kQFp4ntQcYqJn8dpi8IzlbB/4/p/7x/pUW2imCggXjm5G
FvIIFI9VVbDGTP5SsBU0DxG8rEelubgDcprlNxgFJE/scVUQC+wgaR+raXjCdt0A
yHmnqjGFt99d9PeBl27kOoKDLzqRjE+muY2bjlQH0DbMDFNLPKjV8gAn5rnfihO4
lX/VDlOsheq+60wGw394WFThKXdcVcwLUYRK2Gfxd/fPkWLb/dyCcuHeVBv+hfcC
eyVdRolRdYL/1Plg2gxHC0LNtJ4nwlhoKJkqRH+VJfnzFfewu0Q7nrn/6S+Bvd5c
KSNtM1lgm+V96vMiis7gjn3WBJDu+Xv3Fiex22MbLz/6LikuqYX4X1chyqxOdGao
RIJ7K8/iaMYCu54+JFLeVsgZn6LogvE4s+nfyq7B8JlNHsbzgbRD8rWhRJY5U5J8
+81dwVQWiz6dNIy2hI5xuh59p8yWesaA2W/wtB9f6tn80sDILYHngl7MSHQ0zO2i
V0hh3jRLt2E+S2w8c34JieDmIt6ojWvyLjBLPpLfQqmdYbwq0u7tWq+spCR2QOfS
wtN4/amsaJL/0lRbQjPq7BcMmi190I4QEM+YK3JexJoEixiDKoMXQhDuCShXkwPw
FWXqbOUeSJe9ngM7FGvpEibWINu0vc1feuuizxgNoAxrXL7yazQpOxnUdLcKIBJ8
6OvEQiV75wRsquG1YF5l4ZQu+/wFqPp7BbVWOoIz4sQY26N2cx4iF/MTm2J9EXcZ
znEB2ybh7TCSM6j3XsWJ9JY4DzWMUxb1RRuUvq/R1AyuDpa5Skae7Wxx5FjlPRtk
US8xJVAvaxhPgXkfei7nmM6kj3ZHZBJ8gbif80PmJexbUcVnHw0I35d7UW012j9v
q6x8b/wTrXILXl5nPIrs4NmsVqkPqrVC+qFJOhQgFnCwzMaoHpvzXjH7QwJ4q4ZS
YERB+/oi0aa2pXeCksSf2ov1kZwP5sBt32kHyeK/zEjCOkzr8+y5lflftvlylfjT
IngfhfIQVZog7zZVxtedhRE2bkyh+MyTw1cLypguKcqOQ6CVybZVdJJ17js+bvGd
/KzW77r+g9si5Y7dURFmIognnZ9oaks3kpxyFZ8XWj01sUcz8qkaOodBjcW6GzvU
tsK/oK2Jj6cVEsHmXPXWmwTOSltrfzC6IZJFPcJvm7+Q7iFiBwnf5UFEmzWvDY2p
CZH6vSZiCO2o/wa8AK3+F2Dp60Mp2Fd4Rxfmpcu9cfAalI0yiWrfHAbbQBReh8Xs
9d8KpycytJuYfLpOpJWJev/jYoYl+J8siiaHT5oaUq1MfLgfqWscPtTccpE6SAU1
MSuJ06fK90FvbGyGVvoMLbQoTXQFTlYYx1paygxnQdbbKvERfjOITWeq++F92RyR
32U0G4RhXUEXAfTdCPi5j3o6O5qX9hEpWVZAjsyZoXPsqhYFpRPDn+Ml9CW5BgQp
gaPWgLsc4wXlw8nJpbJmwqjWGxz1leOMCrfkAinYtlL/9/72gB6RfCK7eXVR26ge
2BmAIDOQ5cYjLLme0NCYFygt7e7WaY74UAWE+mC6UyshhPjpsEPZH56knLvupWqQ
aJyROvl7MKiaxohdVWosMK56xG00I+wSLgygmAz+Ub8mlo3LbzBy6s3rLRdexXWA
DgjNdK8iZthVNDggbWm4073HaWQDhQ1MbP3rPleRNx/lrC+xd5DklGYtR1kqG/7h
vUWPdHX34S8D3R9UtJR8TuhqT3PDJgmvaR3/qhUcBWGT3wDMgjbkTjpN93viZ+6f
7fii+j7K+ipz4nQ8+qtrsZzCrBpGiQpLe+nRgxjYrjjaN9IcmzIPH40SAQjYsDyN
Tj7hx1yXkUMUoV2o+wM6VEfP9jJnQbCQCRBAzQWQEjOInzPBbRwUeTFyYNVKJm41
At9IY1rZLg8YrGUQvBwa5sgpU7vy/q8DL+tkkQTLwm5SV4lYk8gWC2v25Vn9uJ4j
LofpM9qeQIEbPEP11Uv/EuSe9fawBJMemoJ5DMbGOmNJ+y0Cbg+lzQsCKaDoi3Lc
hl4pPHNPj8E4y6bxC7cXwxnwm/6blCz0AHSP5r/x6D+rk3sxGyHs/cF5Ed5KvY85
3m0RMr34Wi/bAe1Mt7TeoLCwV9ZZTJdyMFAMSVg1aJic5zyyaB7qg0776FJZh/jq
AkZermqz30EQ0T5K4BLDXn3hpK65GMmVQY9Z6OmUc0SEgoMxMXIlevA+PiB1ryeO
rxs89gKzsI5Q+R6vUiydDl7L/gWSI+aaIjM1BPHeIh3MygSP0KkKBnQvZ9OkFU0W
61xnnROByPrAllkHKWTTwSIVgwzgmimXqr1YZgsgfsVI7k6a6bFODIdIrG0n1Dck
Zdjcf/kq09+ngRFrKxtn2Xs3TEGzQBgReTO/DZFIyUV1uuSPlglmnm8z4v0ZIBxu
sxcLKFskPTAlig4jHRuBHSHAq9qyi34CaOUFVaKF1fNojp4amoG83S5sJNrwiUTB
xPFznV/10IM2GSoGIKXnFePjVSd85J9fHq+3MIn0gf3RGef2IyolkgTuEb49qv8T
B0BPczK2cNHBmqbZ4mg03hqPsdBh59brB96rC2jCsh50t1ME215Ea1jXhsQrbEbC
Ux8LQPjMQNAeThAHe5B65ai0vPZ/BJWlCZxYNSJCyPrAa9Lk49GF1AIeyUOx58PW
kOs+nWUQBRwtcOK0Jr/hUDR9tlo7+RiQNJkP7m9j8cQiJw+129XZZulnHxCNN58E
32JU1bc7TYuPRFik/thQ9OZnRO+eXWDNTdrS6cYwv9/+ccBeFwG97+PBvnY1gEIN
yqPtk2ssr105FGSoJZuy+Xl4XAXx568d1OUNLBt5pDSiM2CDeBTs/elEZLt6PHnU
Zkx3Qchk7cfMdqPVxP+MOjTBnxuobR7VGQzrJ20jgVEWnnfgv/Lx5bH/nl6xoINb
jxzcUdNZKp0eeez5aPAlbyUlUv7ePawcWgwNe8MMKLxxKgN9aEGItqsXv0h94Tz7
aP0UMYcNBKZVbidBBvSjS+8jSHcrs5bDJg6+YbVuq/wDQQxIIpUFaKQhbW7NupE9
W+G+oSZPWTOYhpT44QCwmalo8IcKTo/uHmiOAMVptxHgGXsLAczsj70/Koc8xCtx
yv7/phngP38Qy+XGWb2wPWVm30btEmmcjPrWSxOveLuBwHEUPG2LIK1mg4rQRXLC
P/8Ma49hdeHDSkU1DvK9BDUObZ//FBjfArpMPw9hxQwOletlO2K5eNI+6sboPhbI
roXQXoTwBWehbrrREeM+znc/HJer51vcYlox2JZgOFZq5NOW7E3Rxjg8XzizFZNh
5kWcvSwW333GxMxGPEaW+BL7yPWAv1eYcftc0m+vy0a1S7tDl2Piogdq0IbpYE92
6Am+nbadc1H20PZtq6TNqcE52Lacze9BJSsj57T4EvfYn2zjeu7Zj5CX9gM9Z8AQ
qd/4Id8axYyS8pfwaC+aFmEYEJfUdkpskbLU/XJAbJVhTkPuWKuaGMwKxRjb43cM
x/sY8q+KW3zVN18rxcaHNiPj6eVfYLYAdlZSMgvtXkpBpK9/RvVv+MgIw3r8cIOa
d9JoQ9LHmKTrZNIJ+2W4Y7RCcFUuUrJXyV/eKcZY2MsEWNFL5qhtwSNKEEYyl8Eg
L6ko/RNdSzAGwHCF0ixB1GGMQH3gIeE2Al9aKFCsfJzzgl1EJpBKDWRaNFtOpqDS
/Oa58TRFoare2seuLDitOzlNjz+TOfDBgO7M20sZjLJsPIDjhCQ9OouPm9jIsO+m
r7IF2eU1QwW7hSGb4f/xUhO6z/yrFE803G0Xqeps5cQ0XdhoAtFq38TAkiGEw2sR
/t8fSVmqseTMraDWZSSFh/Cm8SW8K6kOoper1+UcLKNdTCDfanj5GqPParsqNDca
euzrPsEB+SblPUzhEQCFv6ukPC1WhY66zDhdj/xrTM0GDo1P5tE92dJ8x0rIDVwO
vkDTglVC9AD3bNri5tjP9vgJPxJNOYrI+HJQfKxdx08oIEGEx7DTws309JMttbDb
5JK20xYNOaJP36NxHP1Rl2yPgKQLfl3Vs9q5+LCsel3ct/QdpL23KuIgSMDHfjc3
aEHhmrBpgG0+Jzt6CN50z2tx2HYhy5eikXc7GE6TNwG660bFaDpD0WJRnJfmLglz
f70A10jUZoNXQnjCFXZbIUN+vOT/SghiJUNsYaKHkKWqckc5aPh6u0y2xzJEhKrv
0V5jtS4G8mSgidniazvfOoDjOuZUfcwBCKka7EvUjtOVuKsQCB00gcq3q+2P3KBr
qS/uF+dcIReP8XWlVnz//pamp9ccnJ9u3g2Y5EnzzMeBEM+Uu+MCcorbxqkDP1iu
IKoEaR8uJWNlJlta0WsXqgIXaDIKnpwsBldaln/TUumbxghUe6b+yWkMB+rV5f3+
/mv0VlCgbKMg+sQ/pZTo2X8tIqFBr2LEc8s54jdpCkQKUSxT30gqunh8naeJ6Fyn
Sh30RiuSkYZG17cJNTthOoBwGJpyuBWpPKfNlrJT+ZkwjQ98D7QzYjF7bXj8vk03
kwVQXzOYd84i5Vp+GqP3JnOQWtj5qZPBTd9S6pnNBPuwSLC/s6r2ZOuuavy+T5hx
tzCf2QJCF5qQtAgz9sB0reC9VbObyi+U7lZY4byTLc+QUh8LVMDcOEuHSgnOwpxS
TDFmAaCg+k2yDe4JPp3O7LO4IvFesj/nex9+7BZHPUjIN/xlFawDtWa/LqRT+1xR
vEn3idIWje4pZF1phBNA0AmZCsuQEGHhHytBCeqZHSkgV7qrdECcFPoxFbE/cmO1
ZiVLK+HInHI0hjPLe1kZhZuZE5Le0q4XS1sgqp9Qc6HeyGKfIEBmIBlYYFp+2F4p
oOz3P4tn07MIv+1ohizs5our8MH4WzEryYcDO/fE/qJunz2b7dUVGmfTtIzukPfY
aOoU1f5aueQ5jW+Lwgi7WnvxtjjnQ3NFxSJ/aI41hARjxFFcTSp/9fsrW5w9cLRM
vZKeWAZFWMLfnAhwd+hyVZQwRGW9s7Y9GEkpskNVLrTwh2awMNEvZDPmNVyi/w4a
Pnc1xAQ8TV4JKisSYpNnQEUzGFjcnOABwB6tJ0qsKvgQIF5CALKlwg9CsSNfALqg
Uw0cZPitvOnetoXAfXyZy/sJVU9MQR3EtFFkrUiQq4UaevOp4WTerYhkwZ8uLeND
0rogAUdSZ4hlPtx1n+EZUAv1sPJO+HBlgogOCkKSShuLmv2z9YrRIdrIfU7Li4Uq
nNkaYlrl8dLH7Hmm0/KYrdV68XURKm5U5YbnKNvtkwfLZxgjIaF2iIzTlEVz5kaR
wrgKJLb0n1c09UsbJeHCz0uA/JzpLGyLUoc0pwWz534Puu2OFKK3toZybRxrseqp
Yy/gkd64faXuEkcA1YyBAG/NTFwl+22TNrp59p5e/PvCDAcS0tXnycnO9scBaHGl
lWKyoZ2pQYn02rAIaXkyi1F/pj7ZqvurNajj6mf4yAK2wN2nPXuyCtKCJsd2KF2s
dCescPALaGm29PtlpzxRyp7wbpOWPzcgU8JB+YstjtYl2g7GsCqJ4j7jcRxGoUF7
GgnfwDJcWcXqn/scWAAodhgQmkejBBiVJ5/TgHuZIcygOrH85CBImJDHaTjvNZN9
Xks1CAjsKpZnaZqV6zb2MqP+axP+9TdbJ2G20d5hEy99s2XlLGyqc8tQjT+QYITE
/qMraJjjO/Z6q+guPB0RGizLN3Jee8WHsqP/tXYiBE9u6PwHCLowOQeIdO9TbU/e
WqE7THWyYmtgUIkhkuOsUIbecG3Re5EAfdrNZqd+1ACEbc1RlaUoJqFTABLBaa7Z
gO9/IeEzK81cUSSVd0RGeJfnhqpBQafFOS5wCWaf9Yl8ErPPN/wpDKNtUllJiQej
J6sIhhuGj30pbhHtmJRwxJvpe1UuMlmagk3Ch/eDcOm12n/N9W/xcsM+InUVf9kc
Jcjf43mut9DpZalbzUmrc4ck6eQILFtyXrq3ZasJliAm6txU0BeLDgGTp0yrBEi1
tHMco6l8KI38eAaG6z4FPJdWPXT5Aj5Z2boh9v9Vbr/Wm0DQXjWDVOJPJF471EEv
PFLZ/uIivEFXQofLg9iHRa1ibVWe+Jfd0qEvg7dIooC0ywR+oWGbx7B2WF2AhH8E
TzM2mIKBvh89qJ5guNrgTs63uTSZXnBxbontfprzHEImvsaYD7mu7A1P3ArPWHEL
+pOLxnPvIiuERMfuyS/w1gRT27nLM1qM/3PXdM9jZ1bLm4STjKOSd48vhkSSun1x
yDW8PP+QHq65WszZxBAtqnJC5yCk8HgXBibdRESc99Xl1ybMay9+urWGWweh+BEL
p4/VdqJPYqi2ihtr1RGyRhkHbzAkZ3bkHRYbjgut9Jg80U5FNJ7IvDxGjo+rwXt3
8/s9YpmtJQvc+oa0Hp1Xc3244Sk8y7Uqc1gULvQT2ohLgvoHu3gth0CsMJNFxqBu
mK4S70AWWO198b4TT/f6QrunsfHRaX2Zidc6YYCNth5dAIAI8zG0ghWRk1rpC6gy
ELTUZ2XAf7WRnCq6ancN3PJuHIzu5NAemM7pxd3/82BRVkiy3FTGYup4AqKk+BD7
0rl1pygo2QixuSJM9PlUXPzkNmswLvOqrC247P5lxpwNMjjow6P2Rqu0dpjRnPu6
Oi0tfjhimhd0NiOg/JD8aSvEV0Qo+FBUUAZq/hBmtAJVz/4w1rhc44HlEjz3b8Uf
zQ+Va1BOx/a6TInqXzhN0HFeLQsXVkAymWKT7rEtWOZ4I2L96FhbrNhbWIOY4gXD
wpb+PofEGDPMMb7LaKzSeNIKpecDDgDpSWDR4sWRXA7mmxMEVRZ5EfnxjMmKxoYG
+ETI1O4+pgltTqEvJF61UO7rWHsbjjvwHITSwg/RQD2qH0D6ettRzWdjDoGx46Q4
cnqJ9aEMtNVCzYILzL4M1W/uYtgT+niXz9iWaHH3B08z1ovBJ/BP3kCtW26FbXVy
rkfO8mjVQRLwNnyn7OKxm0O7IqmsujilNiz65H1RX4oss/0y3+y53No44CGxEKxs
CALhx/aI4FojQiD+FMdjDhcWJ6X3aEDCiHRk3eMNbHv0yme7l8brflYUsJjndaTL
8SP1BUop5KZuIddmZHL/WYNje8W83iYMDe5kt0SEowh38NjYU+dzFWBPSuroEOsB
DOd/5k5ytDD8zEV5fK90lyMK6AtEeV8Sn9tRw0Gn47VQcPUvTPKC+fXp5DAh4TR8
iRMTzxom8h5AbONGVbtoCnS5Iuh22iBS7G3QLYatUd/F86Ffx7keGTmkjUXAhjJL
RUkeWJpkmmcp6tIKvn9dCn0eHH65BtiXxktyKqQJYYpilCqCiOgbNbjayyREHajx
GEW658PGwZ6i7MTXyut4TpVGotbgd2J//bLSUI1cc1Pmezk/+IMrnR0cdnNcPDbv
EZpzbyHUamMEA3ydYBVsDGp06VAajgVhWJPR1zOfXRW8j8Y+6T6kunpHvfBnWEbv
6E5dTuEuJr8Lfgg0HHnC6pyz+P/Ywd1z9SQIqxSF7r3exPT5shXJI1S0TaaXhJ5N
8XVGsVdprgisCODMMSImw77L8Glzv6/GLRf6z4p+kdup2qj8Hlq2M77Y6rO7mFXT
DSH7iFkto8o5I6aC9KnNtfvCNblck/phm40giPYE5unz/L6gIV4JnxkCNkTDpWLj
RyJRbs5F26J+NglPf7kwCR8J1e1xNU4Zr4FQ4OuT/lsdu0ypPj/bilQFAEcXSTi9
tkI6zihR+t/Lz3mrG+pmNSPSrYlgzHyTgeS5GLCJ0KcIAmnluNjCy69Rg2av/x1j
SONvMYmiKL7bCLir1L9/Hn4UkRQkzHfPPr2b2UOW6hQcHeDXwM90MUWu9AH/RBfb
iMY7d6xs+bu0qb9GJLPF32Dl06E6ZxembhysC9WawwGgZaUQfC9ExKrfN6KKpnFh
OSh0GpQ+v5LPG4Mq6Ztky3DtglTzIV7pgBXOnPhWrqVhns+zeQyrgKFxdyTO1Jq8
z9VUSsmUemWvd730gSM6GyUgP6PZA0pmeARfCQKoW7IEVsN6VdsLsTOpqVbR8HIv
XKL4E5Y+NDP/Z07JluibB9lvCada7kXptpQiyts7qCrA4GTYnGyx4RKufWJmprdP
5prPZV8KS5GBv0kw5CEXAwCHrhgu6Gfnzar4CZdTSMQ1+3RQaCuRQ6GrZAtK2ngu
71AV6x6AtQ50Zx5ZHhUAZ/VUU094U55+TWbv3ReX5yn5g5ZSe4W0HJpKmwrxmVU9
+ib0jPj7r3hNHGMCatYx+MA3LPvd1x+TqTTAkzaHYm7xbBZWOcfMELYuRSkxtCo/
RHBT9bpbrCntL6gtNcTlg1TC4nEkqzGh/pvIDXQin8rnUKgO/7WR28YqGnHY5uyb
/22t6QD9AGpdDvwyiNqP/aNI5nLNWxfmYzYoP+I46BH1yrZxOl0w9jPuhmD61z25
QKu8W8oU71a3RVtW1xkcB3X0fsbR6xeo0/i7h+EtsauNj50KL0bFlpnjS7Z1TduF
70cT/iAbmmDQbQUaFNwrzQ7DRlbsMNIgRRfXijjTFIx43RhzU0NegUwmj2Hd/bdd
+RWbKDCFciaCVKDH3cBU/GgYKmGtHMD4vllVnW6OkSU0oSUjMrFi+UwtEyE7wbXt
gWLxFxGdqcPi8gFJ+8RrxUV1BSnmKrnJ3ZA7a/iEESj77ou5HGFNuprrkXkne2R8
VK8+TpkiWtsmHvmG04ONUiUWgDbBv/FU5UulABCZ167eko90dEOPcj+9xKT+2u0k
dfR+X5CQN8jW79NmVNdzJbjNF3AwuqMMiv0t1o1JBgPc0zsT9NrpPep5VMesRE0B
nFwRSOrTTl0e+pVM9mmW6qmihh//2Smy+/a55PEghqIsem4LV8QmBnLi7ykf6N/Y
9gU95bqCeG1i56Epf8UCTZ1leoDIKYGbp05lMNIJv7NzyDuyQ5QZhhhtIsq+O4Nl
QXl8qzbcy+lMq33P/hPPwyYKDV2WG7J+gLt3HMfs1bmf2waJnB2shx/er0qBO4Kx
6W3XLvVQyt0Nq9fZ3D3nwC3pI4jCZAE5TRoW8terq2sflPJe/piUaAiEWR8qYfoG
ZAylgv+cBhR3melWFBR9nVGAVgVY2d4Hhz5zI0cPVh50pWjn4bk3wOYV2ao+0Bcj
AJOkkLKl/EN6uxnv3kRyQEhg2y3x+hL8Fbl37L30l3+Op8rY6qBzE9dvbimhJIPA
63Ff3rq3lrxgGeE37KI3LFaE98iLT+IKf1SH5SDqTa1BtR2lA/iOU8dGi8t9AIlK
k9jf4/YE6L0yK42HT9xgWGiFbyjLySA8nwo0VvtbjBIi0LQwnDhITXvQWRiqvS+l
qtOO6yO/evhRgMKoHRcnhdLVCwKqsJzmkyTjct2hZaTMOMsRQekepZq/Z9LBQCbx
ip5VC/qClOvti7Y9IZb4AX13N+UJi5vtmiqGIUqqqwk5hcSWYumlGm7eZMJKov4b
srZHjDV74+S8URgWVbtOue2/Ssx1C7kKrGPjpQJ004qcDmMfaBJdqOOjf2ZmpkUw
mWWpe62ypYIP7hn2H7MmaW+A06Cdh7EhsBi/xqwXxvJIvS1mDJBeuUWQ9ZWBfSQ6
F3B3uH2MRud0khSXo1mHwLP8q7Ug/51h00K9pJ8nr+DNaskx9egNXHGotaLvDYZi
HEfk8+DB7jR5XkPbkJHJ42gKZ6MImKl/sKYa6wlSsE5zoHt12WjoiRusMRFeeZj7
8/vFVXv5daT7PhDnXAzRyjZ2C/WyfVWeR5pZRUJa3JcDit2h8tPqRz8jTwY27115
55DkS/uWmJ+y2PeXQG+3sN++HvJMfgmy+E54lKzLkNnUWPYEYSWqWdo1JyH+d4xg
MIqN/Q0981Cxu4s1BbavWhbGBG5oNYpgfzBbj/rfWqsCtqVSihgacjDDTKdpYToS
nN8wricBRUL7wiu40W9TvIzG5GnfTEMBdvcoa3OFjtetKXGrBUZR/VIARiMo3QWZ
+jJdHrlLum/SUZBb4mzJzpBW/FKyULNSmksOjp+qrx1FKrbo8nHe9yVFtTFjX9NJ
HIntRyRqOST03ySkH/EgVg9BqZ5w5VKIIAO+9YBaSgRzlwMWMoETc4gBM5+j09sl
5Mi+nwa7K0n65OfQseV3WOP60cJkfOlnbKraByq2DbpRH9teLxnVuKfahIkgVp9h
2Gc+ZGhqeXhrofBKmnz6xFlcKUY05rkObrwVDPf5mJMK21kZQxcuP41m6sGtwS/t
mtj7hKWd7Nfptugr0o8KlybxoG3HVwIiHUNWs99WYeHpN1onc3afsqPpeK0KPbFt
58SACK+olcOgw988e7E9R65LqoKXvKm5f1/AkvD/ptuty4Qn5afcXpG+shZsbemg
bs7wcqdCNqsQNrBtGQXx8alymqOxUmkAe9ONn5VxSd8W1pgSs7O2FVbzUSo6R1iR
MtsKIJiWHpjSMwizkXnCHc8X0MsQqY/g6wOJ15v/F2acHeXs1+S1KWgBuJ0rHl5K
IoXpM0BYBZVs0dEzezcs1tcLyTiqM8UGjv3MeuRBR02JY2KLBkW65ESTEi4VeJEd
0f/BUXCLFNZCUxRo1bxQK+iUANEMHMGtQSZPB1Oxz0gvkRwxQvybmEa3nThBIMJ8
Wr6IOaVQY30m0NBoY1o+kbwWrVthy8NBZ3qA2RGK15prcXNSYPw02NymTbCDDalp
78GzlnvMtAbze1snSVrGHa6CWnRewlv5GWsvns8ec03HHO1PXefN2nOdjOqbNIB7
/+raqUZvDupSkrDGrseSmu/eu1tHGXzjFdJO1/LjZDCHT3Qq8KwKLVTh/KMf6zNW
kL0Hcd1ltNl8jhz0GpTCgbHLNnaT+PRcak6Wb0XkCL+JROQGx69gOoSJKvYI0ait
i1xYlfkiLcrPy3nWPSxjMEO7+U9h/1v3n17kErw2Br+0z1OYxoVSkEd67/Sl/HY0
eNFLDnjebuzCRMCLAU2g5+PX3MtbqOFad07YXAqRD1SRFc7zoePm7IiyW4vM3ah2
twVeO9nJtD0OjIDJtKpSgpTJui5uLDD/8YPdc981mDTShtQiqTon/s6ULSfivR5L
EKLutO32KFOzqVNdcZDyILrBGwMjXX/YZtCOIBMGHm2fxumwzPXUQ+5R05kJxNe5
lWd2yIQdRj4dqgRA0aURqTYcdlK2R+swII+6UYJ0rh1HYrKirvWfrjf95oZzXlf/
lvwcTvfPhqul8W95HslSAifDw0sVXUGQ9iZw97pjDyOUo6RlXRVE6Wq+uwe1k4pH
oqQu7Zzl6Dklvd9mQqt6gnQmNCRU3eQWtlEtTjgo9UTosLvYUOTA1QDzUu/L9keF
pvV1lNU3rQMsz3KySw/uBqCmvjz699PP/BqIp/6fjZiCktlM2mKx0nnm+vxzBjeS
2N9hZ0j0oOpUTGaX/8FAm/fnrfc5gVBy1qChmpaUDsCYmM64ruRsnmLvzNkex05P
RdqGaipfeM7x5pD5dZTMzRLXDfZZIlmhhr81DP/WXWgvOqafiBqqSyOwuruOdl0t
ibuW/hkxewwEtea2JM1Ynbc7x8XZ4J4UruiRDDW/XX1Ughw59BYtOZ/70469Men5
JkDsJAWRC+neM0C/hYc5SFTxCD366cJVeFq7/YygMY0/2lMoXn5/2rb7PDTQtLrC
KMkbz+dSlOc7GOx4fphSy94+r2rRi9T5oGrbDbS2jJyB8QqJSfz293lvWeFUkG+v
TFDxXmjNYFdeyspeU+pKoCMPY6Fb7XEz+FKgB7SiYu8WNnvjnxeUFh/Bh3ZJZD2F
GgzcGKTzeRMNp8ft0HKdkI6d9Lf2ADNuvzMSfbxNe2yqMcCjeFBRe61niK8StOeS
d9g4JMtulXCvdh67iLE8NaJzg/KIwi1rdAqsZjpIrARKAOIhDepygJuWbaypG6ms
t2neBVBO34FQq49M24to6ayClZZOhNnCSJtCFbJKGbjVaNHe42aNArHIeR3qPrln
DZvc7g6yWL2zZGo69BUDswblNtLHtqRV8XCvXTkS6v977WaUYvtgruxOErlpWREN
o/n8eNiv49dnYQ5hxX0MmB3GVnnlQEEXiOu3Sb1T/Gd/rZP9sBhDQAFmQRAMUdzW
pPoFGpUUxuMPN7Vtg5CeY7YDB3fSPz2WPm8NXl429e6Z2f5B1SSCRkpqCxfyDfaN
bQmgnpxfcBPSwj1XuMH+o11Dzr8Z0u0F1XkN4pzIppJIVlqgheyab5iAT0TbJt2L
khbME6HFYZGK8DqLkjIO/LhTftqjgBlrayA+eGHaTdbeOFz3jvydyKqMrCju3rc3
Omse5dfEsBlUSiVvSZJcZiFvpzEbg8H0H34xRA/j0n3Gcqu+FX4sPwoPGHs0KOns
8qvKLIghzlxvBa7zRCjF+OS3bDOrWxmp83PPhrgL33dfzMMEW7nSFgLlIg4OFRwF
P0lqdWnc0W8sRbvcyulVcc6sMj8o+LY4k6DldIgmAOKHhBAlS0TiGpN9HjXVxhsU
cg9iXxYyRdBbnHa1DWfD70Y02ZZ7t8eEzYaNQfT7pXntvk4FvOlTNACv/QxbnGV3
q1VvZ+zFpRqihj2W0CtBsi/or+eP66QqWLv+BKCBpigEwcQqLSBZypazVZSiE2ai
q7d4iPF9XCGGl8VYQOEcnQE3cMopo2oHBqPdywwlD7DMk9OpEQSM3USBl3mO7c7w
Rviv4oDjuqCQxBYqqLDKzjHfJqFU5SNJh1D9XNnaDeksYRyXIcAxdHGgYLuPNAWh
CqhL/j/VFhThmwcqs9x9bb0YAzcKaBSya41feVdVQKS14eeNlz904kGQOOcDhHyO
8L2ix/xlrTkX1IscjdUKc6nUI+LZKuerYAwHDFq6Ada8LIt6uIugC2+oEA4KaKSK
KDbmp/ecdiIeXgKmxeqOcSnuvKKoQ9dhRd+388a11mY8Ztbmz9AFXiaF4CILnThz
T2FwLsHOWMyJxXnM7cpQDef4RgvO9jj+KW3AgIdaTlbGnjhD3Hhqos0qg7AFcLy/
cI9N+adBmMp/nlg83A1uS33uePRP2ZB5UxKe4q88glcXmWBpC1K2K/4avAGuBQI1
+nIl+rW2JwnUcv2muq7nJeevgr77VTalzLZj1BsKc9Q0GDc4HFw3TZZRSWv+6kYt
cFf1puhwRe5W4fLZZe8jTNTh7pnVfhjIrp+uWY16smoDFR7IQGhY83LedMJIhkEV
rCCYljCQ53ihv0mSvg8s7pBH64qQm6l/ae/Gu9ksF9VWaaeGSybLOz4es/Hxm9ee
9d2ZI83ifN8Q6vv4yW43d4pyLxUjDYEaoDnTyuQD6WPpZA3023Ic/Sb1wHGhmnrc
Ex6ZlXoJIOrVgUip+VeUTUUyiNA4e8KufDSQKybRGvoB4UY9wwNGmd7H0WTnjNVQ
qWDt4nH3nIvwZAEyfSIq5Dt0ii9+LJIfSDBZUhTp2SANVUtuYfb6ntuWCDiEFk51
LeczzMEgmPojKDYqdIUM9DQifAUodu/0SnLj6tk76eP9X//32opI2XdQkihnf2SZ
EFuJzyA7u7U31Wmb86mrPOiJ+wYQ2EDBeWdBCTE8HcQwb+/7/ga+Dohg2Rrq/Jwp
8ywjqw2fE/dHQLJx0D5RgASlwlrHQu1Z049UCyv7CaAGs3Dmc7wHodTk4kdFXej2
18E+z8vx8C6hdXm0V7DHwCSicfCE1J3mt/11nx010HOV3llYGKaZEujp9TuzWY2V
KTlE1fDzD1lUapYF7YxPCkASOdErnkR4TYDgUG3IplTsoYWDjCfahHjNnf579SIE
d1JMyav4vT0ziEH3pBRhfD+mK/HGHuDLbhfeEOKxPyjWJZVzZzmur/jk+H9es0IE
V0C5CkUx5+Ibq1V9Ap9PHi5q4nVxs3bzDJb1AL7lpx361XXQxwvtVaM1E5wNlJaD
jAEURmdwhcjoiEnr1hlgP1X/ugymmjmiRHgSrDm2ccA7cUQXd52h1KOXYA3NDEbq
zfmXMPt4z/xuCeFymiF1W+0c2HtFTSs8k74ZGHPmG1nPk0UMvN2GInAhat7DW4Pt
a5ORnGZE0ncaa6sD7A5XRhrCNIA5oVRb+0W+jzsvvpBooyyQgkcNjoX9UKqTC/v7
Q7RuhLHEfO8wiISH+ISRJh2joMgwrzALjduN6yDfbtNYDn6O7798sRu7WUN7EzYV
FlQIxuyGeGU/Gt66JegTfUCq3zJMh6hQ/l0y2TCN+SpePgwD8AGwbUwtRY8BILbt
lahEWU5ecBNfq9D+p6VowONPOz9fqig2YrMSHJp2axAc/ixgjtvO3GySl/VEd8zp
E9FHqFRWnDNzmmeg3AthQGp1ZSkyKGIt1MC/Mw7uTlBz0XNIFxJ1lJ+5o6H+SqIx
RMJUc0eNhDHCDqYX2cOKWAVd4Qox86eYtGoeVXifl3Li4ncvA82w2RfVtny4md6B
axOcBlb7iRpKKtvh6c1YNwEiKf6Ntc3iSJz54BUmUeiwMBGf55GXS9NgDaWouC9a
+899OBwEhiihbIuKpoUlsmgRUqvVhrs+hrkBmJb2+n2g6eagByCZMtPx7y0dkh/F
TH9xwdN5SF13Tln+TbEAmXZ8Qg5EVlaP8U8C6yILLRbxVDPD5Hh58uF3oirhyiGi
XpjEj8HurkQN5oDvPXg2k/4SoKGOYKXEBcXRRYRg76lbJfCjy2LmvNu/y/eWpV7Q
IYXDh2YftUy4+UPZvRMpMYzuCpq+XAXb+sDeZkV+056T5MDdzcQu5B7ayqWFoY6a
ZaLWrmN+K0Xk78hrwQD4sRxAvTHLyI1UIn45e6cHbGCJ1m8qwiKQU3ECdQ62GI9y
QHqPu/JwmeD7tJQ2izxWnfD7Y4uOOZNQeaq2TzLllC1q2VKuoeKeRr56DwGaqCuh
y+Jgk6Jq7pfSvrmciJND803bNhISAQ9BlOOLkBty/r2xddCMlvG5zuyAUAUMmA/z
fdv1CzfqOBnVPLC1pMmJqnobtKYrcVKOKF5xS6w/L0/EZ+FGrA8AIujxMHaWKIOS
qU6DPGaNxGTNAcAlrh/ZIGPQ3A/rU9j/MWZir6L/XqUcaxNCsdkprrV3VAJN/2U2
GSj74nurliLDMQ2gFJGWjG2Yk9JF159cCJCQ3abkGCJ7HysO0tkfV3+k7CFwjp1z
4DZNFFqQcsYagilH1HOKwR8pmMcshHobiTA8eQkKpPTroIeD6WNLQZzTe6f1XXVs
YM9UOBHJxfTw0Lu77he9Jb+MN74emadkioqsmCD1eszd46Je3Xdar8gzx5BetxNz
2baYB/xmCPFGu/QSl+r7f02jqkT5Yns+TF4BcmmhND4Y98GFQ2SMORrM9LH8L8E5
INUrR8B4hmB/u+7jR95Olx6BnwsB1anCxDcWTI/iZcMZWyiP4XvrTPqQDwNOCf0y
+o8B62ZHxNmjsByvgn9ebqUBb88yzpUNEFukRVN7LXHhp9cTZUJ/63xqWTTy97vz
FV21P0gIBe9WdV4I38YhRoLQEuGUGi2tEEWO+kI185g+sq1+GdAKf1R1RhDSykyD
qAMWHEyokOjhJben4cyJrxsNlZOodSXOOPt3+4vp3IItsdIwoX8ECUpPN2YLgtAc
zDhMqipi5hd3p0ZtrOk46E9Xh3GrYa0pa93DtCWKTmAN7l0fI8l08S7oLn6y2dxC
T7nAdoYY8TxDgqX7C94fO3FrYsc+TVIiA40FAqppLYQWyT2OTLbwQvAN99acLPiO
UB3ttbVqhFxY/5aIPJ353HfmGc5yyVD1vvlln12MbHh6UKVAz/CLgSgAHBI5t1qn
I9ksjFPMZ1dbJc9YyeqhSdVWw4AIBjo6xS+5/S6cQ7GirdRuSIM3a7a8Od9OJpeN
tBRwhkJfjxPFxjbqfa1Q1+TJxXp+UUz8qaxwWWnIm5vkcPFgNRHjkOuEWFSWRHVz
poW4VjxVtHKEZQwLy5c1D+KlsdB34ikHnWT0TkyhCiOiWYZ6CaalArcwZMRJg9l7
JjMpoML0fuzuZhJFHVBYUinKhxZbZrEpRcvFIVWbdaCTBDq8qshD2vywPFOxbL+s
uL6mlzisyDThSbrncXGL4Q4FRigOlbTlPzA2ETcTwmIjv8m08ZgMt0jKFUD0VxIU
szcLEDltkwSts2ncwMuCi+DL3z56myfeAUhyaLN6ARbMu1/rlYKLeDXHv0WorGkI
nX71XCnFTMqOzYrkrahF9V0CMiEgd3SusP5Tml496yIT9c6ID0SRHTd9bsNjxWq4
TYr/dsFYEzee2aTEkeV/37qrbT9yrAkcyyKvxBuLxscsrSaj25gQdYQUtNY2Xqww
TDCcTB9fBFWLfR+5Oa2pFX0msC8gYlEZEnfqsD11YJAGaFh3Et+uh91QzCwD21ZI
YvE5H7NsMm5KoR+hfajRZ+NUzL/+0waIrqRBihULcHhNlwY5ehwoR5gLUWRJeWKn
iedgaRrgHl/PO8weY3aYpJVl9fCDmcLMdN+5ccr5Dg4UcLAvlo3cEzASKinU7xYw
7ttju847uEEMlINPupuTh4adwzyc8I5COcZKanOHg7VKVian19PowBlSTI8SJ379
onV9QjlppweErg0u6xs1QSl/2n7obrq511b34WjpEee5OWid7og61n1P0jzXiOJl
JmkGO3MAswcrSmmH7XIgwfWl9Ppv7rciFJnZPNxtNPFKsscu1mNAX86Ag9Zb4VW/
WpYijkmaf08+1piHCSJsWrLKmjsw/B8AAck/oLA0cN4ACQ3GgV7qgPBfzJEeySoO
XYD8noQdgqJYf2VhStmvSm6AtscedMhBagmmfRgZkqmkeJCvc8M7r2O3JHUbv11J
4pI+RI39hyu2XXOcDO9kPXFstzUqoi5GPJymJZOzLe9+axqOEPlWj5O4yaSUpdI/
h5qRxzteXLKIRK+25xjgmUNtYX1WGBl5lbAuxT2xZovz2OF1x0weqkAD6OtgaGwM
p/QajtZZqfweWW0XCgI2pOrcBqahaxZmAcNbpRwc80xUco6P1GchH3zoYUT6nSTZ
oTn4X70d50lRCA7NpFyLqManx2n9FU7BSvVWxyVp9jTjmaVZ4e41iadPbGYbEw0h
wZ9h0Ye9vJq1NNU72GSJU55s+ePflYMNXqFxsjXXKH/brdgySS/4fm1GH/tAtuo9
RGg/JhWoG4or9wrxQN6Yc3jHAdRVqt1+r0Nz8Ib5XWpxVna+coGOjrbHWPObkrjv
qdMPDP0BeU0YM/K7vkPYDU9rr/D6t9vbzWY+Jf+O0tq/eq3k9qHmFIzqVoKpLmB/
0fSfWAzRt77oBUUpqGppzDWUBgxYDrk9/DmuDGDyFRdA9u5mJCvD9xpcHOdOfiX3
X0IBVFTu82gbRvQDx0nTG9Wk+71H2LXvoU+eTUN0P9tY3lTxEXf4hQ01fzsySUyW
XwTFVhFjmQ3akrgw42UVJQI+SFyRhlXDsOla0yd4usVlxRSZ7z8Dj6agOshIUJ5s
WYDO2iqgf10oI18FozKe3FyEeDiV/R/9VDYs1+ZNw0E/HS/S8yqe9PAs7T9nOCvl
G+KBwTT3hYOMvH1XN6fWAfVx9y/7TNTIdUCYS7unq3mEvxkgzFon8sNF1NMgmqPT
XFtf34o7wA1xXDXsvM/vnpI0rokGxsjKYG9IwJYWp2PmwS7Axj0kpfDQLevyMJdJ
ZaMoMHVruXcN3QI2/MLXSPYiijdgUTvZtCMYgrfcvURkUNk7tr7GAGheTHMG14OG
xEFWHUQzqHrjfAYxvsjQ9gnPIrf3A7VQzs1Y0YP7l95TF0x0DAPkplbCtz+C2ify
pUoCU5DMR+CI6tndpNyznSmr1dJPb4kLZUu6iX2nmnvzfVUp5/3+MFbMSLhhd6e/
2Bt1bfR7Z1c6pPqVa19DQVM2KRfOiUuRIRAjp1l/hbTCoM16u7HqIslJ+g+IUBDR
J36SleXr3Onw08IFTVOI5oqW4xJxROJ3UUNt+IYk7UXUCDpMuxj40uFbnPBuzVyv
tUA3ANXURHLLgDc2n6ci5rj26tCxLc2bM5xyrXnE6Py41Ca/ym08CsUyDR4pXP93
1ciac49zEZxGnula6Ewb1lJE+sRhj7/NFhsNPiIHmxP3KnGXHOq2f0cksNfSaVwz
sW2BtBhkSdolQ+kYOQcic59MVenBS4B73d1OK3isRhqxgAdFA5e/pBUt89pdZWfa
YVsa48sIgRFqnPCHNYyXiJ4QeazJJoxnv5UP4pEk5WjT/xJ75q7Y7QNePPAQIB6b
KYYiceLakQPaF8BfAH4Sha7maHQzA63DbRRSjVyaHMyXLQvsP1DA0GfequarOqN0
hVJ3VBIm3Q1ojP/f5B+v2l9re8B/Fdedm3goaVyaujuuHFi60xyAoFcmVAh4YOZs
EAmQpp2m/Gk4/GbAhxOm8QULMTsPedwQgtajGMU1FxO748gzCCjC42pbVOMhO0ol
jD7mTdbgx3nIkvnBWPXfWNtiHRyM4xHfF+pWtHQaOA9Mg0zpcEgsprBjKMH8Ig+U
KpXV1ZMQo2CosxqNxbm3XT/rf7id83oW1as50NY9PnDpyVifRwp1lW/GGxJzW6BJ
WEWZL3lVZ7yKYRA/8Yje/qI67ARNBCGLGkWaejfaf+sGGDLCOCOJrJLXNZ8+OtAT
sbHJlwRMDyldLNlFtzGFpioPOQs0IHbssogDmLmqfzGe3gT7o0IWdQrsipPOTOcx
lrSY4uU+lRbcXyTnHH7uaCtnKgXDsRtN+1FKyXMood5Hm8j2RFW6677wjP/nw6cs
dhHCw1RX+67+3EfDWps2fTb1+a6xlIWIOOZHdZ+K7VqoAEP9WkpqlpGSp1zEtgA+
4IVc/WDTjFLRPRnixAPINu/+GcRPt2+N4EKxy/HVgRJ1eaqzszkEHg39EldpKIqh
gGdgNmALf5zGjrR+u+VFyvlWV3lqtGv7ZBBjYvAx3tcL6EBW8rSNH3rlCs3sg3pm
lSFUs8A8nXTyz5/TlCJ+deV83FrsNCG3YCZ5yo0dQUVXxy4fqxQ/vDwsT8isr1TU
+RJC2GR/JdyygjzbkgUafW6kKfOlvOZMPdacZth5400X8tcQwn5drEum9hHo3eG7
8TmPSmrUQQEEz82PqlP7nvo+UmLpalxW+C/ZLliTChqRcxkjN6NZ/QXec65MGBDa
QCkUs+E8drCFwOjyZ+aJ/BVGkD3w6s2pHDh8K/ngRVtQcwWe9P514r7LipMJSBnU
k/0n5+fOsQaxeGXP/UsWCWm5tWNMVvXyd3RUq78It95KrOtp4eRpRYyMP9FI21rL
i3QkF9dNzRQnqXUn8fcthcK97Z3JOLRqGo5d/+3ExPHdl0QaiGb+yyGtwEVcERTX
dxBF7R9Rrunu91Pul/SNkVm2Bo9FdTaR4tfNmySZlTCK9+xFE6aIF1wv8Y92LYIs
szFgKJIv6SBCwkfpWMASTZmhC786guJKHX5f9v4XIcUHhkFPLOhcyKvBEUMXESXs
azK/svRvfZJ+N+jmrf1OR9HNOYQ1OOltRGhQ78ZdGllDpp1cn52i6cDM4xF6WPL8
I77Xy4iiIaFPCXk3GgR1LB4TimLmmLM9dsbN+hzkwXnJqCMUGno1EKdJG0rThX1M
rC9vzvwmbHGRphzrEBv2iG65ZwsEEonVLm4XvNHuuwQKJLCExnKHIZHtw3leF6bT
foKCqomEY+2xqQYexVrxnqByqlqZxq1/Fbooh5fPnE+ztAxvjAc/6kQIy1uYYfY2
w1th0a8rU1jqFjrIRzMAfjZSZSzLxzayomurr7ki5ANljh8M7WH1F2tq2WB6IWXw
VrT0RWqj6HKdjW4Mql++98ELu/XSYIVtpj/GLyEcdKqrFmn8Mzc+1RDbvhTvjJUg
1Ob0uRnAd3lyvi/r2ZJie22x0RQ9RxVqVr9Tlf9wW36nc5H52HWeTJmbQMJ7dsn8
iFUti2sY81SI7hlfF85Ml2/03lIyHiIXsj5xUwhamU4V9F2Yd8pkLFiufX+3oY0D
/jnb/3ZUpBuNaiLR6WXQ/GafCFCG3Ue3cXhssFRFmANW/8TGLCol09gfD1afDtcG
8ZVrwfESGxoIcWO4Kmb8cXRqaejo7Q5PkafFtc131AfLpJwuDtT9Lbe4/dAIYAQi
n1vjW1PCLZDpQf9I4bJUle79dW9F2rAAed9SorsaKqdfgP46BxFoiql0Jy8QiUpZ
hDjAeaHMaWbnfXxWXL1gBI53cn5zzDfv7KaA37BPI7fmxj7uEQTk576dt5RsZzd6
+/XcA5QcliFPy3YWk41GcYmJSIzvyaZxAfl4sQHz+HfonrX2+mcl6qqRGBOnXoap
AobU+bWtv5IEfkqdN7gbqBkyisto37X3svlsTNE7uteLbq1RqbMJLK1v0qDSbL9z
40Joj5ixkqzZb7BLyVcFzzRQFGWRje+9r/sv6Lzq54ZzRAHiJfKVMV5g7ZEYZUwE
eUqT2mH9xU4I+YZpRf3npZ2wQZiGrZr/5uTTynTeFuY8/seDrK2af5rW9BB4EQPJ
F1pRqoPEDbEG/+6/k0qbTdagNszrUC0PivDtB8eSImPGONDq3ioY/5npiIBL+yC9
EXXj4b7HX/HoQEhIJWa+nkBDqwaC265XrS/M4bii6NUrypZfMwJyAZYcPKclXtt8
u4txliFKRI08MeEfanQ/xkwEypOTi2xipEGTaby3Akdw+QCCPrfAA8AsJRT2PQnp
RBAaXagJ4RRHldJRmwCX9D+bHK4RAGe5XpYlkq5LGjz1UG+pVhO0zbiuXxwoF8OW
962gNcI6eMqUrmjBWfJbN3GD9zMxLtbysScm5QbRwCEWYTJHqpSF721eJfpLtO7f
xLHedoX5RrJnITn66994vazn6W51x19ElDSxVwi7xBoyy+4xbDfcc9eRdR1lSlpc
lgNn/L94HIbJ5aloVGI8xWbhBhWeG/4ov5jwy09NTogdTBczlhv/U9NeKkY1/D6b
5AAE+E2iVJ56zz1L74sBKnTLblHkwqsvhQ/fnb1HgNgJfZqdQhg9RKBrDcVpW0Rs
eBxpJdFz1LZmClI8YPE6Hlca98Yvfg4xGZdwuuLrEMogwHpBtaOniJ1qjT7x1hbI
cX74GF6V7fYw12SVUaxgdb6VvVJqaVh5xICNhKrrCHPqX1Bi5Rgr/R30OgOxHOWu
NPM67s2EjG1kwQdZ4vVX9L+FREdgTBDnxZhr5ronty/D8L+hfhsEM4dS8WCtmsWk
O7aST+3ts3K7jeA48eQA8meyiT5y81m2IsM0BbpVKigsNK7/v+oRNSmWV4CPh3YL
57U9tOXKc3wiZ/FeXgYby1571d1dWL7Jpf3+HJSeJUb74URq161JWcTY2UOLPpNE
0om6SNHQJMNQn4I31zg2PRNc//kbED1nSzLnXoNE625+plLYGNd2DcO3ED46ZukW
s5I6AqmxupBqo7TsIgpdVPUSHyFqkqpomDWPc0xu2kb10qYmv3WsC6iW99Y45g+i
OaUnxa+k2uk0d5gxmQy5yXXkNoSyJIp0KnI8geL1HmN1ob81ZZlednnCCh5D1pSo
26nlSLQAR/xcQOLYPYPzS6KPIMvg/IZdjyohfZpdH8DjP7BHVh0TjAFdmhIHotiW
cLkdqIYYmt9qfdol2exWm7FT/5ycDIBYde1/iZyomaKVDkwTl27tz/axlNgIW0sC
ACQimvj1s0PTZ0HwAL26doeMZaFp91M89zD0dKylxiStGt+3CE6hB8rPB7LMZTqq
kb8djAewQYxVhsDQArjxqDUi+WUE1OGG5Zp1ythQ67/RBGtwEyuGeXMCcdfIuy7i
bQjLFFi4h4dbcjjEqWxmEnPYbmg+mXokUDAaqEjtnpzH7jV+5QxtWOfROZJ4FsxM
ZdyJm13UnsvOnz9l8ihU+GgLwrB9iREFvtYLHLyF84iOJF6k1X1s3VVgz7HfkQgB
ZZ0kO6Y5O6PVdSMiZQJa9QPxKgbK642BysMIdzOZhFHD2Tav0PpQcCIaX1Q1PoBp
QwUNMe95lZHEWCa0FnuzB5WGuW8TeRkvFrMMFTImQqDR6odGY6/mUvAKuz7eTUl2
sKOSVnwjmgnRu2FsZWVQ6+Zu+4dhTIRRB4355ENGq49DJkf0AjOtiHegzqj4weZk
KZMlWOCxIAaT+N0B+6XY7saFAinaSbYHo3KKedrNW0FE3fnFBbaOBYGpOn4XRgu/
vSVBQTR5NjCdDuW7AE05nBt46Fc8Qi5zHKYtrFnWEMRiLbJ1gSNC12xNAsfK8qCO
y3q/eA9BrB/j/ctTXKd/IYROopq4g8Kk6oYcqvNDzfMBKb20dE/dbvjZlL69nLed
Ot3HS/wy2UOVVy0gQxrWtAsnS1n6G0M53MppFby43awB6o1qLmU/pjRxUU0hP10k
NU04t6XNHPIGCTmeG6h6VMjOqOpDFVwD/Jqd7vzJTm57fW2DhPQXNZupdp7uXg73
N6O5cwW7wdril4tJkDrrzCRWruIHpNIlbUBaA4ikBGFMbI7W2WvKFg8db4gvNzrB
K7LO+7uwnw0QxSoq30oh1+e0ZlxnfPeAdpbpgYWX9iC8pVgLjATATtURHXZghSeJ
REZy/3Nl12fMhnWdQoZU9k5jAxV5qaXDmHn5kCDxoluas+Du3QNXLldjoVJ55Hxr
JCCbB/mUe+GMY0m0ndQCXPXifJM3+M0Z9WjQsRAun9Z3n+Q+zeFwJu1g6ggkC7b+
sOjUqkuAxLoGl4iYb/bO1eL1fp5pCU5qzaOrv6RQc6ur+3Ve9ne28kR3vyf87MRR
MQOxkbCGdffzUy5JVTYOuKFGaJSObX9e5goj4BO7AGWq7dp6i5xV8KeLWf5HFuJi
Uh2QOTvKO0KkYUnf4WaZuyrS2Bp28NKJmRIwQhjGx7hALG86P0ePj9jnv7QzGhWg
Am8nHRLJGcICrFT/BbRji0G+eUEYYPwfHh9tpxubsfhReoO5xKjMslDwZ/6CA+EX
+okADiZR2YBg9kVC1S0iOExluOXNdIyHNOMgCd9JuRsVlg11RNPU+66wtozAt84L
lg1daqSh8GarfFa3bs9+iK4Fngt7ToFDfloKCw7oe1UgtLbzpo8uKCW6ZgTEY5Ar
jVK6d81Ko76V3tYGx2iyTZ56esCKJAl8lDe5ydzjcHXTeZgXlqBSgQ5/0ErOy32H
aUdv0r6sQvO1t2edm0WzpJFPY4pYlSYLsZ9bTKQMt9z5rRj87k6RMNeDixJ/zaED
nZc481odbnF6dVQjHTvM+2DkIy/T4SyCjCuyFWiBR5FYpYI0sZg/qdsqpaWJRyT0
mSTWwtT/rfboMUDtu6UFnODefeSRooVtXMZUXRiHPOPT+3TCSfE+yjxq3cuZjEuT
hidCMnKo8oFskHvo++R8SuzoC44j+R6IXSP6v5KUUXVoBuhGoxaaFYe2NDMUvIy0
cjvitPngZ5zpwyA0oCL0X6J5ki2J6QRp0Ca/5IWHeSHxDeL8M6Pyv38r2ZoOlyij
UvZAM+hOxqhW2fmh1yygXeuDnJ4VyjHZ2OxN9ZJtTB7lOJ4/kJ+jpbdL9kLFpe3w
Cd0UgzXSU7SlUkYiAPweax5Y1KQrD53//A35X8EQyjpxr5rWBfZgUI8riuNLR9KW
l17j4SKg/Q3XJbNhLwzgD+0I/A4I+MdFXMdKkxOrIRaj8lpjWSpGsjW01CFYPrYa
GVBBGdtmdRCZVYu4ITl0YHgXzM3apwHXXm8gy+XjUxIRImBbkZ75fs7AIsiF5bjJ
ynW6n73rH8d7uhZAQ52/cKorF7VYyu8rRc/scG/hsIabsL1BSqgh44wMmiPk99nU
U4i3Lx2B+dOUkYvEmt2iZQjzZgkHQfV8Hxh9zTU6WxBdTspgMsPBgUaUgA0VYEWh
Z2ijk552pzI1ZtpLtbVRxv2d2XtSfHXqEGj9sSWGSxZqZJdejSBwklJZj1uCWNPx
78M/57GGqJHebs2sy2TVU5IhswehQPS3kjZLkvN6wtJRHvJ3po3uUY2pqV/QR5VA
q7aF8Mfx7ZmM4vH+nSnvM/aKG6gjyI+3EhMmJu0Ja6QE06dutxEE////NQkX0Njx
JFaT2XqKzu1Oxr8fJStbE2I/dXHxzTudnvAGSe7TYmruLeGLt5KwC9Oc13K3a5yy
+im01dAx6/wtrZHw910MU3PVnLJw8kWy3X9FrTflPTf/6/4GWVuxgatk7TlUtJDz
2Ii7PnaHjvFiNfPa951R9dXwbw7eBLksucfBa+S/kEw04PmGlSC4zdc2go6nuCn6
+uwo6hwkvToop2NkA05mXyr3x6Ytjg9GkYUOsGlvFubcvY8grt4qeN56ApdaeojQ
PIIeChLDfNsLyADkj0mr5dO3/8R0W59G9IFDK2oMaNR5pZuXBLeJES4rOxXvHqj3
gc9JUf5q/c3+AJMvRZKCk90zzF9ppqEbaxc6IFVMjKmdLH7J6lVx/POCNIoRxgaU
nr1DejE7Qy9p3LIesnK1u672elHAv4eJoKA/nrG74FYAtus5oGpZBEI3J06HqqUQ
Qesir5vafuejjEZwA/frXhbM7qvVLnsJ6BvKE5JA15oxgl5AsPoMU4+r9otyL0Kb
BCjcm5bEbMedbKDNBKHvW5BdIDovr4DZDcGht5aMFmeBxkAyo5yVHDunnW7EcY1G
HBb3tIwKDhLxiTAe7kT83ArnosOtCuPBatz3KXzBIWagnjTJCY0UUfEABNJ650D7
wVL41kl3hw/V7Fd4mbB6SpdfnCQpTUpC1Osn8xkRtpVdRT2j6cUwMQnFWhXYdWJ7
+8lRPPnRGKldS5ZBLHxwnGVtaTiHMQO/CTViY2VFA/7+RtY1z4z+v65IAFaZHTzN
HHIGTZOeODTu3dmss4MVE3a3aKCCxdg1iQQ5wBu3WvnJKKiJ2t8YcKBb+Y6o0a8A
xU0s0s9UsmWTofPD7fegeqdhT6YTRp62B25nUaOYVHifIUo5/Qa8GPECoYwUzXgN
vKcA3/T9aKWxbnSrX7fPKj1ru+krjSLBQZtfaExt/iVgsewEglVPRXrCkkL0X5i6
+DJAzaq75LRl2yOi3KnQ0uYSWwKkDU2qtwkymmmF79OumXzNIe92tnIsm1TjKPr/
qH5yd/YRw5B7L47YKLLhTLK5uIckdyjD6VZpmuOy5e2FOD+3vt4+WCxSyGROOpJc
nKmv38qEnwX17KaEGrCDl4Hban940jI7a9skSQB3Wy2nxTuJeVrgB4/Y0L/AqQ/u
CBFzmASpdk8Cga0reJjJemgjIAWPNjffVWTYNc1S0m73HinsJVDKRawj25us0t3K
vWVDyG/gJuxDALx9ljmgTmE1/MO/t67xgsCDqja6Ru8k2/MHiobuR4zFX7arLPJ1
/LsZ0EBiGW0VSPkP/gtr/Lv+vDkX6o3zW3cru679jHaXJAh6eSV8bR8gEpotLmsh
5Jbpq3+CHP2hxNUzpqIAtxoq4sFBiv/AXQBN2zSEvtcpyNzsQH4r6t9cDuAOOhs8
ij7If82WgtoGrJTXZbCEbX8qRxABxMQYskjSX/1JzwSg99tdY5DFqZ7WPLfXkWra
hE2NOUthPy4fO9ztEjS8s6Xxto71t9F3rs5Vv5Bh9Wo+uShOYN5VskkIVUBq3HYt
UcPHeoOwT0RQCUw2iDQ1flFsKDuF5vJp53uVFK3ucpPu6nmnJdjKw0Nro2Z6TEne
BzxH+2MTjvff5Gho6WULY+8bNAuQmpaWo2sPRWqQuvfbrFWb4Gd/Wl0+pKDdp3IE
qLQL4q6ku42hEJVLKjJabm/3r3SDq199XzvtE+prYa8xU8tiRfwu5JZXKh1gauRv
ci+JF93MctTjuYnANDN7fdVMBBtC+cSxfrZn9wHzhluaIzu0slpTKOF27JnSdsa7
og6EsO4bpkGzajb5883gPIc+4MoZ8tTV2GgBcQTVJPU2X95CG9mxnvC1p+8PC+bA
MYnqgpYex39gghtVwhd1TtBeRt5k9oS2ogPxgIAUfO7ekXoEgNb15Ht5wcjQVm7J
fAlkfcVqoW6bUnO9nci2B/ASxgrHh8mly+ASOZLBj/owUZHomLxQz2fytyYt+3Fs
CUkRMXECwv/ybK2cEpaxLcN2pNpP1tpjhI0hPHonpmA6Z6WXpU8OT6ehPnshCV0g
qxGFVIOaWM3qYl7UF6voNw/nWvc9Gzc85vlBHWbbMQd5/DCg11ynvCDOmzIbgQT1
xxxCRjsRZsq/CE/xeLR64y+SyieObG+cAsRHN9a70zJeouzm+qhQ/PGTdKAqVrGy
4gg+++4vVKpKdoQacz21zWS8fk+v2lRZkjG9D0yFwQWmhDuh4QhiLoyKTsXHijFX
G/DxnyHjrLZqbOLZMlmxN6WbCnnBUvcg/UyCBDdVO+A4GMo9WFlnrFZK5jrdfVDS
d1BJl7PdEGbF35M/qDXP0jR86ciic6Ts4S3BBCIEuqQ85g+6AkBn3eCrAmrO01qY
dyzx81aW/2rp+hty8/KEXlxQtq60XOHhTxu/b9vsiDOjBCjB55f22QwNTbNt8cWU
q4dUq4c9xZGt/U1ownpzleRyh2+NIMQ9oPRsCMw9ACWZFA4Y5oOQ/Xv71CYO0bGF
+hEvP4VtzgMdeb5HJP8APRXwo4k3rnZxnvs7Y8rZBIO8mkBLqk90BOzOn/b5iy2r
wCAU6UuPl3I6P9eWQ5K/I8XnhXaXqqXBXvXG5MRx5mv7XqS6CUaG4zL+m/q1Z26R
tjdjq3Bku+DmZYOHrAGD51qPuPbrzZcaHtiBY/vRU5FIa85rNjFAjJRgEECAK5rA
ZiogTjQ/QSgF8+4f40S5iaYXpvLfLw1rg92WGv8PMaLnPFan/USkMk1kmdQZ+LW0
3mKp0o33g7Vjhcg/JFUxVdh9/uDGCF2e071oEkEEsgeM1XG6x/4JGOnLQePFyhhk
c0eE+Hukox3+UVFD+oRJkASKqpWETQa57IkgWbme0eEXPAoLWKiUEXFGcscMwlf7
z1ElirWc6m/i4OpXsOYr93POedM21RiLWvTbFQUHm2F/uv1tSz7BQleCQzYM2WXq
KXs6rKh9hbRMMG0WnqPeDTNZLZODn0WZ16XKxWL0HqE4LFd+ziriYtfemLDadvBK
MzdfPKB6QQKAGP9HZxGjDxwdDAlCFmadnEs2b/Fyv3c0kaghVGquzT+lDdwLIDs/
hM4IyDI+400JzSx6euWVE6l0SZMI9Li2QmjUPAJgV5e8LYMmVpCkN9DB/XfORb1f
DOIzqvGh/fSdqx4lp4Je59DdCHJKqOa4ROrb9EgYD5mGjmagI544PuGwJvfD6tnA
RTMsqjnM537nPQOLZCujm9sX8f9mcpEPmza8Dt73BSnyBxz2kYOmre0beVQxcHhC
r4JBm3av17HFtBxN72T3KRKEYf5jvv/kCpUO0lCkV6jLeX2VCDOCz/hjI0R6jWWD
yX5Pa9nCFDouqe7/kY5TfNrpFapoqUK8nXNvTkHHVQaFU6Evo2eqBkgGvGNWrIB2
244z3E6TLZXawY2duZpgPqZVcsyKJLBqvFI9Dgkuu373MhVJVpODqBrG2M5899lv
jCi1pw5vBm/dEULaCtKxYmXo2dCbwe/6+dfLOExosHnqVvKuLc31s0ucSC/Tt8ZP
QKOwhTNqxgD1veZ52gEGiCoD4lzckShOBc3bHIbwcS3fjplZ64hN0p+06iC8mMl8
DeWCpkirmx2f+WYSEF/wej2JuQ7bCJWPuZbEJlMmnrzsZ+JVRXlY3Ul/9lLuBFM+
RCoGuKRfxsR+mBQ+JY6BljzwRhzt0dLMnupZi24zFHz2kjZnZwEn0c5tl5tz+fFV
tKDBKvjyOvkMWScHe00+m/UL0LU+Mw3rgAo9IYy5lB4JgS/MUmZ5fG0gCWyL9RPj
QR30vSuKXd0/2o5tYjKR+rYQK2z7LsS4FWIC8q+/K3gsyGPimwVs6DLWkm02Ywq1
jMJLjJGXjo5s1CshjVmgOuz4s+BWTtZeHlweH+evlW2j5JfEY9t7lWPzQKuF9sPs
BOLPAv+2zH4LhLpJC45GW0b/2QILeGjYb23AoZZjT6jYwa69T9y3tnR94F5ElAKU
t0h2OCEO6y43Tf/KNDGyEn5Hiz7yf5Jr+Av1CUSUb/zGONVQQZzPwCmnmTo8myQH
BqA8VTqqbP8SXrx8uQavZPMz6dWEFcSvYAd3Xk+D1mOFkYonUiePTe9wKSxeIfXS
LLzyJ7cBqQMyFw4plEXz4XzgWX4oIJg3l07RDGGRkyXqxJUhD/WW/38Kdn5/P5cJ
yjrMWp7WP79rrGY0eEoTJkY5mcXLINI/mVQ/KGGdpgpxX96qMVdVouE8gX+bFYFt
T26FEi+yC9wUkP+bOsihYSRPzIUSN82FwckY2KEyY4B15nbolfUN8mJN5hGmSZZ+
a/ClVXVUbtc/3TgXy4uxmooHSKt2YrUiyw/pbtVDm1r9lK4TXE7se9dW0zrmLoWh
7C9y/5Y2VGVkHRhAh88exlgYdZBttkkEpDA5NRBDwGEo2Xy6WK+rXfgd/VzoZpiM
GjAyt6ast95HKPSzVaXb2XKbAhzjTnhYW1JwuDGPHOvamC8eiM377aJ+COxe1LIM
BA+OVIjTuUS/XYPTmOqR8m0gMs2+0s/TI1C7M2oPdrFqipI9pEDF89nCpQT2XgMW
NlCrLtLZvj8fpMuv4UKXYofyQLO6fTPUJJmb89MhTRtAAGDFY6Yavxzdc64LFQ5d
+dd6wqf1Xw16eFfmCwzp5FV5eoZBFFPaoJvRStgYS6IoZDJPHBJBYb39+zcLg6mI
wcVOlmRrA7O0KbUiOSSGPO5SLJ9wyJM9+pHln1XqUSQwIJ8uHydvkZLKb+Wzj8HI
gueFtkCjrvFFLb3AFJ92wjfJ9EktdRKME0i11kSV3y8zBJ+0pyvVWYcz03zTRg0y
mQFqvM8TvjSUH8qg6PCDnzYzffmYRF9JOD8Ech5JptzlXeow1NFiXLz1bLMZNONu
UEvO8u33FBJiwhfYeCCOy55boS5PSn2y4dab4KVyp2mvYt/NeNVbakwD5gOB7AEf
Yn6K6b7nxDQ21JHW+ByXYvmjkqnWf8J56T7NwCmGiooYNYzjLcZBuY0U8usEhMyC
08kQIsDsidIlPf0BLRuluefJYL2TQVAyE07InYNh/o06eXAlVeLshc2Lsoa+Bjcz
Xe6sJuFZn/IqCilCGKmzJK0J7P+++zODJClLkP+ZbK64Ude8uPeSCHsDWY+ehib1
ghYPPXTQ2YqH+wWank8Loos2+D5vMNwrjpDeLLI5+O+Kp4K21VBU3zEwErzRVGCH
U/l+K6moDH6GR2dmrkoo4tEFZg99rzgkmzPqeoigOjLh4W4JDQS7jfkV+lC1KdvM
LYRx0wZmwGMrQ2+GquV2VQZ38nAskx/pJZNrjhmrNfPLDaHNvKflXfsY8//36oDn
vV73pFJ3eBb54+dGyFJO51+0VIaz9zA17b/gwOBLZFNSOnPInxlskJUOEon+iDmH
NQc0mC7KtyiAV/6AmLwf6bBnVDL987RgXFPyETicFurpxDOh/bBlCOEU9K3efQhI
RmxM33NRpBDfBPD/KRu6Rf2AJw8e6jrSeYvgXdE8Ne2jgMIk38v4M0O3OEwoYXty
FKpLOlF/KgpdhSWH+kP0+HbNGyH0ZAkFFZEtjpgGsydKe2Uau7FcmWDIFLWvyxnW
JqexLRFwEsj4uXA+1TPM+5MnH8oyxd1S28Qsd3mddoEhyjL3Oe7fpHkprawZC4fd
nqhdBOrtK8Ybw2rN0laTwlO136pZbUZf/dkeBOxE/AdZ1TLRkrly54vFXNWY538m
LDarrZxE69VvGs4heSSaFO5mAbDilBuTLEL6WOVj54Yn9ajZUF1dkq8vos2ReePq
B0eUoxmbQF9weobD3kAwfys5bphJPa4Iti3g2YrXA7gQc/L4WBM+eDUGmp0sS/Kj
++5CWUVAkoa4YqbcvnKkyD29QiAISzfegis9vdMgdU8LZGrusYvAOSgd09x0vbvo
YPuggXM+i32HM7g6kyEr6c24TOi5ij9y205/TkL9gCALey6VopOzoj02rnOJp9pB
6zyI22o0D1rm3LUiQ8fU2zrTn8oish0KtoQ0I6BvI5/yJdWCd2K0COobRWAmOwv3
x9Y2FNy62X5sOfcmmlWCU3jvZQn6D2P2pnkmyMJLI55zTM4Lea8xzzM5PCoPCi8D
YsHzdjT/yIIHzeExKc34cQtHMsPVR1xGO60n+/syjDBneiRprYJxyUGeCmtYYxzu
q0TIIXf2BmQPeOYiCzuBAT3TTfBeU6fn68nCFQlQK6wrp+eQwlntmJZgWzFuS746
fzXMaTf/+LXVHe2ISH1WdCTkFhuWuxKnKcKUqmCKeJN5gz6cB1CSmyo9Y3P/s/3u
ANItvfiPd76hrajchWczBPNilrK5xGKVp8zXEPf8I+itiz12GLDLcW3a6i1UUtxj
6EXCkXxKoScjlSIlgVzip9H8hGejHW/kzlsJ6LYB63GWfr7jGvB3ZEQMxd9MgRSP
wd1F2AhmUpZUUNuVh5LKfmBMsk6Xw+u145m7b3hpFK4LwSsvrIwZuysnY/mCIY/z
24dcgI+BRAPRx2Vp0ywvldkCr4pvdJm9lGiSYid1aLy9Y2Vd8dpaSt3jVkyBeqwh
hO6ZWQZwceJNJ3JMEgMigYoPdZBea2/3P1d/4ejHLITrTT/r/Lqiios61BKtOExN
chzzrbBpCq5NjovLLylA53TPCK9D8NM/NcmhQri74Lqg/I+dqaR/4xf606PpXjKJ
WS7NErCotNFBC4LPEIpweCIPH/d8NX5ql3HZD+a/MUSni0vw40Xo1rQATCrujko+
xT2ovJbQnb8BRqBv0R+Woujh+nfnJ/gryy/NZB/O7cHeRhdO5lcX0UlA9lZ9tXUv
P9Dnv3dnR+nsnfAUKK8f8PTNeIezn9yTVaryMNAQ76OpEarDFlaw3N3bA+Q6mOkr
9h22x0rJRRWs4aWM5krGcZYPNyeCX/RNnWElZ8N3Yf/Y1G0KAYqrakHNABVo+2mD
RQE5KdoniWBzfGntzRdWJtKsiUdJQCC3Mj5dpdE6KcWBOjz5/rEhSw/ouTq8VO8M
uGlprPGD4vOh0zsEPHEPE9VzwAJY+7RF3oSMKM9DqNBtIW4bQ3Bnqai/LGiDENG8
TueGd6a3JevEVmQCj52n0MHWrOMWpcOVB8wm2xMu59+tkMajo5OD1eEvItyjPWtV
tJq1nMRUxHKYfgwCIaVJjtC2VQYzWorn3lbh2hpz6Amu/uZp0j7W6Si32nIjl1NG
um+5eEqQBnyIoJXuOHHOS8Lzza+tmqj6r8hyKE21LcoWk5LktaNEUTpxYOQEBP45
a7qujPYTJKQASMCAm5/cLxZvVq47iw6H775tLVlyUwGVKbO5P+lQozeiz+76idcP
XAFs/aVndLOlDpt/CANJxIiLvQMnZhes6/yh/rQtzCjb+ze7qGSXw5AOxTreeyde
xiLQdR//B+BES0MyQ9Mi79GBf0G4inEY+9VxE3Wc/VhFDAdoVnRj5PBppYIItQjU
bfGc7EJ9vAwkDkoj+nG3wjBXFqZFP+UXPb7gz9emE7vT7vHHd+hIvLYxSKUlWmag
Tg+oUMTgMN/4IIAvvtATkKyVrgN8l5lIRMLhMh75tQp/eYDvAwIqLEl3jgvV1BXR
jOnDQWTSUGPCCu9nnE4T9WE2i7S+3LGWy3M8qqwzxVMvuNahlmDknEc6K5uI5TQa
/Gd41wZGkqdQnro9tfQw7aHSgjzhUAlbULngwVutG98zMXo2ZaPW1QibjUN0EJ+F
H+8rdsuzBKjUAM3XIxdFPL+lD1WfkyNgHMtwZPnRCUJ/PLH6LkSv1a5YCG5b6Vem
rqUAs6smI5Nb70GH+Zi7rzmZADt7Y9ODcvkB9Fhjwcdpu7aPau8fXKrVWa+PejH/
ySZg3Ew9mdBQISFAmHIXeKklry9yOsKO+y9b+4dEAT/d6f9OLb1JzV1uhmk3w1dS
7BeuqMgqaoY3RnTF5KXq6bWubBKaPewtio131BMfDDZvv5vOhZIosbU+jiGrYClo
F1sLIVTbyqgkp10wNMNwqHbrAg78kKXVq/TD9N/Of08NxTMHcIj9HHiRhldc2ZrS
ipDgqmuFndvt6M6aRsSAbLrp0m7poRuOo/ysZ2wDOuKrwKyQWhnCf1Fhqa8rBJj2
yvNYG+SrxX7cLgARkalML85WW+MEdcAb0krsiySy2h4whIWUeJ5cyPs1jMV7g3e6
z+YFAsQHAv5eYFBmAXdGjS/AJVOl8j1Xh/1raFNyNfhlSYHL/t8m1OC7stZOyqg8
DbP9L6zl/KxPPQ9WlpttuFr93PY/c96ZrHaWRawENgQ69u6IJ6sHVh/laYa5ao65
Oy0dB5Si8G3r9p2zQ3UxCXoF0tKfGPVQs9LjZwWHW4rebmW3AWGfFFMJD+HEJsaQ
kBGJwLsatVWeQMiud4e7TZS0Urg5nxSfi9JXNyUb/1VfDVbf0wuWMY5jQZWkK8SW
iMYQ+MK4WNA7B1T8JDad7i/ILJC+XzOj6DYs/IFkxPbvfe9NX4cVYUyeMAitylr8
mCAUpiKcUrgHXjnHX54N9OA8EwE0HjjJyQ13KGazy5PrXkKxn1gJyMldcz1tc39r
9/ioEeJA7lII0KEu55q75C+KxKxpfYNOpgvTaPbKMR8vMD5IiygWawHJzp5pHlBt
Bk9PVM32Qe8CNDl4zK52rMJwBReflXcC+CgYXcT5sb3lhKA7/ckeu0wQtlC3iQzJ
1MnoeHKkdLJHKK/SOVX6Idj2QSqboq1mIYjTMqDQapbXxrlZdA9TGmillHKB//H2
ytr1CAq8LWcRenk/OltM2pbX/aMMYBdD1ouvz96pqPpaLfmcwmGXt0XExcsVgKDi
uPEWZVbtxe+jUtuO/87bTyfaedKxQOYVuNhqGK7Qo2fMtU2N/IvgNyFb1w/ysaj7
9cbH1TiM1IUFZfqL9IxjpxMIXx+zLukvUdDummhGVuHOwiLoc6eGI75YM0f8RYOW
7lssMt5K63B4b260tHktRjYfndDA1zFncs7iKAgxxK3XiIxVM6OT1n5g/gK6yb+b
ooXcRVTm+ASdtYR+wmZBfv6Y/XrnJfAHga5+uKXdPU/LtRQu0KNVPbdsCqmbFapI
grhWdBxp7fZliZS5OiXz+dz/Suxy3dgvr/aR7PzttIsh8pR3h1T5QaCgNJRoxaQt
992vBPFW5tp5SpfFYY4DL5mOu/fGGki5kTOeSd+sRgeXYj7pXlk0+iAjkNejBRS2
jsD4MhTGSq22tKixaKSvAsdlv7XScn+BsUUfguuO040DGLJuEPOwpCRbShN3WZkY
Is82uy9VwWA5a9MSFJkTLLFrw+pDdeICfqOjLQNn9RUk/skqFJByiEKStyOVo2Pc
rznBtTLhpooetyUHezBQ3KPij5jXoRp8hA0pJjTJfSdQ53wI6v8U7YDeLgDUgBEA
fPhAa8YpQEFaW2lcu/Wg9PwAClyNoASepu3m+6JkiR5EwU7J0sqMMRU/LpsxmudK
eJTlJqHb/0iNmmvI52RrZA4C17KoB8YiG7ndadtdQstjYqjIEM+RyBA8u0F04zFe
cO5FYCoO7dMUf7z2dCof4QulKeA1Ursfh2WgmBu8AP617rfgFzVJ2Wz9epOs1Bma
x1SkCod8osvOyIxu3ymjh1Om6Dh971OT6pCZMTYs84hUc4YkXtWFpa0798nBXD6x
gzCr2Xe5MJunz126O4+oMRSrjqNFE2/CH+Inxw2zPOwJ3DhEM741+X/2lUBddzMN
BHQluZUw5DINtN2MdVYcXfE7tWj9eS+aHpeyTXRfMV8kIolCuqysJM5gd2TO2VS2
ge5paMqTzU5iOP6s/C7r2uC+q67aOLJwn0A82HJ8jHDCkMUOIs1ccmcvOCg3iBk6
xX2GoPvC54GHq0jACa6t/oXAdNnumBjMLN2gwT95yAVig4uu6+bSLgPfPxtH4LK+
gkWEBaNbtlU8htixzxiz6TLo6k8T/eBHMnK4dT2ga31bmGA9a5krPkvazChpSiDA
tAY+0LOlMozloKRFTMVCDi6lAIWBRaQ8Z+rkuGTp2igog2m4qGJyJ1Js68mAP8GY
kn7rZIpGn0MFg1+oVXGCG7gPOAkLv1Ydzx8HiMfZrUZRvTpVItTOcwwiXIjMuDFl
snDnRFkwrm5OETwRv35JAgK0MlZzcA1GbiJAfNu39x+NAIzZWl49k7eztSSOGhgV
0KOIMokjTnEAbab6IAP6awx0VjPDBAjL/odnN09E3B7kv9CyeMx3dwZVqaSbKYYv
LgstRd+fHf2MR90l4+qn0eLQoyRQ5PYvKKMKA6YqGAPYSgujA7g8YZj/tMrXJZy7
yb0U5xmgJ7TUqTcpDnvFMeVBeOvBf+EuXBgjkk4a9ZDZq13W2t9AGOHZGhEYYpd/
3HAymAsh1GZ1dXaBW/5s9baKZt1JYwdANmp6YQv3QHHGu1xpys9cW6vB1Satd6sf
tfg1fSzHbhgK1WLjLxR1LLjuwRTY1rEPF2GDtN/F/YdWTgtodCXhGZBmb7f2fohH
pEGNUUexxQl1/cNYSMtss5nKyKAb7BkCSlZVL2QOz4eQ1RmYbueSNNS1ib/U7Xxe
/Zexh+jn3LfXiqsUV8iXGJrIAIyVSYNN4EFwZaguLNi3MELa0poVfPNsIgeb+L2j
uWADxMqSv6OO75HsHjlYfsIOhunxk+ovLOmPTOXNv9zSWnp5Mg1D6yyUPBsZ02t7
/JhHuvde++Bju12nx9ES8mzhub2scY+51dUS1Cwa/TRaKwbsr1GNIqXq3zr0dEXA
OKZ+6w8fftb4JWPTLepjBpd41DpRE4s0O0TL8+/4JZkv6ENgNIIEEZkJ4YANEjeh
ZPvP6O/ynviPTQYa4B4G8eZPxxb0Nw454FjY5yyc4rNjWFItHib05q9m9eS7JpPS
kmXqYTiruCK4NlPaA+orfZ2LgssbryKYjiIsooQl9kOXu3+csaTsf5x5k0J8VO98
Lumy9lUGuxdrkrjaaazhNs3bbNYcDs7KbFCDKHS6I4UB4L5h8ewYv/L77LQLEy2c
/GSkVolSLSOet0zqRkhr9e8A/W/kQc/bAgUyh0G7ChLtZcShudbMEF17sV0tKInB
dOjDwguBx9B6UnTcqZyPQcYgFK5cUUQjPOXJyI4VQvYOlhgq7LjQB72OGJ1ThJZx
csfMv7wFN/3c2f7qUMg+scXhnbzgTJ2p/xBzuAZ9xYTqKE0oE5vuC/1v3qDAwE4n
au0ahz2HHInnCwf0drhoI04TsTHOpu5a8cVa9UCbhUo5GbKdAuXAsUFMhWc8sdv2
23OdbU7Bq0yPUu2TFgz5/amyJ6CgrpXA8WP+gMJtMwxNhJJPsAcckWT0+zvisGFJ
LU5o0SS2QUV3SbHzxiaCyhRinO3ss85wnqk7G9sG55mhZJ13ZzEvnKHCG1RIWXxi
mE8HSPX3k1XwU1Rb8CVbK191ISzmYdd9CZ2YPmV/YQfNZjYaJlumXHeZ8nHpCtX1
JW90TZuS08waB6aut29RE0fW5F3kHYax1RDIBr3mRIEFkHdPB6655jz6Md0ANW6k
8Lpxd1tAZTyLX8LR7gwWvXxBLzqwQm7jbkA7j/okW80aBUEIMnznIRyrytvn5s9+
jR5MAorKafFPXEzaNY1/zZNmq4/dSgZokBLyDCmuqw7TDbyiEfogwSWNrlzmjShz
BNSTsuzKwSPvHihzun8UPhMXPfWRrQPGzWiFDMCHfECzUWLOU/0ML+a/26nbVHQ7
tkTRoLQba0UwIz1jBPZ4EILBgjBqol6WrdcLEQE459IpUXVQICwFDI2s4IoqbIOk
IGyIX++4DwqpNTpldvQM9o26uLjUqRnkZTp6TomleTCKL2tET/ITjc6x/oPBp7HE
9VoNNnl3RFkGtlvX5/J5N7UNqDCFEogST3QoQv5PPrtZb9+11eERDrHSKRWFuQhT
J9S+h1nvUJ1e1QIdLuyqsg+VzOIngOafau1mH8rWypzYEHULPepzfJ+FzHBpz2nV
p2CkKRHDqMQ4rsm9AqDvFhQPBP+jcR8PNQ8znkwhq5VKXxi7WlhLhuRLJfZ8z4v0
sQtQcPD86UCdqaj5DjRzdIQlFBv94w7tzqAzY+NyBj2AHoQfdUPzaXKp/b7/cf/l
A/A9zwDf/wAfAJWu8hGpK5uY2YW20J2JN+2knoKSwsfPI1SfzEW7CwWzlv/6JaGk
cShNmy+oFyf01wb+ksJZh8b7BRP8sj7ajo2sSMFCaIk1K0wbQA0HteVc4aVUSfhC
lLLO2QKYdNfbecn7cOUTQOWKlNOTloDvh2bUZiItSHYMUPYF8FK00Djwha9n833q
+emw0tODGx6k5HfPqZnHD+AEAKvO57/2vkOZBkPU8/WkJSlPWFzCysOm/D+JyKop
DDiEos4MoAI9CwY3Oypwb81rbtFCBadLYC3VTXfx5tfATiT7nmTB14raT/E6oz3A
8X3LKjOSmoczaUQ6gBrlRGO/hxwdot4KjRILT6pAkoHAoAKFIwUyQ+L8W2BlCN8p
PEK16WtbZ0ZQE5+7PG71Lkx4a1k1+hXy43C7WrA/g4yjL+I/X6H2fOArXHDWiOs1
L7Loo5oIn+PEvDQr0ybnAD8ffbfBbtqvxB+vCzr26LuA9g6DwLb19EHRFxHV8nfh
oBHkYwLJEd4qCeeypmB94LtCThZNcQ7FdW5zYEpC8Hzv+8b/EJCv6jyzQcPwF2IL
rSed4WB7Mk7g2HCfKAlBEpL6ILR5zID7s6oWENqLBaQQQQOsC7hlIb504c91G5yC
R5g3XfLRtlQn5joUrtU4kXQBViNqg4yd9e33LVpUAww4JLTtlXfszks2+A7CXOOj
1ESFHGoyhboOuwLuNmdw56Gg2gv90bwyl6WfyGNqwDFgCg998QV9qkHH722lxC5X
iJibNPU62Aldnf/kDshrQpOr24/kniG2X1rRfcW3w3RQY3GslVJKnFOYaMCdbRQC
n7Nu3RkAQ67JWMlO5zSCatPoyaxrpT+C9gW+6gjYQ07vup7k2nGm29smD4xoH2EG
0fbO9m86amkQZOrLGOR0A0zFwxPFZqewIorUxS+BrGIkxtlE3yaf8RbOoAElbY3P
sLrSAXd6+9ABClftl4WeOMNUT/Jbh3nEi0iYL8cnecuUYhEKX8svrT52Dt3XTGxs
D+KdZ3SSYHc3MCbg7wa4EKiWKMXOb/EF3DW6PWZ3qQUqeCXe90ROOmOHPqZKS6UP
OBYTcXT4LRaJzzH2JzUMz8m6UkDyUjATiDOXbMSZtW0ET6g4961wCvWxeAQH3jZo
cTyEk9wVQC6WDFM0bh5LD8dzAxBKwUd6SIaFImYhfHx27uioWDcN7CLbItahPXr0
fQT9C8RB/gflUyhMS4pGyQCfMePhiODix7+mYywK3VaG5YSgpJJz09xlq/E2/2Pm
esqt+RE//wicut584Y7U9jm5ih+5EXKd0h2w+O+fa6MOjaLDkmM5riU6IPjvPeiT
xZPHsBNo8TSWbjpXlgGMQLg1yS0yN20A3iBBhJrxS0TZg3h1IFdGIGujN8FjdUE7
4TUDKrKcpG4gkooEMbQk5u1GKrY7vrVyXV3pB0CTUPlfgUjoyIPMy3mB6wCO/UzX
uLR31YXdCLVhvAoX2ScX5yRkhdPPTTSVBmZpWMjY7mCUDjD9H2fFSpvEiMTuH7yv
03jcDMqCuaGJ4Tx8Ig3BfGy2jhXliBHml9zbiPuBs2cIUF+QfQghQ4L8OnakpBch
L7G2sADyKVNgDh0omrWXholBHw0Gx0lphWukTlpDEl7BLai6Xkh7523Cr8ENBZKI
BeAkH4ab9LMWAcnjuw38w+m2V7hVO/ugjcf9nKxgULLHsgsjJbXDjGsrykfHlxik
i9uYJe0TdWBxAKzgsAthf1RV7/hT1wnUU8bIWXVZQDdE1+HpuXlkyM1HstaxYchr
erGsoX0wuM1APdReZHhUNzaQdoaYwiGnv0INwax7recVWGdJG9q25I+/FoOtGlBf
mlymP0QPSVEI+d4BA1xyW/tvSLPunA7z1SPvd1xExTdeURGZgcHy/EZQlo++o140
TVyQXqod4WMp+EjCaFyYsO2uA4ux7u9LDS/sx1b2GlJR1uDQKCSq0Pr3h2Jt+ju2
f2jjXTqEYwTkDOPrT6PbPfGDDwCQPml+pGV31PP1avhttXK6pP6zkgF3iomoUz6x
1CtVH3sV94kWdRFgvloS0DWGyj4bVx727qwDKGRwNiO3ULuxsmZ8rbyaGmdasvSo
kZ9snyAE0sGZs5DXzYOZOV3BLjUeTYdUsPwYz8e1mcCFBC/gyvt1ss4J0bQdu05f
6h0kPUWwkJZjSyqwBX5XrAVBwZQKSkXYTIRt/oKBkVwzkNJUhIC75qD8JtopEoW+
kecU1H4ln+Us4LXhD1lWZWQ6koaUycFtHhwdwPzDg63R8qfrJS9e0E7OH3qdokDE
wmifKli1kw6bAFtfmSjmLVsXnIE1/kq2cHpILddjb992XZ3YL3eoJS0jai7vKwID
yD8N9Y7dUqhBCju4b/+DFbCiuB40y70+cx3iBN+lPBaqVVAVFB9aU7zh3orVrbwy
iQy+xpYoM9iljK5JnwRUz0AAcXT3zaZwS09lhXOC0V/+OYBv7fHgran5Z+SmhR8J
rCV/t4Lmd4ihqRcVLb+RomIOd6zqChEF4DGtkU5TSqK79EwqKjPecxE3ae4h1496
yWghHzZQ2NIgZf3SEvIbh/81STHyZmmSprFI1REqRvtETnLon3Vkw/8/C+y5P4aX
qTZVaJvUXrEwR94kR/dDPLkOO6WufHPGsj+rVdgtmFFM1J2ags/nrflcJW8fPHuO
/Sw6VuO+AgYXEQPGJO6CBQD55rLTF34haeGU/9R+9vMFeS6KkII9tsNmlYOSwPbf
yCMakV7WVihmu9AZPK/0upv39WSoSx6M7eQaXZhJNUzEb4C70RsuJPZbKRBBtUU6
dBVlmA/TLSOR/YjxU3gAn2H89hfrqbNpz5RU26XrqisWomLHQ0f8C0mEAY8V/okw
sldjnHalnF+hxMQ6egduHjjtGT9exDX51c1fm76leL0iiunxknpV8MMjQUDzPIMv
QxQq74zOasJEoxeE5UVxQbvIwajUWxb0VRoOjWmkEOFKlfH/CdUxbPwkLDXeU841
TxWgnwdO2lqeNXn8ZOga3PCPq3kFcoXFl5jEXWE/wGaHx0D9HLAqgJXo1OnKsjzJ
R2g9mY1O9Yj0DI+z3Q8Fvci6wCSWe4vZjLR9tOwAhl7dlrOlr3ucvmLSjHeEcstd
ApLZDWkJvspgZBY787g8hjW4mW3ln94cSZ7Mv/w+gtf0US+Rpt1PrtEKZAr8T8gR
z9IMTu55LV5kpSQDOKRZXoxYTsOzGjmn2fDagJMOx/5De/Pa4BmNJM61dUZwypE/
mYpfvKdcJlYa6JW/4RQsTe8Vpy21745ppy1Zxl9NUoUS6mhgDdLkV9d4VKNKBQU+
jeNmr2EZ/mua87xYICImvHY96W6Tg5r9jHv9olvjt8e0UWqGCqvwA5Du60v3j32j
TGLDZ0I12nKOsTFsPIx5CSx3YsRPgIBVABJ/IYD7sGwqWxy8PSJlZfmpb3BfSOEI
292dNrmmylhUPUrOgemT8agqs+/IvdRbzOWljcc9KdWc8b+FgcwsMgxM+5JjxxuN
j0XkGH4BeLQmYrFjy72ZK66ZX82WhKNjoc9XjzEOlbpBbA3aBnEvw9tftGhCSDYm
G/ooXpRIdTTBrSjtOT+UBJmWck3jqUKSTNiyHKRIXl2f+z20U0GEEas4l7IxZ74B
j+BxdE5ythGYvNEXIo5bK/UBBFiGvVC7QcsLQvw85Kseylznnqg6rPK+NKnidseE
7st/214PcHudbuWUpnUjaFOA4Hudok0ygxBckTsG5/PpXcQNlUo3jHruyfsAX+1D
Y3uRbDHXn007ytsW4G+y8XLG3VIPJTYAZniudhKlEY3ig7ItWKFZ9KcN8Ukgkaih
lo9rsXOtjCtE8f+aRa4IzKvdA/1dzIzIudRU3xZqm2R4oAhwUkOgXifexS2vT0UN
zh5yEaFTsemhksqXwFUTZGiUMGX2Z6NWsSfScAMhkJ40f5pqO0T+uMKYx3T3S6ER
+qUVEnbtWVCz0uVjSE2fFgs/tgLFgTcJitmzh21xvzqA1GpE4Tl6jHSQjBYoY9Tc
0Ibf03RC9sBkh1dIxkSEkE4PQGRm+phZqiOSDdLqtR8scj3xOwgbHbSlnY5su3K9
mWqZrVc+pimhna+pILGg8EzxPjoXUdBwTX1AHOKdIQmzHgawwHRBBVeviyDji85J
gVx7NlCOz3xPU6g5NrVaM9ot93JvzExPXqr5ytRbi7hePhCNgI2rrq/7DDPeNeM7
5eYawL/T8MuxgPvNgfemDoyWDn8kfEBzA+Crk5FXBIJCTmOTxhuJPnHtcWnbnt0t
Nf+4aPRzvYHmXyuZ9vBKMjM2BzORWoYuSdrh9k9aSAKYFOblpV8WTa4jH53WUbJ6
SWoEqLc4miQn51N1kb/af1U+YSeVfMw0OVXtTLsmbob6+k9h21/EnKLCzvyu28PL
KGXbGIHHpGsMXIy4pZQv2o2SJ0euOac9l2eDy/3uIbOGJvAN9S2IEa7yUBjz7wnc
ebPh4m6/+3LhvMs9RPtsLm+7+t1XSWYgJwJKXuzkW9xMjbn5eXH83LPSEGm3PJm+
Na9Pti6NCuJVVZNv4aYa9Rvu14s5oO8hDnMxiO0GVqtCv0qIAN0bQBQ8XNfN/3te
O9KaZq4iarLAongPUvXvLmd4B7o2Base7PmNJ7DtfdtTQAKSg/zBJsYD3wEcrxoh
BTX4/DwKwQ/hKwWtjM3FZfhzlHO6t/aDvrravTMA1ZfZNezZrCg+0FISvgjYk/g4
otgdxN3eLzRZJ8i/+F4fxO3C36Xs26F/ajX1hqwqYtCU4IoBYpxd+R+kiQK3iYHT
UHK6fVRL19cJSOQqPS5qdn6139ZQfdcC4ZSqhxSmA9vmCNhoHQlh6EAKjZdd9+Ug
owM5NyiNs0vLmjvRyIgDyf2FMMoKBIbTasj3pZQMVVc3YTzhkQDRXOdCT6e8Ohn5
fCi1Q2Zxx6xkvzaZ7S0h+cKIghYtS4ChnqiRUIzQIbpaTwI0xvJSla32h67td3rP
Ui8hj8IHbPdpU19MbBhbm3UxEadv02ZW/PhApaflaK5IHLqBAdc7VA5d8+AXjrEI
/I49aMgWp0oktuNx092Lu0vJ5EEeUW3Z+uhJj63SCNK6/87k4BjhX6U6KV2nui3G
oSotTrLvL00ndOYahAXXcyj7NL/B3a4Nz/natvwqE2XFGtvGKgm0vXASB9vAPGy7
RFhtzhx9K3eLw9Cg3ID8rxoAtritgo/yFnZzM7U0WfSKpLvMYlBqGylJ7ExB+Za1
ER43H18IT7JFD7Ji7YYlRgbvfJK8hk8TWxqyfTretYOaFVDMoNpArK4vEbfzEEut
ip9AiRG7XUfpmVs5FV0HL97YkykVvngFZRjGmwvEhGA2Unyb3aZMYWfnIGELQpwR
TFQqqNIsNcUqQC5iR7l4FKZvYqSfzmg1vj6K+8uhNVorKe80hfvJZOgjvyssmnTv
iIKIhHA4ltf3hj0jtOfmnNSyHqDMc37NHvtFtNT2jfnd0wutUdPUso9FxYURqfXL
d3rUCM0pg5zffeUcOm2o2guHHBVLcAwEG3izdwnO1isncrKGUQbKhMknUDLOMWA4
1LBXW4qyaBW6awuRAaRHLUPUnoUp7CJXr6c9nyfqxXeXfiP33lrbhV/RvZI/RfR5
EAfMIHRhMh0EklFOqpUaA7ai0cxF5QC0aVpUKLfUEcTtH13D2DaRLKi/Hz8C2sb1
R033Q0l7z0/t6IAKbboTqVsqAaI2LYjhaL0NFcCKw2Ozw2mvbp8CCs9zggCxx5iK
JAUyAdKcrslYUTxyDAV0yN1d15p+3KRx6f+8HWi8kgmizu3bEcKYEjtpGDN201sO
WS/mx+guOeMGP+ZJ0sxpy5veKtFW2kBQBJKhXmQ38ayItvITmO8YBN2ukMzCnss5
SHZKsRQy14FAzSBBoWoydR/f4jg2WFyBNpdyAlEGVZQnLrndK/rfdWwMnwiwYb3k
kfaIxB+tLAmmncpzgvU4+dDGKLcTveHezlbjzZBkZy/hiXrpa5XNJvfxIRlistPL
LFSJLqnds2N/kkhZaPSZvM2mfbMLVQRXBKx1Xlz/Asn46WdoMBS88oxMLhWtWwwJ
SCP4caEA9E/N1Seo0kmkcPllJl4rpI1mk6yBexxC6Ij/vMifUsK8G8T4PlJF7P9N
IEdGl8ejqi1Vt1Sh++kSXnxIgZgNxY6VFfrQTrPANTxYagWYFoMKeo4gFoO2TBz/
qa97KuMj/hJ3thWk/dTsCGusE4OX1EfW4qknXW8zqDbX8PbNsqyrJ6J/dNcWTCYu
STJVR+5o/PBot2tYndqKDrw+oSryR9ig6r5Tqhjo5sjkDDS0Jexg2D+HyeNDUNb2
3vFcv3RxCSL50dE2Wbf7PtGsDy55PMD+Pn2wkm5O7DoGYZzn/uxtmopbavRsHbjt
eBkkcAnV9IA0iSYpKOrzC2xlH2IiZNwmnnS2lKowvWFqjkMQGOzp8LDtFnwTRlto
sQJHGphPObcZDFA3cCIFcUUovHnfBoa4bYJyUdXH4AgtX8yeZ3newbqSmr5DoPdj
chLJX3SSNm1zouEB0Acp8DdlKsy66/NhUl7UobJHQIvEpjwYgNmE9fHL3twaazmD
/lt7e6Q6H3FAkaCoyo595jgoeEywuVjUePR5tQWNQvK01ubRvzEUtsnJwsVkZtUW
b90BZcc1k/Pz9HVWwCZuaGT0oJ+CS8L4Ek6oS4t2boFlRpoal/+4DsNE6zwWYUhK
hODd+G9ilUeL6qC4H7Aj8fuHKo4W1yxv/S5Rq9kGNc3ST36moipywJmwWnltFTIN
VsfGwP/48UYX8zELDJlVdG0rneKLi8K+5D74bTeRWlExuJuDRIjdj+a53pho1sdj
qQGPkDFCfX8yw0dzqS34Pfn5y9NYCa9BuE6zy0C9Owtyg1gtev9kyLS6hjeqFkpg
Yg/dU4G/oHynEzu4VyOLEAjmTmPPMDxm9NslxneD0SS9SIqgU2NcFdwul1ZXcwda
eoVCYgsfkMB8jPDJN1gW3/CV8sP7CWfAWVyg7PqroN549+Zl1NvWrLr6WU+mwPRb
vb0TIRhueTs9mYoaSaLTFukIe0wWcEWMaVoaf1+70qi01Ph3zni8Bl9SzSxVdR1q
Pj03ZhsVdp0Vm/K5TitqVnMzDPyrldMwIComlmzCLyL5csFRDf2BOtqzk5PqmiFw
vpKxkEvwwk3bIoxgQIFxI+iJSX+3kq7RNv8kz2KnG6yg9xclPALuY53tKYSSuIL+
KE2tZBUFCkvCSzQ86MBAcC4g8+kA32N0zz85qG3WbanPNWDqLz01dr6Vr4SSyYE/
Ac7jr0trgCv2GsSYHGS49+AF1nDu3WPUX3l1dI83ViVOdxohucM94CoPOZwAT+FJ
Hb2UaWKYUw0IyXst7AvcdU/YViF8pMd3pVo96IeBzk44MUUe4egzBSyGo3pSziQb
X7KFP+QwD7T0suXSJse1SwFar+S0D7LhNNU6rWEE6vF9ytOJMoPhpqDUjZf9Qnbj
gSihutQ2xl2ud6aR1bWHowuDtyOStgbjWXkWJxUkGGzttFsKPLUzLLwVy5OEtQWr
NifI5KVRLACDkKCb79+F7jG7Atz40IFPYqwDtdSG/Of+bMSJWLxdMbVJnSMeOEB4
vaO+7iZYUzmHlwElB2HOzd6rtV+sRfCdU9mD9ggdRxqw9z9YRYGRrh4rn/RPSCHr
IsX1Un9Y/Gn/o9j9tHg0IIA16EKemlZAwFEYreypcnebo9w6+P1kvtqPWQFilFV/
zPUxdAHfUhap8sFJfTTqQJxY0uIXCW7fzlM9rr6LFZ3s4IJwFm1nLMuK03eoJ4tT
HR35WDXAbhaxr5BWXv0fyU57F5cIqm2iE9Ge8lDIN4BUKsuAMwzlN5XBl6IpX0EY
g4Pf0d/lofjcdCnah75ict8xEhiDaY4jgwiTRPLwmAy0/dbNDMQ9gxrP8vjXgzTp
VMvfqQT9Jw2xaBfLgGcKMl4rlXGaXRXjWG4vqJo3SxQRc5Hfkgf5gOl4/w5ZlLO8
1rTED3pyvceOsIIk51+yzH1E9HoXkcy8gYRg4w47JfnnJSYL3mL/ZFKxfB9tn389
HOYGYgy+A5Uqy5vahTr40NVih6lZKDVbSg5mUlOKBwyJtvl7AyA8qQZRVT1hgteQ
PrLjBWIlJqbJf+KvgkHq+7LyUzhy5PwU4x2DCt+ML+wPf1LhYJ4UHKSm+FmIRWFv
9BMoF4al20jYfhUOoTEA7bYG0fRD0aUePzd8aYZ032AUx7xh5NE5gur9I3GoTU9Y
aPvMWohIbfbC3RGOhpC6Zb9/Gkf0T4H9JpHfWtsNx8IWXlIfX/HUdw1gG7DO58P7
emgXIOS/0pvnijpPykz2zSNIUv5TrMmchiDjn1Qz+9H2zr1t6J+Yu+K6OqE55BR8
Ho2uTCi4A3d3FZ59Qh07qGikzJWQ5S1S3emCKJZVziV42G/2W1gtFy+YhatvESBH
wAqG9RYa7BPmEpqx5Xrr0IWbtOX6ml5X6Okl3UpspF1Fm0on4eCoIqFOWY3r5TRo
RUhEL6SPOo842TiQQeQOoSWwVnLB9OhSowYJyD7/8yz9pIQPJinwYpT0WGxAO9qN
ZNxzEC2FMVTAMOASEdPGIsReTZJiDL7o1Wqd4ezLIafxSXbdJ+GF8zeDnQSJbirS
ljBfgqFS1wKCDBN0+Yx+sHFDrnnNvf8EFLERQphGPimpTPar60EpRAmlQq652l+Q
k6CBGeuqbHZGGQ4wX6OYF2zAkQBQWDVlu7oQVDqO7otHaEE5D0gjohqivTyuK6Vo
XVP+81wZzcDIWtHGg5oijJQOIdW37NY88rm9tXBwuz80jRQ4FB+bwoz6aDLMVzuP
aXzG2PDKSXuS36PweK/MrroAsIQ+WVYYXz2ScDiPcj2hH5HTeqXhsAzTRqpoRe1k
aoRtgXaUJ9nYvGeLMY34ISQku8uGRfrp9v3Ni297PO8JB4xL/GePBdTGOZ6h6Uvn
4PNXAtD2YLTomuUn3fpVlbzrRlCcqU+Y1F2dT7MGxVX7pFOTQYCuz474e8t0ZrGN
k8qGg37MKJKAUn09lbqpo34yaJpMCCIGWeMhBFXpMWmcO2YJ8ttJibsaP95SU0BN
srKxOCu3e71qdKGROoWS8C2gjbfmXMh/5IwKWf+z0JONBKfNI6k3ZptPg7v5rnjc
jRZzVhjo79nQgYJtYr3NDJXRme1stGJ8J6ln1sPxh/1Dy2P4lBiWAPwAy3QXdggy
Xg7P3szSzepNc4Jy+4HY1mAAfyVrnPyGcWTJjzC/zLQsTlAcv93r2GJ06Y/1EPHS
jyFP5LAc9159j22IC9LJbjEIjAMVqHufkwAId2KO6wyl458ImEsRBxWA9iqq+YoI
VaUJa3hx+v2WBX+9GZS0raRfbtm1zPUYxoT72PRbzUFw9nHUNmbfnCpanTzi13wL
LzrBTBqSM+PSODpGKP/n90nusmhyUmWBkFUfKEUZ3zkrmeG0468UwfdRspycVreh
yNI68xFwcVHEFDKrgw1b2TtlsrcESnM1RzoAJwQavlRY5VaG4sI+OFk9hfxSVokz
UxGFNiZ04aTRhVSS/WCBp/I1LH4ZvppjTm62tL4r7E0ZcIb4NMlLOmYwAnOpNdCi
hrPSSkg/ruzeNMci80upuS14TOnoJcb7OC0iRmByM64OkyZACGsYgr7XRt/+HAG0
0bVWZAw9g91dNIDQkdenHGgcYe1zCQzMg+1t3YvRLVIM37F6gG4sY8bdVvDaH4le
Uf3Pk855fsndHZv10NLopcOB8JLPYrbFMv3UDZqJetacHZrWnHk7UCqJ1DMmaMjk
7JQwNq8q8lDfTFoq0UUnC1rP4gnUsN/3MG6o9mhGU7potiSH1sCe8bylb/D0LZ9E
KwHmFO/xrJ2LD3j3Q0doTbajKF8f3tnxsg8+cUWAi7dEYNnt0P3XPREetpEe+8di
unwu2ry3nyvfAdk22nwkFWmi/CN7rx5i1Lgfsh4zUIVjgVA2unJD1DBbIlLn+mXE
s4WTPJmIdQg4XfYXtVeRMzSkjxPnGlFniIUZHgJm9T54LU1E7ki6ZneVNKsKEGVw
/qHLT6fv2ATc+X9akzSKRQ+37OadWXOzuPZCNh/OU9+QwsGvkx90e7CyeFeODbqP
4h9SpDLHXqtEobt9qcBmlKs4bWqtRD2NfutxtJ/uZg4raiuune6laC2VhhRqshb3
/OpwYsuShNv+YyPIlq19F2FawYSAJ631e1hWl7tuoa06jbcOj8NgP5nY2gtU4xwf
7BJo8eNxAHtRNX7ARz1evkTw4ShN7++AMdDJlGZM/iDRYQg9RpQiZAgspAWQ0lYb
b8gml4p3qVAuakWMjvToqa+CQRjufXGRRCPsBp5IDDs94U1KbW0GjuN8I3i3s+kW
r03h9CMA7ObHjata+qq+wbXYJhomS8sHmkMbsLZgEbfmFwhYbYuLF5QI/3W//chu
kt2t3DlAKxaF+vLNXNQ90CIShxAAtCVbfrqXYzPgsojypVieR4Swf82eTvbWEtAb
EBdZ0tm03LfM5Ba0RUj3NWiChPP2VpOkvQBCTL+urq9oBu5ajyv2Zc5ACZxIoryV
Q7cENHfIt/xco7kuXrz7Yqn3crXSZgNP/ih0D9xL70tmSyq5JoCk+KY9vMmglpZ0
1OYKVPQo4LOOnF7DUMnvhzeiGOcX70YUgCx8L+zs26y6Z0uSBcCfMp16aygTXffu
vH/nWfEDZbehGLjzOPdqJEkqO3q47Rt/Un2S+H4hO2wx1S66FySSlkLOqwE6c46s
MDz/km8DuXT/sGNqjsaTVKsfnm0jCXIb94zOlwfCEWkMpJ0YiYvy+/F/TbfIKRev
knc5Tmb8rSIX/XXRMP9bHb21LLhqfHwJmH4N7OXRAcAb10OFUfRc4HztnANcbD1C
6RVcDgjw+to0Kwvn/yJq/DjFSC3xV/meUF+Muzs9fp6vB16z/v0Ad3auFo4Nf+AP
dFWr94jSYnW27gfgSgjg2m/x9xduzX+fWb/yVSjrEBsA+fC/J4t8FnyaUX5iUoFr
WBLpkbogLk2L2JY5vgWQxdgdiiWAxTSAsCG1Xxf5nc0/0hzASSOuQLFl6rPaLefE
QG4iUvwSv0UuNn9P4zMGaRioGja2T2kGQz9E2dkxj6x26dW/5xcg3k/OzdZhZlz8
i/qhliOBe7G0tem1WaJxQsw+UHHVYQ5lpgWMsldnsXfC8cXW2G+pLy3/ZZtJkxnU
maVWWbB135q0JNCgoNrLSesOcdzfA/Zcm3Jgvq4aAa7M6q6Zvxoy4zPH78tUViRZ
jE8S23Gy6hBR/xPbYul1OqrWIW/m6D2+PUb07StQ2ohnL5f8v2B1eYfahaGwv6lG
vWNmS1nQqWQx3j+4R+CgfT5ATJkfYPVxX2AzNXTFNCukrBH06B4PlHX9+NN6efxo
1Iaw7BKiYzyH2NHfPt3jG+npn+LV3jPG0d+fwebsHl6Twk3dqMuhyi8OL0GMY59x
oXvcnNo96BUBFBoZ5FSpf+34stPFZVQ92OdZu23ks1ICOVVJWPXZzAay3S+rV8mj
DfBOH2ZBxPEKMuWGbuU1j7OfSlr3NFTju8SkLvVkRIGkWIey0B3R0AjJ1GnenHUJ
RrSxyTf13zb4XF0w/q99zn0UQ6rP4JnDVGO+H4h9upAwCAVQgn4d73juPbrbaOFJ
dbAxHHkFsy3H1hz/ZLVp6joRyeuRg14UwsT106YHznNMqwXldPwLPsZU1jiDQbxf
0yIiK+ok95h0jJ8/hj7j2jKq9iGSDkZWHbHE19kr2NXxg9ztNleVhS7SE6hLu3wo
foVZ5lVgsMpdoxfVQHyQo+Woevenns/CC8WwOtHtCF78ckZUadkBZgbP/sgl59IM
rrx5NXZTdfvSbDqglciG1C4J5/H/x1L2uE565sljiL9XsREmzm/zhbnP7IIFDRTf
NRR7fPrC1bxAdWbsOMyYvKb2C8p/fbiKyQsitjFGdB0Jbyua2Q5V/p/7ocpUASV3
Ya9/kxdf9znhdrvF0xEscPPSlLaDTupjUnR+W0lIRm2WM8dQ76dMZ8l9FT2nRVxF
S2/Nk6UE3DMll6wkyKVNzQnbJEPfzZ0B9kFX9nQAOoOrVWy3CGu1jdZ0Uef09JJD
COhKMGbP+CLKO03u0Lt0gt9C+NY8AFRjyVxbw4dlHXx4kFnBHdvrm56z2ezhQ3G9
kO6YnEdgHBNWvAbVnI3F45V5I3fcdv3OXy+wLpeZUUiyvj+E8VfG7rBgZ7f352gC
gUSDtcp0aDJSeuvbIUrr2FH9O+KtQgfS3fgGHsmZDg4s3dJqxrgPRsz4/XjhbLRi
2Pqam64gqXYnOzmGLCb8LCEm419q6FtQbtliEHYlPUE9gDlnVB904X2u4mW4Rwl/
TO+IiWbt/3CaVU1ZbyYSYbprGeXU2jOoW00KO2JH/nY7aTU/YnrptJzzYDQMv91p
OqmyGOkTDm6rO2Ir/0oIY/HNfhIriQoZJLt5mVw+4aJOYqMR60Up0ypc8DbFnoJN
s4KPZf61girKEnSJncsFi4mdnIi6hvPdMX4cNCVyIi0idd27trDTCZAIRthdIG6a
nRuvAoVPfIDXUVgOagAJXdMuramyD/w5HWPr5/EkItWrgv22wrnS7ikG9OHWkJ1T
jHOKqSNI9OtszDsTE0GMlAG41rWY8DhCJJJ+IifEZgBl15/3RMrDIOvf3YYk7oJg
4JZ8t8HxxklYN4ViJRpuj3ZZNBaapX3BU3pG8yosPz7UkTsOIYOD6mYZvhV+Vm3E
bfzGmfEzbBzTe688PlieYrXcmUEV8PrcPFe2OY3+pKL59tRtNhY4Fv4gbNur+FPb
0lQ9AuZNTAXmMtcYeeahVZ4daxbiJZ7SZ0uyJQ9SDASAsJdyMFlYusOm5dUkiLa7
J8n8h29E8M9T6cdxABT6SnTs4QbvXqn3ErZ1PU62cUiFlVFYl+VoR9R/32HBTLCK
xp1p+u1ulNTZsoh/TAgTUtF1laKKSuI4NiVZ3rM6f9MlgDuseDuSZrlCSHIeNTe2
A1ynSQOpB8JeGqmQ/cZFNVpuiqZ6lBoZYxIWy/DPAVe+pdID4mha59TziVgQquum
audc7DOqFprU/VpYjPnanlXFpVUXN1/qCrm44fnb8zPuZbDuszcK3ls58apKSKsD
/DqERpDBs1DLAJVQyZ0ejH+LmWFihTUwFcxxIIXYB2/MedgVNsBGFafbUx0F2RAQ
mLeDFh0FcrFvPsdv7LaBZVTnM6zQTf6THnQOtbuGFelARyrR6415ZMm2CeOPzItW
KLpP8ZnEkuCR5qNJ9ZT3SiuDGLUbdawLildVfln36TjbvUKx7ZehqOeHAzSJ7lbA
l+YYUVKk88KA88qt5U/SebVECoqxtbIoYfPCA/DIyLObEcAvxoiJ1+mRQBxIXWAa
lYkiZtzOjml1t4XwdSmpD9zZV3JfT5tK+e2Qszu++hV3wW/u3t3xV2im5ODKpKhJ
jeqVlSPI9+cu+JspC1asO3MgcJrHtp4+T1cJt/YohtJrb/db/uiB9YhlUtl3JdNX
fFHbQInKBHG3qkcmFdOcou81uCQ3mno0CiF0Ql7AL+dlIjvulYULTBqhbgHQ8JkA
M6Y6U2d3kQWXNQFNniCTBLodjG26jNWft2Xz8A+1DEvFjjg03UBaIrJ/gTjHBLc1
dAAbouA4w60nIMBdZvjnY6k30OzTrWIyWk2FVumTpZX4kthy8MyOe+kaYFZLKmjL
Me/cMeLarKYu5Znynf46KCm2UUrMTUbLFCRkX8270F14Wg9JMZzLcR4EnmyOc8dg
fj3NaFpkYztJNdYQST5HDM19gPysWVxsFQVpB6vAdkI9mKfvEhxB+wMb5PWBfkvJ
0q0EbbmKC9xBG76d/i8CP5FfP9zcMJ1ISiY1kvQf/pzMGiB+VM4hu6+orgg7z1tN
Gdxvpcw+rx/SxtQhR5bdrbimXk6L9xZ4IGgqMcnzoCMc62VfmCrNSKJfWv/mCsMU
kyw5ZmpufzdmHGVIzYbOZko631qwq/7GV687TWGp6nvIVQr2mLq05iOp7bu03sYG
QnZvjLQ1UvdRVHjyU5H6jfAzkYiexk2Gu4syiu/m3zGPOF1Z4UTIajF0FMDzE0gQ
fWpLSG3FhlPbiemHTz3/74nHeU4vJoLDvfhQIyi9/R2CVifB0BC/tebIeIgRJFzs
fm9M5UrW75WIJNBiNoEEhK+aUjhrD0tV6pR8ux8si+Es1t9egPgP5jZkSaaqVwK9
yDj1kGNblh/mO1EAXCJr6ZYYZmeHIr55rvmIYOkYtiGwF5+dvHY1rFmrcuoDsd4/
DkwF95Eatksr9DXOeINV0KqiQCWxKXwd7f+qUNMIcIrv0aKuKr3iijurf3H1tmlw
cv7Tnh2+cD9yrvrVS1m08P5HMh/3JMoGFwY1lAwkQOdQORmUTB26qGAcy4otZNbZ
O8F1tjl1vbKChWkUleGvBjzPZBVyvj/r6uY8jzd89vUluM0tKIhis7+WtF3H8Ibe
bY7hCYtrxZEAO/sXTruO+lK5ZQrc0BB4enYhA8lLKbI25WzdwO12KP23lkiHXZKI
eLpdOBd1OmAk0EzySkkhDncMsQBXlhsbHAl3GmrCsdJ7JGYvt4UGxPcGV5JXG3sj
IiiQU/Fwz50xRMdLVbOTArh/GwYjhHWrNnWgyvH7MheqfllJnCvbTF/XPrYzcAc0
KEgQwh/dqV7QBLGqwPYJSPKxmLAzbJLu6mqmpc5+hsDjmJBpWGW4yLLRkrQazdhR
woXkCT5dklJI/NMjZijehRQYgDhAt1/IzDzMK8rE9SgMjmOGTcGfDsdGBPZdIF4u
OB0cx1q9Qsve/23BIWoBCUuculWe+5MOI/yIV8G2HczEcWjizXz7zu9zNIKGLZOp
Gzpdy6Ei0DFWjAd4AoUVaQr6rd+AenDZHRLY0lOyG/UFmEjZ4Cc2LWGBGtqW8JdD
bOKJUX91Uxm+0jSvUucFR/phBI3okhKwtQyzn3biyk05hHn74Q3KyBLBLk5nG02V
3qqQsF32BdNv5fHQ9vK+6Wlg6oJ7MRtetyMWuZa/Ml69F8fj9B2ntO5YIugcYXbw
/qCv8u7UdOqUslNH3E/4GCoWDUkspQT/6bC/QwqAcPaD5jTJd81nKePwM8rMfZdB
UbQE/W/+s5Q3T57KfrDQ38fBrCD7pgx+9alIpT3+uryVz4y5LiajYhJw06XpRV9N
t/zNvMYKAE5CPHWoL6tAGS7p1XWrSQZR9UqyvefRxU4rw8IaP9NJsXQ5zrAZuUNK
6gHThOsoEwHvO9kRbYSfH7wwzwQTt7KgCTHozoshM4HtAjexR6zKR4m8yepLgXTe
LvpIxtV4kMkalocmOovnrrNhd7QSebjEXsOe7WmJ8mHX0QCekpshySo6sXhM7cj4
kKPPqOP6btR0UZF8Bsa1bjO++eqU/NGijbDKnDYGrbU3HcE9jVZH+Q23F8Jh7cvc
FI7nMJ3ylLNtBbA2Pt69p0EV5XTYfcwOTwg4HKsf7IIDGsMFXqjZOXrSMaSYSEOA
pFXOEnIc48DS60dc/0i+0gUIGgenA6iikZKtKuHi8S7H+PIPngxRTRPhXvurVE5t
EPSAXui5juY2DC60KYq872pE4pB1mSPTeKY+Igq6sPCfSrYLN1gTXwUCzvFvT6i6
jiKeJnTD5j6Tchr0ilv9y0p/PYQci2SityK+SmkCuzvM/Eg9iLQdZ46due5Z9+gG
jZ8/d0FHEJM3BnzVhiAINvo5o7BqmkYZVRFzJ0AX7u/I2iyVRrN7iewo+tD58H32
o2NF2hHFdzuDcfLy/c6UXPZItMFIL37nPEFHsqGLtflr8ueTBI90DwZKeL+vMVzH
R2j8Rpbu/rNdGumXw06A8sCh6k7zBodDYUHg+gqhEx5FTE0Hs06QqplNPlYdaVXb
dINrI2fyYJZgvYuqpYe0KBw0Jo6vNVnwcBeVwvgSfgFeWcYd3bRL6913SaCLwQv2
cDXwJOOhlILm6xR6w0FddOP6rz9+JnPJ+Aa7xEGkrXh2fAi1spsOF7aDik6vH7ee
C+OWxkNbTD+U3cMxyJsQAXyvAOAaZwyQNywwOCvpEDGklfPTV11x3pPywZBHQ4VE
WuO5P9hMWc6w5DUq5lyHgKYRPtYN3DmgC8uP+VrYJSYoNVYk+Oe9l3Qjh85/WhV1
k/Az72+98C0Bylk8x/Rtk/0LLKb489RyQ/16a+di0k+ZxLqzGCylOFG6SNyIHxgC
5qzLpfF9/h6cUr7R4SvsOt579YafivYfCFpJsxJWnEwbPfI3GLGNi8LQsQ4rI1jg
KOQ9mN0fq0lYzTonuVTn3fOtLIKkGDGOKYKv4JKekeYhGCaYXtkHMsYdXN8kpxtL
yPaFeGjAKgZwx63jbVeASlX5qSuRP1x7QTU+0QUpvsQH5DX0Wu64Om0f1lKTu4eT
/dgEf3asukMjoLon6TDXY5oX9+YwxBFL3AhBa3vVvHFnPM8+sPFGRywjHyDM27sw
envrb9+FMiN7+L9xagGNu5E9JTMSmnNYEdPBNYTtzVHAfeV0zg2ZMPzC6xZ+YPjR
+QNG+BE/xYbAtkZ0CtjGXjj7V57LztMrA5OXW5TBqq9YoY9ewXzvV1mVlpM95pre
Fg1z0eWcXCdQl8rwjeCjnfXeAEon1e1adT+49xc9MjqTlcrNgRsJbaXF4grZ/auS
UztCVLMWsi2w20d1Z6O0CHFSnthRp/zQhpk4Km9eY8yCzWnjUkyTlo4mj4TVfYWG
StjOeRL7TKGjFbWM2UEnNoFoTUvHIWKTKDUK7dRrEIzzB2MRyL5PzQR3Zho7ev92
TyEP6YxNzaAFLdCfDEGoE7IeI595zBFUK8lOJXboQAMt3RV/QxQiBKnJPaZDOFjZ
DqRMm+GXH0grMhAzHhD6anSPz2X9xFHxMdOUUjkz2MUl/Dds1pNRnYpQe2bRRjai
ltscp1DpWdkHJQUkatwMluewCzakvMDG/HsjgnO9DhyG5NjmYUAbTxbdQsO0e586
n0OpXZ+Km5Gxi5CxvDTHIMeNGLGG4SFh4OnUyjaWOZRo74CE40PLl8e6SctIfS1v
AvKWsMpey1Zd1zzJootkxpFdA5ePeII4zFglkxu33D+omvF/CvsJHtV5uhkEBkBT
uCIuur7PPwf37ymJlUreercG9sMMVLV3iFUpNxUu03bx04M6Ctx31c04MBUyTlzi
z+Rw5o/h5xLhIRAbimnJdSWKo5mz9cjYbq97QooLLcFQePYCmN0kd88uVPCSI5Zo
jtKl5J6q7NqFfTTqzh+NebR8LClAOd+ez+Dzy7r5wqXBH+eyAmAwRewTCoyGiReq
TzoJyj3RCS2Mkkzw1LFAMbhiq47wFvkgHuikXGkWIcD65aQtZ6veiZ88VUuliWDI
wKpawSOXkR8G/HwFY6v/3XKXQLutc/oIQ7nfo/lZY75WwMIwaItANXMZJATBnw7p
yi6WUdGHaC3RHTxxtYL+a9qU1/gto96tpQFP0fFVUl4TiZcseAUjgez4uFYWaMA6
VOI9JvUzIvHhvL1TQKR10vztHcjLwRhf8FtfuRpyHITL/nUbvcTZzKxnskbNgv3V
yuQOHobHHU7MzbfOMctcbcbhbaSqLbBHfa/dOLQ2C1fQW0NSlM9uQCjtE/CAfMGB
dgpcVFrdPLIEuAS1MShGVSJygyeMfHQaeynVIU8P8SjexIssfjreQo9Tq6Ag1ZpU
QpIt/DIt1MKKev8qg8550jCxE98rANmaHLy/72CqIsFIYciZniKouR8l1U2Fu5xg
kjc9e3P4poG2xKH+wHTKajU+hSXUbWdpd5LwRFC93+5RWafFdL+AIkaYErIXeLHF
9CwYfeb7dkX05J4bmX5vU05LeMAaJRBjrYR2KKXq44r6JmjUucV7Q7PPDM/KC3yT
9yGhlTIh3Lcz5AxhNB2E8gMsJZd0uAgxtFJhiACCEYya4DcWoAxA2OsJaIT8sU/z
B8JnzIyuhq4ehYIWMygy1lHXR2G8u/kQD7cJ7U0/FteDtTpLbtUbMTaUpacIk2zo
t1v5Hijz5zSciVva6uCYYqPB1gAmp3kHKKa1FGxWUcklXfusVbVQSh1IsfumnVnT
qp1C2OQQKwISk+l0yzedRY0nUIJ1jgAMffcU3OykD0uVEqCO0hIfygMKzW6R+6ML
2CO0yTlrm4ePPrOcVqwnW2GClQUweOx0M3zTtZj+xmuJW2d+mHl7sqZAnPMy7Dpb
v4lydkHfaPBdrcE/qgZQmy8uwOEKyEXz0TAviYbg3+oWsCs5ou4bt24O4LgRJ4V8
DTiFiIpY+gF5cb8nPKYBz8LC5NOCvR+roXB9WmSpOmGqPAc/u89IKyahME44oKRS
YmqgBA09EXGiiCInGNj1RtYuzSGCSYRS26+0ZLzOrey59bSOrGPkOxWMfm+wAGiG
EdaBYdacnbxDeS8B+bUv9oYBCqop8rE6V742RnLmXIn5+igSdoTf0Ycxm3JOqmKu
ek2oHeUJR04cQkQQkqUWz7tmtxxMXIrIQ9mWV+SVUH5t/MiFJIQnig3b5DMdbzX1
jpvpykP0FmyYGYdh1ahVpAsB0k7ADN2lc0qJjYlEy3g6DIzwppuWFFj5U7a8RUFM
5Y3d2daf5EmeOrsnfWi0BJ/altqMMsyo5fhh8Ia9xTApSS6vXuCIuoVSweLWgZay
kEc/7iZ1P9sbgECuyDWGIabJvLPKVX9QiScODD+XS9ZDvURECVRsqIkFYe6S1goZ
grqyu4F7WT96EzObEDi1uw6jBz+m2wUmAAsnQ0sGQd1F4ymIi4Q3qC813H/gtyft
g1WRPrNJVZY1bTRwbXM71cHv+7tl/bXPG3Y32fvBrakF5ddnst6l5FPjV4BqXV8D
kz50SkDbwJPEieiF8SE+1p/7DXKS7Tj++9fAiV0KqaCBGbQHFs5K7BS0P2UNLTEo
ntwXCblJApiL5Jql2evlejMzqayikBTbYe3ybYMh70dLNvoQrpV/YS6Ii55E4RCG
OK5BFI8czcSTXN4Cd23GR/Raux4Pre2Bmc4jYdJY2Fo+Xn7d8ex2yUHpT8k2J61e
vtVv6GXH13rOjY458/0cPiskE39LWfbNeFyCs9guuKgtRgS/0MCuW3ptjZpgD7q/
jfzZf6Tg3GMwHWgf0JoTdNrpKHHfKjgqrN5OOO1w5Rtr8ex+Kx+8iYFIBaqlIdLA
rn6QPxSdloU0iE0POVv5C/MBkNjDrGflpNq/nztKeSAsf9mgLE/1Iivw7vFYVhIu
KVhIunz0UJBrvRLSHiv7mTZBFyKEfQgyuwbfKIaC9EeMVkdh0zb2ih7In1yqu+UP
cr9jMSZ2egoU/qkDtvsN0hIXjCBFDhIqsvDALvXcMqy+P0bNB/gqhkFOVVN+BPXA
kAkcTi59uXA//nm5ukQ1IC6rByJZ+7Fbi0wKF9t8UTcbp7VAUVQ9CiKm1TDTIbwA
kS4FFZtgMOTqmS0RWHAQJm9sYmUVXbgJX3gGrzhdB1yAU+AOwE7lhz2CQ8GzQjLC
GFQnsJJvRpK4m5lYCUuzs6uuzFu6yDcf5dp5gadfFK7jSGBZ6LuE2XXIGTXCtbA6
9Of+h3uxV/jGyWKfgdKGG35R/Ik2d3yGgYv2+KKbhZ0DFq1Q3a1vm8wpDt3afWzu
s0Dp0MMDXGHWAkN9eAdI396g3ZpK7Y3xMtvlewtW/NWKG7rDLZNgdqR4zgM6Q6uw
dbf/veFVUdjCKKM0ERw/FDIj7C5qx+2TMwMdGV1wXAQKO3lKlIHOF5FF6h5tNPJE
hef36Sc4dHEwwSxoEReDj/X9DwKyTNpM41uFpKRu3+0IkWynB/db0s5k4tcxhyEt
WMlO8SfNnfYUfDzKx9sNuySR+O7CZoDhgtZNzvEFnBLozQqGO4Y8SY4fruTs42/s
TMxQjI4tGQIZolIKSL4wYT5X1vnpLctftSBLUkdtesdqruvPT8GwBAITTfzvSDR5
0EcuR7rN5ljXYJ3Uc4WM3s9HLZSf31mcBAk8oA3olou1hCOSHxdxf2gOw401naRO
li76rg6mSlyQnJ3hcgvC7W1tcuvjpaVbV9ROiKibiOg6siOgUck5bzvVRDpvY07n
Y3g2wFWCdBH1GWum0+ljPq/eW9Uj0X68gWNkUXYypj3bkDRGFgWSebLhgyqdNgnq
hE+Tt5m4Nlu4ZxEzDTd0t0oVVkCY8mxN4R4m94sIRO6ITzW4vdemKDjgqvxwlRKD
QhCFFNE+8Xdc2+xnxS5bnAWFw4NWebIJ08Tb4nSZUjEqCbEZZcKubdXD023z1urE
3TO3eDDYMawefLRxQ2gu/Et0DvYTqDLjqnUDZn0eLmhPSwUnfr5CX5Ecz2vjQ0Gm
gjPINe8MHo0XXLVKsaNcAeKnQ68ra2HRIgY2MWcfKTUPSz0saDC21u0hRVg0XsPm
azfe9yoVK0AiXM0i4bnHOVUeSmKUff6Cv7W0WX0yEBNl44SQ69rCprZ/LiTv1UVG
EMnXN/DUlotaXTbJ2s+nH1U0d3hB3O/29fbuuKArovfpyFvFt4/1RgbDjkKL76hk
LIHKTIikd4Se9mG1tyXlZ6sD85gDgU2pWLsNCUzBsLRBMIU1tkDMpMX69/JLyZHX
4IX5v3f9kqpnM64jYMLwW65F+AG3xklzCGk0VKBn+ihPZDTmihsIeCj9/VV4ilR3
Dh43rvqtkGh/YHK0TYrxZKKcK1uLjClyzsU3jXIshccysFdlON7H+C3qT1KyWMtf
GwiVoPhChToPaQo9VJdOUGD3wQmsggy5myi0X31j9wX5WvRCm1tc4k5GXYwxZ94b
2hf1vlEJf4BY9VILDvCxey/iR5zN5L8d0huI/qjhfySj17E6WPRg0+KTuqguh3PB
dKIE3xVUUuqdCHOzqG6uWPLsiYtApPXplIWzc4maOB67iH3HZ0w9mjwuBd3O1fQ7
vqRpTZtGAo81aEuv5f3HiHp8nauZq7mzBZF30ZSh6poX9KG/M4SQu3hvb02bUbeM
2l/r/d3abAHVKkNdtEwV3zJXuhj8DlzYdqmMDkFdLb1rygYZy4zADIYg+ShJJppn
0JbdMFnurkjJtDfFg94JE4aXbw+/jTXQma+QZqtvox3YQK8ND/JgT0CQj3gw3qit
35zIN9BGq9qGRi0B/TGnODSAMt6ViWac6tRxaOibnseJcrvtMSxuEPXRdNs0FMEv
0QFP436r6terITERq4E/iw4mcDHoNJmpvg2f9V6+kBEbkk6c/h/Yc1O4whkXUzSl
I/1wbvCc5ia2nrQTE9VibZ2I11/r/hytgePOBwMKnuVRaJOKlumXO+kQykZesJ85
ovuDJnMDljLZie9vfaWLAnk2C9rCqRes45aVcf9sftCycVlsQzq5VaQv648auaLa
wtKRmPW81eY53Rj1S8QMDbhEw89UyHyE5klpYaG9tSL/3zkgfvPv1Yt2SSFmqxEi
nrMZGngNA8cXCZHcU5Hi67tDgRQLesGqoYWiRMhf46jtbaUQFZgaGSl8L/e3Fddx
wGhr6WBl3yPLSlS/F+fApbSEw5yKCT6XfQmbmCn6mQT6YaMCyv2CvYGsiUY9S03u
V2HYaCiHGsG6CWeaRcH+lKYWHjtBkLVIIeSwlTL4AZJdwOIVRN3iKZ4TJFXaZos7
1Oh7NxM9oHdFCbtUXkLuwbOY2YMzVkx9qMHup5lQUGmUuF7rMsLMdvH52ozJ7kOj
kkmwUfdBZRHvo+XKbxT5vgmrczWRoIPRGRLUfGCAF8FBKDHoBb9Bw3+baVzQxBxj
pGYTNF/rsljq6dm/kTkuAognH8Qm6xc0lSGIUjNiJ69Olmnz5sYzbz3QzfaXY1DL
m+TIQsv/DqOtqQG44PmybZeKyypqI8NhByb9TREanWJAbPM6z0umoExPeicRhntl
l6/FOB2yxOEojBlpjELYLOq7IAkXbM4x+LBRxp27+jkupE8LfCP0CM0MPRLjnZb4
zWvrLhXwD/VeyfERp60ltpftdtov8Jel7AWELVSsXaxUyPcMBqzQN2Ea6fU5hm5k
DrKXoEi6yLv4DRwe368En24anXY4TipCJBVNADjUEWABUdTA1R9aJl0tqv+xnvof
wdWgJDlkziVoEU6VXexqD8/T9rSWS71Qd0w8BgJUndKR8GeNsdVmHG4zNvEdQQCp
O01tChpWIobfTCXTLwiuWJfmP1Fwa2wDa5RrjNeaUouUTO1bJsSEPCYG3Qp9oK1o
3uj1PqGzpx9jz96GoVN/N0TaU/uxSWuvqlR2EW+G4Tg0Nud1f+/utYN0QQXMwj/z
NCmQ/cqHqmsRaPyvdMNhm9dnhzBUNdKW3I1q68nX0XccgY8dMDKV2pk41Akd5iNZ
i2YItp/D2k5VNaG25JwTDke9B7TRDcY9yzXRyiTfpSIWdreMiH4uw0F0Fkpn0E5K
Rrr53WNYTwG7b7kNh5RUEilS/0zXfjUh4EK4WogVN4z5X4Ogwsu7K+vLuv/UJ2/d
Yg0OKtncoreYBpK61vjVromGcuXhx5KdoW2JIUMxmsUr6c7qtpss3Bq6aUHRjDab
b6a4ccYgqSGbFvxjQOUwig3ni60jSmOZKBuLxM9KZbkdETXrSo6pMxk8JMYp2gFc
cQqDSFM+03HAp9IpsHph78IiFFRAYPI6O6KNEsOsVZeCfuk3OJnRnNyG3VKPVPO7
O7ubRtNLytFMu9VVvIFpkYAL0DWLqmH4gy1mUWhpHHXK7VzFibG7+X1KjacQyteb
gMf8W0VDnryO0iHp5SQ+f2tDdQ5ec8dADL2e++8Dh5mMIGZwzzcoKsba+rB1bgqo
nveVTQiyelxSlbG8lxC9zASsBXoueYhLZ9xgRkPFGFp8JpufEqpNPNAfEpERDTTW
8xtFgu/wa/PR+8RXcrfrPPYf1WLFFvHVG9oFeRpC9HxwOHqkw9/7W7rh91o/5Xgb
KSQmm+0PFCTaSk4bMAnuUoeE0KFO8Zux2Z4+eEtqNA92K+OYfeyFzDHBDfh6RRWt
61YDQFU+Xk3HWwYajBfByOyv2DBscg0Bq4HOI1jP32hwW6G8JPV8tHbHbtWOcGTK
GQIHaC8g40HxophB/iYg/tMh0iEbMlgcDWOxLBeJiuvWMaq7dHcRizdvWFwrBOgq
kzp/hCJ6Pu8wFaIiuM3JoELDZLpYS45VpnIdU5HxiQ4cD6PCBXqFRs2xgU45pUSB
6JfjvhZ5QTW2/DHl8kJtIYTRRicJGtSa50flGcPClNOX9GD5gM84MhAY4ON8lput
ew0r6EllsCw6a4M2O3KbU3FdG4TsdM+5VlED4KjnerqZX6kHGRbSDFeTPAKlpmLs
eLAIOiQ7oLOaQkeWG1Jo8VaUdhzhyS1xiFmoe6E/obCCRcWtpEAHHI7LHHKE1X6l
8d4aDxuF5PDM9az+i960sYC1t9BPddJOPHjLUOOAFniJNAOF9LdLV4pUqPLlX+iO
hx371t06+4ia19tSgdzr35u2i5AqAgTZzRifsRAGlgssaU8y/6M6uIDYB5nJ8hWW
uuh9hRcB59SpHAqR8MgI8FywI+OYNODHzXQD7CpIvEgO4cTjAoLBBzZhlaHyQDra
O5t/dRg9/noP4H3TslThxWz7ihDFR97hLKlxkKflyhz5WREdvf1hJtWfRXfJY5WZ
NboN9l5orffrEXIp6zSglTVTqE8WbGIe/c2ALj9fxOBQ2VWR1W6+xi8CIubc9wk8
vKEScXieHhssKBYqGXdXnEPDFnxERjlAlGdflT0HQlXNWiFl/Rh3jltjh01+xYJm
fn9/XGEhxoYpy31o0k8mjeWFh0gTjq8Ig4M9WulfmlaGaMu23Rr0NL+7lXF5uxnz
VsJRbuy4kbVBf++/BaYc11QrQw1gq6+wMKox1Hh0MU4vHW7fWyww4bKF5OZQyMJa
3sK4SMcKCQOBaatpb91gNKZ5lXY58n9JuGQt6y1KSbrGkgrOPq8R24zmH5+96O7w
gfDaSOlii9FQuO6rh6m5EBZe2Kng066yYyyvvQbxvFISMlg2O8b80oOqiJRGn2yb
HS2XeVhak7kDjvcVSgXA/NxoKKAR+Ck1P117dn0IaTij3q4Z5UA7ZIFZ3QTyrI3p
vStzDBCcXUU0iEPh7yjsLVuexIFPeoyu8y5c4akeKUfvjt+tOXRZtl/fwA2wCt47
/iJ8VyiWmtXxZ127aWSKlaJ1tl++u5SZwrwEYmO3E5STfusa4IZxD8XrkSiy7rju
72PiqvGtM2WlbeaQ/tqyL8m9EG4bGt8VWxlXg8bZwg+tCWw9VhzSBORqZwaPQv7k
Eq5+4e2J3+6q61GW9vD+P2susikKjUO5OEAbmHACkYzD4d1LyW/v/0Dy+mE/knGJ
6wnuGw2ZsC77wIDcvb3RBsvNAJwfQwcJ+9Xb5g6XIn8A07ByHxnlEHpLK8niLf9T
VQcgFWj4Ir0kc6wctwQvOgeK6MrExP7w5lZ2BIFoDy7T+H4bvc6ZoAF2B/rMHS38
aXk6OpdaI4m3owhxCxU2UnzFSNMFDfXdhnz8Vo/eQJFqHgeFqCtgJ+I6e3Cw1BDe
gY7veiTAs5gH6EHYQKAkmc29mBsdT8ip+KqmYwJc+5ZMWszM9R9L71TYhryJ2Hwu
NgH85BVtSX+qDrvpSaByceODXSZDN+QYatY3+yA/DjPStHfdfgEru1ONR+n6uaef
p3upn3NXFctBCHQjT2N/pxYwuAWOKQQkO5o4qQVGEqVWzJOavyKkXhFpKgDEUQxd
4aZogYuTpoVjPV99irGCZPkDir6Gc2yX5QLR3ESbRhgPTa5FVBtQjBDVqrgfFEac
8GWlBJWZyZBJzRfGYFIrc3/7dznNPeTPVzadBFFQd0wQwNeTVw4BJ6u9v5VS6hub
hg/B/NZZMSiY0TCEy98IeoDkWBR73rWKnIS92faBig0hRi+7w0FDW1FJiwFlb9x4
m0H1JjzsgxDWAl0BJHEL45Q7aiFBw6BOVMlRHVjQNKCuJclu/YzT48pSa6dKSIDD
KfmEbGG1j1byK9pYM0CuXpAjpQdh1opoFZjOHsOfOmDP6lB3zY2JAgE9kh/UVLeb
hwqubXIGWOBe7mSQqPEN/05rWpHudsiYZEB8Rvil0WohRZtkGi5l/RPmiA7wnRs+
E+99W3113HXrD4s+IrultOnhyys3skiNQXocd8nFv6siGgIQbEStidDuLp0ij1rU
GNwm3c/p/+xSeGw69wEjAP3uOYobxISoeNvH62VJU8QAUXZXsoP9Hh8ido/7Ls4C
ToPO8eQn9GJ2aExKeyvodHAHkt0TTWzsudqYZWXlf9FEsnClkdXwy2FMAoocb5lQ
GSrlvTcxtEYwcVT+5p8NTcpdZrjxpXptIrs0ed1ntU0k+ckdOp09Pw2z9AopPzN6
K6U7ITrt3DV2UioQzSvu47+uXSAVWGW+L/M1OwdVVGR7eccH4YpPZodummlQu6DN
hAAPrWXhNrW4o7oczf80haz/tU1HgmO6mLcUOtqyxN1xi96yzSKfsKTHnp3RW1ke
ZIlW5d/g6EfCnU00Z3Mar3nbSd40jADWSnixI0IPkdT9gwmSh5ncUUNDkOvrRZ7B
qEg5YgYvpZe7nH8+kKa3t9ohqhK/E9VzSQQVJH0H/s5LlDQ3RbuNiJPoLxiwx+z/
ZKYJeatH3Kl2aBEVnViU0PaDqu83fIudrIpehmKwJfKrs6IcCngikrloUZzVMSYt
bmLmNzApSxrkqLLr4cXUqe9vL2xFJn6VF1VR6Kc5/gZ1NcaO1y4mbIJja+a55rVk
qhz0ZiSLjTVFaVS8pnXbIrwrdGzEceJ2VIAQiB0TaMe8v036jkAOa03RlwRGMdGv
SUNBe6qIbQzC8ESYekikaSCMLxqYD6dLBsrfLA+uA750v0lyhk+2jciZKCOtqapl
h1FBpxsox7H0xJLQCtZiDkJj1/NjabG1QwhXpcCak65pk4lyhosQq7i7NmNm9epT
Ebn5DGgm7ZcC5crB4MPcmN2iCGtU6+kvUbCOvJXM9HrdETpa7a3D/BAMcIDsjM6J
c6VRLNFLZycw4tsBQ4qAEplHTMRBsBEPxKP6De1GrI0F5v02B1JGCU/FU1mEI6DE
wlxYL0NtAwTAk8AqmAQ+jo4Swy/MBQ8uecB8hzCHFLmK3HdsexGAXYEglmemY9Se
4OVzVImSPFKt6QcWE9NPuROL8mEuPDEhWiT8kopPOY6qUXiHFcefRpktunUB9O+Q
I6/rGvFbk8cZl3do9rd8ZeqWWF9g4Awm0wsAxgNwUo/2/WYlQHftbT5wgSRRhAb0
Xj80aPgSvqNQ2O3Vq06C3nfV2odsz6yFJqu4BwjQ50ivorl4+wC3Tt4NVYRUb0C0
McOQSRM9jilUzkcUP/iZfjnimKPJcVklRl+FWPpCWjyD2L4oD6fAuzIUYbDUhbR6
zcgZBC4doaY6F1aoTHPDmYNhEJEvRPiNVmMwVO/dxaI4lVO7swLqzkUZrtMUKU6Z
ttqbkJJJuOsAbL8OHDREkFB0vIWvb3mScYhu1f+ysK3X841QGYTtzF8b+ojPckMK
wCZuzhYioF1HK7whmG4xpV6yqQ88Yu32/jym6NZaiqhy+bCOTsvxmwZAFEec3k3a
8/m23aDtCFsLPgomyRl1c0967wG1IIhNWFmX2I3g7FaSzxbM7xUUZsNES7k9D/VV
fmLM2/MK4aFDFuscspylEtvQGSTOH7PkHF3PUAWOdK889e/sXhgWrrtum7GL4iaR
fXv4NPnHX2RsojEdJzoAo7qyHPXM+jZKa6CRu8B0Ds18++otrTf6OGglPnp+uhSl
6ovprK8YsV1/LoYvc8iPHAJzS38reMGWsCpWCGjJq2nHFgmr/bHZQ4KYyG3jUNnJ
TKHLGTTnOO/5E2f/KnN6pjo1G+mj06gqKIfuD38Zg347pJ7sYoM8t3xg6G+KzVzd
rsavxul+awgeWSV2YGYr78kO+am1/ANuo1R3T+lNG0qtn3vLvB2wKvn6heQkDcBH
AWORuIiCzEg9qeseAIb3p7ehFqUE14Ol8eekHVcjEKJhIEJc6TtY0vzIIZbijiEc
UY+hGeLGkNVaQFi1C8HHqVVUdYMH5L5axEdSycwg5/GvhBJlOKYW/hhWik8gEepk
CA4VdpoLBJq9P6x1iVFZw7yGmPJAQNU61pGBgRcMlyEb1CPMhBvAmLCtHbXYz8Ry
YUnGyvnlHjgzWq517s2lUpGov1M3q8P0jchlJ2hYLRttJla+kwST+4pBKxz/oDJC
IBRH84x4B9nOzgGYpx+0pAUzHo6UNagFV8VTw5GtThaK6kJpWv9cpCEDqKkngbOs
gelwo41PJ3cjhYECCyO9b0gMfpEowInjYcxQbrJqQbkmDpGbplujncNQBaUFFl98
zEAWOAfgFA/+Hvy7Vv1Ye6aBq1On7WaDTDCGN/VpKhKRga2a7sr545DfOqr10W5H
9yNTme40wNze31TcTaz1sjmBj9Dd5nnMh2dxWrZtGPMaFfhRQvr7CpGUGhN/4sIS
qOly1tgzREyGQxx7GLTaBvA92ApAIld1HzLULQZ57nqCN4OnQk5YGfilSkwYsHD3
jHdSUkrOcICQZZgoHtffySHPSYK37b2pgjkMUC7QojGAj3a6K5W14UMVIxVrz300
RA4yG4FNQpheO0JHVQ3vX+pNBIO0/2XrU3zWc+L04tC3u7ItqEakMDQejVo6TlrT
mK3v8xBm55TOInOYutx3t59009zwC8h5EJfq8VX10kRvbZo+eOjBOfHeea2zZm85
wLNZprqGfOMnmCDv8O0vEaqGVFwyUb+GvWR365xmEubsBzmHhp1ugCiO9NuR3G9C
r6GO/ENPtqMr3zpSbeSKG6LjtFBZ1KtJCiCDjHlls/XpbZ1nPmfhBUltNPRLmTcC
E0+3hMfDW0UzVdMOhr6AvvpVIrsP5XllBTpxKysUPO2i5g0/OvUCYhcy+dzC9dEw
1TmW22hgoyC24Yf9dVw4s0NxuaW6YuHpuSw+QX5N0RJiDj2A7705qTvYR1+8oKEg
DmjwBzx90sGjh6JQnWLhnBULfPGDtzyyGP0bjEB0M8BLNAfvHhBTKJsIjiJy1A8W
DYoOOesQCUK3AxuTPelqINzFSaSALOBxk8g8MnWuv8A96tu2ucUur1ob0VlNXw27
1VcPQBSxZ+6OahLb3m/NB/7xxVygbkHt0v1mS/DrdqHv6fxfjRsoFhYHtC7mJISv
x2uJrbnuCFz2ftrc9GBCR16MMrbbeXzqqYOOocY5kudaZdr6I+w0NhvWvbBuH9P6
Gs2+E5Z8qzieJioBP1UmNystFOu8W/bqJdeQQwx0Scm2dXLKutErFn+OzqNisQfx
fCVwsmxdDMxtM36xKvgilNjfrkoxyb3EWuROWvklN+bDuHmZfnZnWHu9reiJfj1q
Mfp+cPjw6DQH0f+XpSePLlolZA/U1dQvHFbOUlE0xo50EX5hbGHLzRwQaEg7iKtC
0O4pGPDJ+Ktfnzur5jMR4OOdkE0+XEPY1xs31/5bbiUO9IFAoy6n50irm7aF/y49
HaWBhukUp/bWK2YMzcfQ2N6vq7zG/9ZkW1HxdcIISZvCHlzWHIBkpEZiTfZRJbUT
hc0loSgKnFa6kbm1ZkXPG/uLhbGrgvSIlPl3l4uqRJ4sHyqFCodjgA/9cj0bfSay
JvLpW0+YtbIFFyMvxkZVDce3NvwkH7298rESf5/cWyejWTPhX517O0eCWYgdoFzB
bSouLE2NXE3qSLuhiWelhdVoxhAJfG0y9a7BKolam1oH6o+mbQTokPHqbnzCaTOH
9nlCQTFtcRFJ8fSpR1WuRronfveH5Jfl4mq5LxHgzeUj5BjWKVF7TR8F5zd3rQJ/
vo7ppeFqjuG40tgmtY/nAuJZ/U5UhKwDXUfPx5fzCIirzgjt/qIlSDTPX5xEhtxn
6Iz/KJusOkZcvMOORDIsJF5OTpXIsNRt9n6U7fgVLOV5biTFzxG0Zky7YhDTE8IU
2szz8dY94MBzFcwGkCH5zLlo7Ov6HJ7glzMIXarzr4y8iPQd5vFIph+9XHYP9bXF
F3unMv0wABDfDKI04g4/KesumX4BmxYyfWzXvid0avA/PnlmmY4I3kqoqufRgR2h
+Nc+z5tLB23igfTH0mniWUafWhzMJoc3pnGWMJuGJLkWFVsj0MViVBr3hZ14eSgn
M9DAx62MSj/4Q/zKXjfEjoJvApVmpFRfY/vc49rfLQNz/Ce+zHoa4eOpGeZQDq5F
hB3W33G4jPvnOgq+MUURRpfqVpiSDlfzT9TaCbXS9u8LGbOoTuTeyKZBoE1+cp3o
enmH26Yn+I5OLJJrn6dkczKX3dYBzfx0D4nln9FIrXlMNiwbpvN6VeX2iHsVKrH5
MPqoswn+rLISA2ZYBubiksQqWcgPN+ubm8oriVI5vjvJREY1/HQ29bKYKatUCi1K
hNcCxSSvhpeiBtiMQVNL2PHTdO4gwJqsKaJEGgajDhfIZayNcmJH2QyaoFginQWa
i8cvCrzI4xrLnYI9wVsDrr+FgROgA+vYO0HGJa4zmU6qwWjEI0nmqs2or1juRAke
/qoo//hJdofCbYZP6pqV/rDxshyPjJIFu4Xg1Zt+FnBIUGsRmd2+TbQbksKqVGeh
jNYDnf6OTYkwP2vDPB46V2ckfEQgR7XG9X0VQol//t5urIYeQvqFzaRgQN7P/ATc
kv6zgRH8R1HuIso8n4aeOzn7z7qnRLxtKnszMy/oJ3kqyNMpPpnLQsR1BYYndy41
Y5tnYnXsGw6zhkgHvsy+kpbDjvLkbxdsFU7GCqvyvjkr9dDfaJwocrawRXn0SL7L
ZYb0Re/yjxs1k62qrwShHGk6Nve2pmu9LMo/3Y0VJvpGhhZal2U9740IIg7FEdze
PeewUNgVZKTkghunWl2lzcMCkI7Fn6499TIKkROQeFH+r7ToLWx69hiz028P5D3G
HdjYo8qfk4PJtC2tXbsMYKgtBxgeAXrEtJE8Ejcjn1qRaqyll4HX4MhoJg3hEdf2
doUHcsmfyIz5ViLcq1w7ZMkGpBPX9m0grwybA6r95skqejak3lfY/GhXW/agLc1r
Ka1tOKiwjb49ExZXdsufKLWXu7t87zojlGvM2J6fW1s++k/7oR67E2lQv3jTTZ0j
4l5W68XqJET425Oa8vNJDUo6uDetP8qnHw8M5jYBwDyx6oupcPgu4+TMOEEgtCAo
ZTU7unX9KP/vHvrWUDMQl0rG058Txs2YnbEVIwSgSJl4JEA+wJSPeqYWXu0MqHj/
PLZWjt2LUvgP+KdTSJGDJruhatu5l3Es12HowWlyF8zE7cGP9vNuv3Gryp6JpEiG
ozCpMfG8M7kPQJJFuhA7K6qv0C/UeEDBeJo4vqURlEFEBlqeWAyBaXmmkNhMNpnz
VYaALjwhEQs9eStE4E2S+sCUX7AkmPYI0nVyC1AZF8ckV1w293uVP72GiapPPEnb
QlHM9tC1Bm2PVKdrvZKgwd+BzMNdB60U5j8NOJCfi6XeOJ78hCkOFosSjDVSZ8qJ
M9PkveAFNto7+zcvtnhcsoIXitdDqAM/zDlSnFf142ChKAyzmscqyXJ3nMdEDN3i
ZVHce8ldr5Wz6w+9j6R/55wJPb+IVRopReKbgIsAqQn/scePDI9rRv1gpHi01G5O
mqde1J0MTMTroiUXRGhZTY+o6sJRsGqu7O0324GIQMZiEn6IqU4TApwxq3fsj2l7
twopQFc1s4iFcahcGjuq8SEx8t2jSCORJiE+asZYsBluHaF0RSQMhvxag7EFVbiw
j4HyS08UEvvOmvPt0oEk5zHLiNPC91Md5REmKYrreETqcR3ZshPDJ29wvHocRA9N
GSjPFt/YYFngOuN9IZevBHpTRuxMXyH2tmUKI5pMZzmrwcO8FjmBgjI+MSSvcNo2
qiKHLif4/fofORj1YbTMRo+VC/z5ew7YKeGuia2m75F83d+T9Uf3P6k5mBwmFp1/
vPQTPeV1knYDZeIik8kqpFnqm6QtK/N8MWZCz4nYBBF3B+9ATGIgJPqbUbo3udmW
bkc6A7D4HnZZcL5ga5sQBrorIzWfjgpeRWR53MB5lKGfhDm1DdK26OnJ3k6GRopT
9sJX5aAUI2uKXngf+hC2LQBhzauu5uB1kve84nkF6AV4tYgFlMMRaHE9yeN4q2HR
rnk+mk0xkppqZd/v5VHxLuL8DxvoWgefa82ExrlqJaad43RTk22ou9tZtZBPeNmB
AT9DGg8N9uCBJ4TYGXMmxOVttLr1JkVA6baPrhzsbDaIRskyKs0Tb5bqXZ66g74t
Q8suODiZicBf2zGqbM2EIlmGd5nnqZEoNbv5GLZhbRsC32FkTrHpqIb2HEqOGHDy
pf7hEgV7kezBfBiFynx9doKH00rAt8LJOWoR5VP2kKbTlRtTUNHnRwansdjWH4Kx
ITcmwER1ofAD/GfEXq0k4Vr3BPOYChVDnICWAaocvLHN+4lAE6hIYd1IVco4qEcn
V+fZ4rD4tagruzw5SCPJMwovL7jIxGTKcGQGJpxGBPKlDrE0/3eEO6h+OHCudRjn
4QZriRwet0l5+Xm7N4i1bEJ/qEwIm16ne57gfuTrPfqQ/krllzyfK9Uv9vqjC4/E
iQaro7dujopNAe8oBNLX0zslD4cQ2dCSnJ1G6Q0njYFBVE85vOKHXYECpjni+WA0
09nNIBwvvjgpxsNpnVTRfcEIBQkKPAAGRCiIVuMkx3os6gJq8yQzI6cA0p9vm7M/
HBu8RKhIYlu0/X+LQgGNmTB6Tk/UFHVx1Au+ODMyFY+xRT4w20b2zRDprd/tJYID
k0UCEXoKciODoYOz+NDp2ejw/6dDWBdGs+cMJ4wTeifDf9NPl/oXs4tRLJgLkb2I
quV+L2hiCUxvUTgOO4/3c/QzJ4Zfog0NzVwg21M+EcGz2K0KlosavAM4xoWvzWnl
AWPrOUVW/6LfcrSI6xk74hp8y3IEOK4a8I/UIHc0U/2rF7KXi8CanPojrMsu8FEo
vAFaXe7pBoBkPwHAqSBctH1AhPuFFQCrOH4I51aVrl8iPaa3U9iUtL1GcJaHEWjF
FksUlGQGV3TyloYFnjrLW7qBB3Ptn8vnw/zePFzanGx8uRmOKPsbFrEls1iUcBBL
IaF+pR4GsmuZ/f7hCnanvnOIzv0Q87X0TjLLtyb/a5fKPHNsVFMDrQ4Knwk58lG5
1gzvp++p1PETagqKr+AHgPJi9w1necu57xz9YqkZmwV5kENwR3g5M/XEvUdtjoMN
C0Lbmv6m0SvhhQK7N4fd+zvXg+yowG8EDnzmUAEE9wb4Wfi4M4kMxOUg9WAeD1Y8
1vBH0OhmJETD2y42CR2pPxXHe6OeLqElx0T/CRihxVKVuST6DH0+E0aD0cw2Et6l
mlWaDytwH+SP5R4IWZWhjifWQuYf26XB7ZzgP7PTooO/45Su/cMoDYx70ZWE4WWh
3tzF+NjX6irC7ET5mH4maYeGVSARcav39x2J4CiIpVBEQGKWQ5UjYYkNBPBIdWgc
m2dagBb+1+PFXPsXWQ3buVbJrOuFvlqVDxQDnQuoU5X+Dia9AsTkDaASwjVcEPWe
uIbMQbGCwY7pqDoeomhw01p2cZMDETu8o1X3Ud4BhQB5gSGHy/WTky1Dc88TXjfx
SIdb5jb+lHjU7G+Sfp/N35Sht1hb68exU01hb9G9as59/0d3xjSO72hRl/atSPqc
ZKuK9wL1A1/xkRBh13UBbpA9sHxH+QwygIpRLOgwn72jGKjqxLCrnUcUBuuHtDmQ
5EWhw04b4OZ2L1kg/kt36wlVSJUhq+YvuQCGCOTfHq2kU4MSPR6NKnAzWPlapcDF
WD2TKC/gvB2zsFvACFVfnwoxrp7wOCVdWRnnj5qVGg3Qri6X2ZTNRBQdqvDIDKlk
NISxCCimhXUOVkQhpRKRkITL7/vO8Vl1uOKguC+pYf2Z9NWTTA0a9hJle4WzAww1
q3hxlZrebkgqCaE9vBlKmzINlw5XG1msU0SzmciEGDe+7W7RkPRXki8aonDI2zYr
vpWKomIRjUEhdAsx7fKBZPizRd6RmVec8AS5xlJAZZZ9/Wj/3RLbvVigzvSmsjim
MXxmIawpFYyfsgh2NsxjlLALweOGY/eJ53S+g07btGrWmdChkY0DG9kj8Wky0FMU
NNLtmfwW9ExtFU+gGYkuYg/YWAz+hj6Qp0wSzQjc251cIGCkpTNItHIDT2dUT9nn
wbF5em7aOX0lFlGJVLnglqS8sUgalPwROG9p7yrSM8L2kwBD+ji48MboRWFyf+Wz
p7dxw7Kj0mx3UhzT3pZyB/N8jqVuiwq9j/gyT4UgSaBMsVd06jjtJEkpEMraZpf4
K2I4CSXpJ01xkYJthXY6+wupoir1RR6F3RbTtDmkjk23/ViTaWjFBU//g1tfxyID
x7Fef0PjQzOPKzDNkUWMz+bT+pQJfiygD+qGUBcTqizxW70622I+dPacsry+C4Wd
xLU5IpQjkUJdJODHtKtiw9g3eCtOEw5c0R0YoT/U2jU1MM5CRfcEAY1Gv7Afyaf+
rIZJiqX2D3NYFvAT+AIVoCO8mdMuBgj9I+iIKiO2HTayMF5nRfo5r/JRAWJEUsFl
PZoZQui47LjcHv/MHK8oq2hcYGT/23D3j25BAjCS+KeUTNUtbp5xloOcrfEGVC1i
XQOGn4s1uwa6i0LkKSSU+6HuYRRutPLTX34CMUSjYLIVbB4q6NvCd3s0hWavhz9z
oh79P8/cCd9ho0u1rSHxC0VPImNJQEgiP+o4YHWbVcbKcP42FNAEjOE+VB58IuNn
yqJVlbzKmLQSjWyak/gKqOdFmzaUhteZzhkgADg6f7FzdXVKKKBViGDvsZw53hQd
lG6YKsbzBzfNz4ByNZ29lYphHRXToDGPyOKSE7jC5cu9X7Jb7m05PEVy0NFfUD+P
klgRBlQYu145eAnHDVwZdygnTSBS/0nKK25XxJVZxdYcms8+xXMcvyHvg/pgXmRs
1Xk5AM6ovn4bYdpfKAphtIpTuNvu9q/qIUifqgibwfbwcZOo7fWlxf5+cVv9HkZD
IhvUR78z/TtCDE987gGjfYyCmTTz59p9A3y3RZDELD9gQt8A+iwCa5A7kIYMyKXs
SGpNTmHfNx2yMaXSR+hkHyasvp49TL23+Qrv0zLRBWVv2csyBiQIeJYR1dS6uafk
6OLJn7EqW7KX6k/umlvYCh9S3hQZ3eakfZy5tbC2VgeLyxf17YUBBcNfSiQygSQR
0PE6OzVFF/KOOXIH5ra/xbISRewHNIKEgC2Mau9I8usnXqOqUbb/R9qacVgLeWAQ
051ORMdqW/wuPwHxlPL9/NXehP7g+RBeUuhS9gifFE9+Rx3MCLkVZ0SVF5U3S1v6
+aqpWztt9/+Zaqd7/5/w27VEzKWWFuKt8xRi5T+npdbT1moHfIHcq0Q/oMKy/3MP
21OPtO9S5fDWyVqxn2cBpQ43Ty+XCyyU82oskH/j0lj1vD32mpsEvQ6jEdH6TmVQ
VmFDCpUN4N171StiSlN8HJpYpwuybLTJ35bhGjA+1ByczzuuNQ8pAHueVvX61moT
YUuHQMuOJ6lb27FVyhiFNdijaNUdeDoucWC1JFm85A/75FFd+PJrss6bUIXaGVFq
RiCgZomTf0+d8W5WMTwBaq6uTTvc/W2WGb2Xvx0Kpe6ggtYhDw2fP3n0eYek3vim
KoE309M8F5vATiz2VaAvsBVEJMtKm1BKJP4QVUJA+WGRgKcsQsBu6zDcBR5DowK3
y4cY8OkFftu8XS+T30IrDW3eL0Fr/KR6Rrc6s+uhUK3ocBnK+NTyUAogPY14YnrC
OaxYjL+VAev76p1tMVGTo+UTtCnGWNc7gtuBY04ll64zVVWJaELLXRU4q3p5NJyr
keDwEfMgKGZ+8AL8J6y8yDKPPwPWJGy+LYltpm9k64tBNQAw0uQz4Cw56/Vg1Uri
Y15APqT3lKz5/APuChwbYQ1D9JrzEM50JIDI3ZN+13DZT27IRjP/lOHHbQug3E2g
MvSugenqOY7qOe5x/pZJZNTD2HhxMZdafgosHOuqlSPuHOVVPM8UxAOG9XmlqnIp
j3JsscW9rF0zpkWP8kVu2wYNWEe6d6SgjXEZy0YhmYoa0Ivk3uKjMA3VX3lFY2qH
YeE/om41IkTwWWi8Y67QWF+jRFmZGyGWWzLOrfUd0rGirAeOh4LLEtW/oCk5Vn7B
/zINu9k2BzeFAEtEC0jSYeae4vKtRCFz7lpfzgOQEWmg4mdAtGXPO4hLfa90e9D5
ZZGGPkj3c2D3xnTmIGvakOegiFu9TiwglY+hrtjQt8LJZHBONhflLpoKy73r5sVy
Eca2m3tbswmXCvG0xEdXmQdjuIsgG/pkuDVKOIenq+W4qndDUoRVJdRInrgSw8z+
eDBk4EvX7+GvCFkmFwFDqVPoBtzmU4blYaIbG0yp94lR8JWjLMW2l1JZnNtJpWKM
CWZ9foZs4oLUalWGXMz1Vp5ECsnBnHhDOERb+3KX0NxkwHe4dtFyRUFEMGwOFGzs
QBtLXoZc9DQEvluxvsX5vH48DbTgVxFtIa+9NDrnjow5veMI02gi0sVAmfYqc9gr
Xzi6jCZKCIHFvl7SImhrK9IPS+sSeJZtjaD9h3KY19kE3GRZWF1V1czKjucE6fr5
zPl30zvHyWzOdrXNnNDum6PrAhe0icdLd7O+LwnKRk9lzusp8iVx9ALJGQeYK2Es
GWRGuGp0j/vSrnXl8MwqZr3wGCCSRvYfFkecn/lk8M0WIjXzqEe0KOFebEyAEhdC
lRJCVFpQpa7aLaQipSrqcctJT0nuWYOa+BA1Pk+iXF0BNn1po39v/Me4zmXBO5Xe
o5FO9pTRnq/KpqxcaHjsoFrvlJ1JYcUTWxJ0URcw0jTNSNEFTnDWLg/s6YVRMEaF
IZv8QYYZSxCj9jMr3YcGWg9+pZ5pMCsTiSGB/1v8yle2irYTnMVB4ZFkMLhOZBs7
zxnUVMV48/cug6A3ElKFsFSmLNO2zDeglC2qk3lp6prh7qdc4GUicCe7NXiTP8Cm
hvvglKAZIcLr3OObNJZCo6qnIG0dl4Xaz+bUk3+j7X111+8/nkl4QuMobOyBoAP7
3DxHvZqd7FmFk+ubBz4DvHUBXSPGoNt2HTXxu6q32aHPo3gIt9HSqGZslWURn2fq
yDWiVKLYv0Lt8Up5dxoezj9wGbgljkiq9zL/mPpyUeo+92a3GjK/K+/IwbkKWb5I
IL49szSGu6Ou92ER7EXZ/72MstbtNlfUuHr3AmcGO0O2rxfMLKwQugxBuMyjzlG8
WeDn4eW6vD/k8aAezYaqGaKeNW1k3Oan10XeBQeCN4c3My42XGTeziJL2yC3NrGt
iuC1WWnjnxD1I9+4WCJ5cM0RmfuJ06w3imB3wVtWqR165iylP6K2UBL4nsXfjp4+
rFO0USyuATjtZexWYuBb9MlUqhTCdj3JpCmltSVqu76T4h4IN7XhR9ZFXRo1IsTk
n91QLy2twNjCoepEHkiBjjQNa0w2XMK8MHJkDcwg4tRgLPZSbOtdcmt8criLvc7o
wvbwVau3TIoeUxtC085KTplfBUPD4SV0pf5Y5te21DdK9SV/CyasgW6xfJbYWK1p
OcfjBt6Sl+BVyYt/04LSH04hSz9QGpjI+s83Y3pt9uU/mwD5ha4laJZWDovGhxX4
xYsMLZorPTY09MWFBD5ro9Kr7TqNihOi9yAaxpnlsDibSaPUv9i9oyYbcWNX9VG/
Vn0mlxQ0ZRX77xoGBCfsxIWP4ELL52PKsMiRSy4iu8+btx/ODI+2DEnluXEOxnmG
kswMpptFJS8LhQBBgJ/ShZ0JOVoVzq7EU65ZMU8R1N6LO7Ngl6knmhRiDCz4GWQP
KXNxjHlV8FU0GDd2RFq8bFPJr6h64sg3lsAUynQEXx9bQ2YhykxBpca0asXLI7SU
vIxTgORtUCoFPdzHn0xIFrd4fQXCyD1jZK9A3ULeUK1MIFCmUnV878lz8CxNLNVP
z4VOtIV+tl+hXvuNvVk3qpyAQGyHSxKI5ZErIOf2T2i4Rvg1ZwW46wvI2edda6E/
Jb2SisJWVkJwQBm2z8ewkE9tyezV4F6AeSCQ0IcANvoyc1qvgJXIZcpAzpu3PgR5
gg1OutT8fwf3kKr+bb9fXbFD8z7RUsujYbZzm5hFI/OaId8CrTMJZpmLPjBf1PiA
i0PI6zSm87teXPpOuzOmtFWiJelxf8T9gXBtz2gOpxMKB9sTzNYTI3FRtww0QQd3
uQ7jCDs4H7t/Kw61CerT2BxjXWK6Ss50grJ6FJt8Yv+cylYhhe/J+B+8g1n4iaIF
sf3vKLudM3d3RRrotPEUM2U4EqdqWL8bD9OCpYI8VPHpy6cswra72FZy0HL5yVBf
7B0p9CumQHZZbBVTjPUKaAY8o1DDQuxEXx5UX3Ixhwtr221BT7DR511BFxHeZN9t
ShoTumPyH5WNEOBgTNMLe45Vb4ljm8/UlLeED1BLIwel/y4DkGYho7RSyh+Pad0Z
bjw2P8pUtJ0pB7a5j7BI6FekmFTGzitufcmoHm8eHo6yfY00XYnOpA258QQFxB8Q
1A+TzKXgP0+LxFCD6zXYBHAk2MNq1ALSOaxuwGXS8Jc/AwDkiMRhDnMiBpvTjFqR
CAosfxpCRUJEfDnf8fckcoEl1w1LyLV7bYVkdT3xXbG07vyVrfKxvWeAA/UW2syV
fDYwHW6UnLBCDNsRCnL37/vRegMupe/O1wsYNzL+I0+H8jac19Ze8xo4imcd3yQU
eLIo/z3gC5EMAKvlkc8f/x1oVCFfW4xjtM3xua3JqskIOCca8r9BD9Bezoh9r5Do
326UhOsFLcMId0PhLjPQH4ubrLX2qsbuvJXfaU/66QXBTKCHmAaJwG4UbU9NDbri
LjoVRSqZB89prKOaPeVaInPlH5iSiOLJyU82iAfSHU7NQhyRrODbh1fxcLiiW3+o
Vm5fH4mwQDCawyhuV53Nh44m8Piy4UthJMrVvG/69w1cAmHqmcZr3xoK/XEo5DjS
M7Z8OU700aClL/8Z5bL78WDz3RtWE88ckb4cLCtCv5WyHcVM5pALqdP2jOSR+1Sa
WAkK7O+Srzf+ckLLLVRM/SlR039gSMzmvrZIubqg7eIYnHfEwHENt2PX8FvGPNPm
5XIwzoMmfax09zZbDqvDU4n4y8OCxfxnkGPKNtlVnZ8kusNJzJ/NwlEpGNj9NOIy
1XhlGmq31MFDfxUXWv4q8QyvSOFYK/a6sLhxLsd6X5QahcaQ1QOsYXL3JdBCqm8O
EIuuWQDWkTNZrIPPedaTRPgzydliNyt+8j9rRzrzU3MEkeuU8pSZVDO3Es6PwMge
ot4H+TCczaAwQ7JAQ7JFShxgxWH3fxBJua9+Lf54qRuhsdbjIasB0Jbrjga82PPM
CULYTeZOBFkCB0kTCUm7QkD6Lw7/4idp0/ZvFGq5AkATWNGF1GDPvAmav6vY98yD
IMC157J/FEbDj1NpyTtcN+gC4AnWLyQtYB0Tp1ukzfxA9XS95CZl0WkOWai9nxMU
1NOltqBfzVBQwm3qCsvMo3f9cvcyoPchP0k7KMMue8aEusXk5iO9Mj5JpWyXXY63
VUeJiUW9NYBTeBJYO+NDZn2uImU3xPNVn6dwEPtTFnkG8HmUa/Ab8drtZPfzQXee
s/WLc1GokLSEE3AriSRvvA+WrLlUX/gbptOL/r7EdJVqXKhsMKU/mjl7Cd1lBYAe
PBw4OOwruwSqVcuosOrw6v05acYLU03oqvE9IdZPrd+r8UudA3REIl1Ldr/CFV6m
5ylYzFYqHDGSH/m6OASnFYNPg70f9PpoRErns+7uNy8vvH4x0ZxnjrZuvMku/WLs
8icpTzu2Nbvv0vCOVNKIPYhNxuyI6NK6EFkhsGBzoKcCY3L3OW75lmyNamThJGRw
g1zm3TB7novQJK4QgyJjFj236MVrcAWEhKF9NWOAVZzoqRc/oNetK27a3KPfqvEB
YV3/6/mCPQzZuQ+a9YhJnCotwQyU+FWAtKAsSCyY8AKkNniBWu9Imn52PdDFYMH3
pLS7FMriHRgDMXV8AbGq5awQqUCFWtmHsoJeckgjTVjH96mNP1j70iUrA40KO1xk
cZyfgk1SM3PeljJ5EP7mxA2bFtAGRjCJRB99ZN+PMjhWPgnxjYMCRXRog8SqnoQa
LTDUte+u7TltjMVJ/3klfjj9X9AcGyUHw/LpsuxzhjhUU+dkogAC03+Ef/6SS0dH
jqvsgFzltYlpZyWDxHV8qwtPfpaLCLzGpkAXKIZJtC9679p7Nqj0zUhmePRw7CQ3
e5d0XZjzcQjbrqNUQ38N30i2ORhXt5aY/2890u0Wivp5/UWzto2cGKWDMzb60pdu
4CdXReDZOaKFqZTVIh52fjHAk2SjYBE4/zBjIbb7r5A2EenbbXvdeN70cAE3INZ5
i780cPZD83q5NgYUK0taL9f4X7lp9DlAUVmHOvpyUMJGQV9QUvmCLMg8wvYF6uuq
8G27ScJSlweAuoYuLFJZ3Ajiz330cJy8AwFnOHxCHHITlU+Ql8LtqZUwHP1gxxkO
U/gnpS4gM7mAO9urdh4uA8KoT0hxhYE2c3ZoxfGn1cUpDMABjfsRb5dT3CMl8Ace
KCKU+o0qKVmzTkEUkKA/LbIn6eqMtgm3EAuxYeOC6ZKqTWpGJFj3wwBDJ+NQS3An
pejzd9wCoy7/cRN0qdJwWlon+557zJ21jWWnWPSysVlJLW4WA3GqqEfUifVFiZQD
LnomofHdaLIn/S4OaGqrnMdUIZNYIwGTxp5nITdR70OvQ3I8JpvhvbRH/Ed2FUnj
wRStQCdmXIdSKQNT2dIgbaiJOs0wQWMZPNKQyh7IpFycdsNbOutqyGkdxzFTVYUl
7kJ/38YrP19dct4u29/jr60Ay5CIhHOPrG+3KsvD4u1UeJ0uow9yKHba7mJQLv9u
T5ouFymqAwVTfuyoBTfsm0WeQuv56/EbG3zGpXpOOLcYZI2DS7kRz+dllEz9uJXD
sRdOMW8MoYSbPlJHRzLITgqmW0xf4v/nb3UA0m3RB4fsAlchtAhw0S7La8mUybob
Df0+yBo3eTXuqn1oC066JevdiRsKFFTZJ0uj1wcPEAkNOptKrAXsfFkFJcyvWnI8
62i3XaouwvkoNvlEX9lv7/19/ITS8LbKTp0+uT7PbKzdg4S8i+QV7LpzvC55swj5
OrVN+QhbY9jAN6ubIAfsPjcpAuy0Z09fIOsz7lLwOcEwXf0c/pE1H+p58xR+yiI7
/lpt2tjBiWRaHuf8AwYZ+7L8h2ZeZDZLgWK9SqZa5txFI8ZblBkmevBwo/Fsoy6V
4xzzmr1x7wVjm16TQTmiY/Fu9OO/i34m19UUa8nrEjn7sOk5KJNpT7rjFlT3eJX6
JVX5P4f5dIUPU8VUmZmJShrpgKU6iYe6sagw1UdIlHXgwwJWaq8fXBE1LL/+2QCX
3sjCpCyyw7PgzLZyg2TaBDfz3Mya8OsSJcfDzWNTL7OBpEWgAbTiaabM09VrkFLY
VYll+Eag+6XowSFNn6+COArXrQp58YvAAkALJv+uQXqU/NKqOYWMCekWPkIvUQ7x
v9tbLm2e+IZUV4cT/TuPzkOdiF9TNbLNsOqtV/giC4Y99wzMipH3ylVnbubqQpuZ
hAjjmF9Xas97atgQGooa7fe+dIG+CyX0m/Vyc8kkkmSvUTkWGk9U6MgHJFqdE/0c
EF6up5aGUr5Ob9DSuiPVg6+duQI3UEl+IGc3I/P4U0pxSPhZ3gdYogNkafFUQrfX
ohXOq6MlWL+sdMFdiHbBbVor0ovbfpcmAGoRfEAs3hn3R8oznnheSKl0t6+Gmzav
kEwqIr5hUjWIqovhOv0rOT+AA3noV0NYxBsrtyu3qBQNxGh4QSHXgCF46f5vMBSw
z4I1TyQm3wGCm9/cOxZHTyFXpbG7tctpv9LIFC34uwMDF0bARDBP+Z8CQKgkReqv
yLWEEXQH6oIwhQoZ2HKkGUcb7uAfyD/tiYhI3izLp/GOv4Ng34cLbjk4S8bDeVAC
rBUgMWBpMgbZ+SB9W2LzUlF+nsaecAAQTEG7oXqXJWr09kAewY93MJJ9VKmEK8Bt
7pu31bqwk9subBxZEYKwNm+fnsKivD4r54wg6kvXaRLBLCEYghBO1qg7mSF4vvU2
TKbq2poiDP6W6FFjRZKUPhddtravnqym9XXZEw8aauxNec3BYyGrjfGR116ksp0+
UfAOeQ7ITkBmCJSI/XsEwur48exUguWcPdM6g16Q0Joawyr0D5PONirX2MEpLEkS
IOoB+7rWVjCqn5e8+vUj2UdMoafiith+XW35+aUGlhRmAXAYzu3aVM1xeLdgoFpZ
3VSYmgLHP6VgScm8qTWrh+YynTkLAGtmF9iC8WKK6OLWuvstkTRwJKz4E/fuAGKl
noILDqgrYHWYqZx/H1fKzfstZWiFauhDuu8nTCHpWtpiy/SILQY5H03fKfWwI7wV
qHWARgHlYo33WBlYFRxj9ElFzUA+mc+nTsvwbjwcSQxQC3ex0W2dRV1dUzCGnx4p
lUcteg8XU9aPJYV/XhKeuHaU3gQEqsXa2tgw+Wxhi2SHQ6ClQrx0A9oLY3J7nxcY
Dd4WqmMBPOSt+S953rBPWUocCByOHeFGa6oScmRmMVKcZ399yQ7L7pSrLo3+xJ8E
nS40+4zEoUG1ccwSuljXtspzgI7uvy5Q70Ths3EwJqqGxbXh0/gmpVehHK8lT8TR
dmjWz2F8pdWHTvtRIXqEXU9etpUMHqJQ4BMzqSeRBrJBTWKkeOgOM3xVRL5vkXia
NQeE4Rj+vTCFChB9v8SkknCXERAhAS+di/I0UKZW7ILSDVRjvmBUpmbCVLBCLGHI
qjgnmfPO3Rsz/RYhrk2sAq5SeQpSMmz68qNuDjbPhqgjHMajClNsNk3YVHKk8v/x
C5Bz0KGLdq0l2gFVFe+GNdTWEDsPjhbg9e5a1OIa+CSxFZpyVk9UH621h9HMSg1x
+A1PvI8eao6lUo0kXmYwS6BUl3Aq2B6kiM/rHGHjVHQDA9S4uZu07EYXk5wltoDe
1SO3UOV7JFBGZhVmEN44Lk4AAoZ88NOAqskthyAgUZ609F4/emvzEa3U2HkKVHV8
cwXHaLm+g1NmE1AnckOf2tGcp64Br4Ez0afzZwsx/52EqYcX7mp49FnsS/AKMQ6O
t8N2JqvZ1P1Lqr3SbaovkYrk7WS6QAzUwbI+qywhCy5t+BR5CeM+OJ9b50NlpAft
v0azyek3gGNWmSa5SE6c8XtLwk79lOr8T+BLw5wb3R0S7j/dU8+T++Sp4vhceKFg
bUTnQCC/BMUrMHcUnehcMOnzB2TlFrg5Dt442GkRWXLPGSBy2CkzvhfHjzxV/YZM
c+hI1qbQrwjauy+wMLlU+Zhj9iP4ktcDIKAxY5G9imTTMu2Y6Nd0hlMCPPuGHKZl
STthhV7FDjlGAf1b785rZ3cLztJ+npS0EJ9Zg01w/yebF6FbsC8y04kbtfWYdLNu
k8BQI6YYl+91yxosMBOaXuLb2E0quyt8h4rH09XkiuHn6M6i/nXJbipgZxqm4KYz
3pTq0cEUwI4xr4F7gySFRZ7guGNbHBk1K812nAL9g3pQfLZfKWDK3kwL2U+wdS+p
mvkLLPmgGVuQdOdBhYU85UOfnESGP2pYuRek89vSS8VZs4VYPUcqk1zGSU84sQqM
br2n2O5LktTHKLNSXIiQJ65E6jAlEqsWPtbg0UkVsre3ddKL3Z1OHvAUYgIYBC5J
0tD5d0hxW+Drr6Lu+Xv0gUU7HUiITV32+jd/FO/FR6JMxSwg/GD9G/dICN0JMYWo
Pu5zkhuX5yutJaQiDNa8zImu6rIcf3asHeTjXu6zSMMsO+2D/Wymh1wWXd7pfWa6
lH3JyjA+wgecZIQJtbjVmaqEOHCC/OUemwhTpjWBKVtZn1RONa0zN1V2tO3NwshJ
lYrYihE5oOaNTI75iwc+UbBrtvUXyH24fh+ngU2E/wDzu22WbkY6UPIYJeqCSH/F
9EwVCK8/uBdn004g6m8cktNFhDlZtWiPCrUUKQqUthb+eaAHIK8J1dWqJ6ioIlLf
1X+AG5R9nn34hf+02mNUAjaoDxfwTDTdVg2nKRY1VfWO87RzYdIgBkmlDbvxpzZL
jBcImrMQPTXp7yqlaZzcNxWerTLw+43oBhhrLA8ndHRGTG2wSkQj/axHGF1m3INB
90Em2/hkBI8ud8vSJ24U2+JYcFTBxYJaWliGPGbz2rBYSx+9tk8ftSJuCLzdigOU
fNPjKKu8EzrAOtNRW1eo/g7+zevHYNnsHMseum+f2zW9XjysKnzNf3Z467lXmbqr
WkPORxrSv3qe6bVco2SWj3uuYRFOWS0SNY27Xe70rYDI2n/Gs8vuk6Rsk7hONiAA
Bw0i7TfGy9xHAlRCdd0yFv9hJ5c7etPxKKr2ZQBwaGfhsE997RK/EwaVjK5uxHXh
zw/qa/QYUuZxSSTADW0S2jNs8qrVs16gxJRX0SkSsvjRo/h1fIKIvBLLdvRWlBh8
mACuHLogieap/eyu1xOH5tW/J986mUwIzBVVZkDh7Fi1kGHxueNGSUULmtBWk2E+
zJ0OFAfheooMbwezlb3XJGT5LiryTAzlxuNspl0yoa+6LrxC7aoSQ1n4ZPCX82j6
IdGVJCHRxxYCNMUid93Euj6st0gknQbFh2rg3Vq0qTtNoAi0gJ0jJyzD2KHxl3Hi
SXCG+3pmg+IRtlr9AJc8vR3g7R9xD9Fkt5eRWWcWHitGLjdSg0yr9MXwHTO7lwP3
7ieW1gWR8PjP1aGpM/0VI5iMwvLtslZnl25XV8HBzU3VtPyfN3LLg4dqfb7EnRHF
Yt2rVNzYKzUgSGJvFXCktRnIwOdN5KJaxaW9dz99CHoljhlN9CwTBbWoxpDSUb3F
OlY3jE8xYBqubtLriKzJEogfEwUpq6mcxy9Eph44ottl28T3f/dineUQrqvfPhC+
Z8y/mOJg2F532PCN8GxulQ07wGkpozpYYtjr24aVZ5bRywuxqfRwUAFYqknuwpCA
0FTLF0o8Pgd+P961UaEPyHs6wYBnazySbhfQYSy5Hb8uEwato3E/8FXbac26z6Zp
Vp/ti5ijoKmvQ6P6E37vPvO1vIfvLPxk/w6MgvMRN2TSdwR3uVDQUR2Aw9Wy07Vt
gm8xlFHCSJeJ+8JlxsuCqZEqDQf2hEIFvhzBOl1FBlmf8xEXOmWOuFY3xDkVpjek
hiFjQbkoCnRPdRGLPlk4K5dggDZbrpyBo1tYtWpoVN+PXlTINMycztAFnWj5S/+I
4yaBawxruplI5qnkYb2piDk6tqSUk085edm9U9uzw23MlEzvqjQk6PLl6SOoGkXc
MCGNN2rx6u1wZDq8ZJxKzatQwQDW4PkxN5ROPj9xp0cUgUzswlHzjLK2X/4Z+UqW
ISa0uWu4qJ+3wAWZLnnQHUxGqRYOB5QLLx9UOQGHIaUb/OoUGE8OFySWZkRbpyzP
bdq6Nf9IgQ+nGJKBdxoBxKBTXrN9Eg3J/B2IiqDX6UjI5HFXCQGJrwh+TjNJ7gFU
Mbxvp99q8sAF7C5mIg81zgB7CEcUJbuJAyVENdJfTy9+Ud4NtrXIrsdb/RgNd9h7
lxro9UhqJA2cfnFQtSatWv21kRaz2S5ggfcozHBIJQctaCDBwwXrhz0AwQsIqYHR
qIIHVMzX5w+MWu8RO0dwJJGUDPz4qz7w3jqYGxGTR5aejBtSwAXBq0ZAEUQD9mO6
SaKpPoihGMty2h2wFXzaoeJktk6g7VNJAmEzyA5R5S5NtOHcb+MYpfEn8gcWb8ML
tTGdZtZSjjFUvo32kPBI4H5dpzjMHjhQ77IcBhzxpd/WFph+Pmv81ENCDdTCZq2f
LCYMRuP8K8y79SA/6ArvN3DlPWWa3XVM6eSNMqltd2PrsIA+4eWB7HbnkxpUy3Vu
vN9Txd21uMug31LJJmEU2W+j8W4pz2R9c8tiBkTuDZM+Q/ke4WZpS7+VtTYoHTkI
PwMjOiHY1dZcRy7v2Dbb2ZGa+hJQ+8Wbj8FTR27PTtflUhhEFMZzKrfUWeIVBD2z
JH3hAgS1aluTYO0SZytalZwAgxL8cAdfX0mBUuV7tLRm7uw6EOkZhL8IRgGoY/DI
2/Gjm3oO6UkwVnivOrs4OpX2xEwGgVDF3xbaNueNds92qCwD+YH9y4b7qCv7wUz/
4KD5Qq+sBrOl12UeSeCDfaDKujYTAuRXgCk2zn0pUY2ifgEEEvVGGf34V5kHtGH5
D/yLOPX3AFx4yxmUPNPyk0cUOHrGb0F0QrrWop9FogkWUleqGJ5mypz6pJypOuGB
ACBmdiAQwBhVKdYbgjQCLmf8Wfq3BXS7z8umu6VhwbopY8XisyVqkFuuo1vwSX10
dk/FNu+Gh2ulmD6D64jeKCohrtbPjpbzVRViKeicsV+lPJSUffpikRAfQVwF+PUf
varTbC0bnA+VV985TIrZtC/IVPHnm9Jk5fUbQjWu75eqnwbjTDsM28S9mDSpSrYg
ymLYbYL00DNgBzL4pdhsZ6X8+XggZj6t5WTXPTIhQCfNr4TLz/NC3/ZUEmZJkB/f
QsPFy+LtGgK0TIxcYS48gX6yfNDWbgeo9v+mmI+YbIavTVhDbxaGDvAeTWDqiz0H
Ydcs9oRMfkChS/di4AHH66SvHav8OdxfYdF5/k1VhcAOfC1VeupzsshMwqrw9rx9
16C4d7UBrSzBM1k/sP9BV97OGym5Q9GJa6q4x9I5QO60fNTDZGBKJG8+gzUk5lGi
yK2OLwWjMe/+C1XFXenVKekSsshlTY/wjhStYWt4KQsgwcO7NpZ0wUKEcP038oqg
ppaCg5+BUtOHa6PLDL04V616IKP3a35m7XdX8gUvQyIAjQoSoifk18ZPzv2jQVE0
sZ6c/jnuurfbyV5HSU6qB8sw3Q1iSTCC89NIO4TPoHQCCELV26aYL2ikaTTNo98X
CW2JiI6kEobsYZ+puUYUGKplU/Lc3lgtF/NLQyK7aV/0Zh07uH/7mu4d0x3e8Xj4
ao7l407Wkcs2wK/5rlX0ln/BkcbWbe1M8TfhaeFnZA4tG5JhPIRbq7ZJPlqTnPDI
HO/oZV5+bj++L90hxTdzdpIrcP6jBPseT7kSqMMRkJwFIHLOofVh6G7D4XJmpDWr
uWKad0YFBq5PdqGn3ug9n1/HLpw9rvmdKgZtyC/z+1AWB0CIxKpXClqnRZ24IkyM
LIERT7nfESV/LoFrqaDKPX0qJYYOgPHC+OuF3SbM2ibqcJWy25GDtDjdVs2L8zte
jiuZUI6+tov1gqi+exoj5l/YoSUU9UXtsoA+o42g/Ux/Wp5XGXEvcjs2z1wMV+0b
2iSnABoc3FefE5Gcs1LkvTfkrj280MLiO/IP7o40pq35B05+Ja/zz5wuH5VgYOuB
CiWwNy3CkVJJ6e1LDkbnbtf3UzYDV7OsRwbP+Cd9YMGHDlrIm50E2r8B0cVvBbK/
jChhbBag/93aeyWOmq78GGHdYlyuJp6ivyXg12eJgADBwNx1D6TjvX5YSoUb5wPT
wuQNg8tCAgPVSOuJbXoD1Qn5e5EcyqgiaSB9btBbPzeNyAYOrU9JE4cdj0pVS9AW
RpG91nVSqvnXqhvRb0gSJ4WC39WsZZx/9ZBw++1mGijZ2VVUx2RR/yB4UTzdPOa5
Up/93UnKe4mp7+wM1S0seMAZ4/hABr/vM+O6gQejtgeN5vR6LutMj8UbOa/Z722G
BqVo4izi69npuZbKgyTrKy7qfZt4rOvw01d6KM46KskN1VZ93g0t+YY8R0d0OUdL
MsInPYsupSR91bwB/MrN3YRzQl43MmAKv/CTQynKQ05dMsF1rdvH1X7r/xANF3uv
8YGsXCuthYr3s2roqqx9jitPMlAUM9PCmfyawFi5WDkNjr697Pb+Nr2EmPtwZW4M
1q/ETsL+iXIOAXKc1bduByoXV/fxFStqVCGPxqYM34r13UID1wHgramPzOsVY42J
QxzU3bts5bnwKEuOCpHQVxZDocyjeJkZmVbdGolLdte0jb2N6DF0HdtU9vqh5uwP
lOeYn/gNvvJS887ZVg3vfzzwywKC0H7cFYvwYH/wtOFSNw2CEWczFypnidIZjPID
W5eLuaNEx0/sxpnDyslweLiqyqCX6n3CAXUX7DhcGMIFfsHFs30q7kYBE0IuC3c4
PCfPNWJpHwD6Jivzts2PKde9AyF75x4wHGMU/SaJmmy/6afxdicgmPm6jizVUrcc
JiB/vlEMYXAD47XwkQuJzG1YpgvnA94R3pykU3Sejptfno70LZNeqEMkQO6eu3om
eLk1vM7/X/24lVLlbPR9/NiymHL/mAUkdxioWwNNmcEb+i4uPtzQLtF+VrnZdfHx
C95rr6cPwO5+VFV1LPjTTjA+GAm5cc6PTB89CIoJVIVnmpKhBYN7Do2tnEQnOB1p
cQqEHE9FeBi+s6HrzhxziyfIVhTklBoMOQqOXU+4aeKCye3qONY38cI50ajQSqkh
5R+ijNBp946iT3lb71IeHziaQVi6ZbCNNrTR4xEPqA8Y7hdUfMDUelr70AhzMt1z
vSIN1mUuxMqNDIbEJptQMqvJFQQ6WDIeYGD4vaaf3urxCMbH46KuTFkCGEFWKAZm
+6rXQsB0ImzBAPNtqm3a3SkV3uR6p2nL64c8b7180QvuyPSCRvA9j810vRbLZ398
sV6Gp8Oz/koEAFnoCK01/FyCHbeadqUIq6ZGqqi0b/gtc1tqA0gZjwySI48kNrtf
3PgtxsV8sIpm5pLF+cIA/0oKEwsT1v7y+nKK91xmf7X/ISUqUwykMXUUsVVY+d91
2lJxATTTLwffZa4rGFZu3XRR6K1A4p3HlHNCM4AV3qohCk6uQeC6Ce2mnGbtKDBM
6OowTv+6IXpQSp5rbDW35/sLfS024zh7gRebcilzUmLjT5AmzMUFhkTMx0ChbyPI
8tdIgEM1Jmi8eq0OgN3HZMNzsCNfl0POjQYCwYZ5V4NTH69xNrUSw6SjdG+Nduu/
QIn19h63o+P/KxvVA5LVkEU8aWHeLEmXhMtdd46PyC8Ot50eeTdcbC5QFcQHco7t
KtXrWndCKlEI/LvfzIcQllb+wTIa5ydwOUPNJHsWynPwolrlldT+BXcucA3cMZRh
7WYAuFbIi8aGlGg/snuXP6CCx1mrU/sLMyKvBabEcjkdUXBh5oX+SwerM8oIytvj
EgIksFMZ2oWPjCTweaeLOskF621/4+uo0yMr5A0F+2XITjodA/XvFvjGRDsHX3K8
F0Ry+XTXdxz5xx/mtw/MPiK1Rwr8hI3KzzAwO+G2U/SsZREgG+ZU2nQ5RhCpkM5i
nO7iWCItpAsU5gjRy4grxcjZKwXjb5+ErVIy9vLKBLOAcZfNym/yRJJZNd3D7U4o
z1E8VZKCfz63tz46WdNOHa6n/ONK8SKYQ2buKl/79tL/dARGek7Sdt3dj46qUNOW
22ElQ/ymwi5HmYGlyvvNtHkAUpCHpyPdPv5Tv93CHBvxftF6pwiROkQ8j3W25PCF
hT/ALsDW05jgilbek+aUM8cBeKkn9frlGw0zciF8Pr6eTsdbrnQcCSp7tbkM0LeZ
XEdmhj9fPFbGZJqNSrJ/N+5Mbqwg0GNKUOpLJLJprLDJkW+zKpeHKxVCyD+c3liu
W0o/osz+poY0KJZb+lCnqFnrA6NUx3TK2wVcaHz6XVTAlsLBF4EMutLf+Kcc4kvn
zcKEqWoW5celym1bwitsx22HfRnseKOeo5v5gEkfum+tyoRT/LaCEu6xWiix0iIC
w/85xCpny5pE03CQlfbI8iJTmcr7hyJ5jyprKAt7wTIsEMyeIVuC2XA/W/bA18A1
HA0zPi3ka4eiwWamGORJhDa/bCSAr7So/WHkc+bCAP4jMkr0nv9VyrwdwjIeij9L
pfRSbnaf6ITldGSYO0POTSYonwimz+wp8AYWiVquPCjYk//UDe/+fdd18tx3ACO9
oCGJREiWyzIi5TBwb5vTH5IL5NQrGMzjPMCTayvk1dYInUcruHVFjLHqsR8G3eGE
0XMtb8/TQ+6kvUfK4AO3LWXB1WknC4h1cVctf0xx9EgcfQY3/3Bg32UQG8K78MZg
kuo9RmqHCsy0TSGfPMOTukK2esXqWsRb+s7osIkQ9dqsKVXSq+yapvAEel964ruR
2iEY5Cy47mD4U1xKbxsO9EWvez4w0DeDM+pNICL9Spx/XvZCcgvNoANcxW2nSdRq
/5cznI5IDGtsCJ+GgwaRs2p3eLzRJSWINpJlLJtrPTRdO1AfQhYTP7pylcNmRhNw
HWSIPZ4SOS8QWleWSnd84P0ZBVNJxxQXeFYUgha0pkdZ0i36IOfMRM11HirAiZYP
dfUhrN/ON59GlRotlSMaWffNPMSGzDBlu6eeQzQVyKKIM+0LLknWDyb/d3Z+e2wZ
AsxunqBVFwgxL1lOKIFYXY66h8uR5Iym/VUkJTWzSsN0fw9sPqIrf26OnrxL2TFL
hXk26WZ3Ll+mw1Rr0h54uNmgHxF5LQBq60Vs71XVqzWLZa8DmHMH3zgZqq0aFOrh
HW5Uvfz9uB9JjOU36OO8uE/6Fw6dQv8OQBpIMPMn98ISN1FkwvSrQSv4tt06hqX9
ErpmkfYQxzkJ845+9JAuloHxabKfcp7y+CWYnyr11VQ2pahpQtOS7yHTlyWDklez
EcSTEKrecczF66uJZe9gNfzI2wn4IutmHTYuPZONj1F2rbKl1/DvaiBH56vOj+ny
/7rHaSIjsHpBm57+65Scr63rTsbDkD252ytlxmezKObOlj9rt//BLQoqqwk7723z
6IkbW4qxMVHehCPGFJ+xTLarptb6sDZUU4aImcsK+1EU/jwQKK985PO7FfSPIBbN
5q64TJdK4aQSpmw2dNbsjV0cJUwWdiyL/4+luIlgOKGNpiI9j7oFQprfg7pSZ6db
jM5dTWDcyTJUGb27NXX1Hq3GU7DBOv0FWdxYJ4VwdLNvSIjic5aapjLL0l3yzw1S
0POou1TikvPVt9OIAS1eJbIUqC7pfq6g85VqfRXVnCfBsFq8fx2Lu+p/dpC5JFdD
eCAw2Y9JliLxpaKsxdsXbKCsOzxV+XMhtzCA00W7kwNBY4kewav4DOwCA0ljAG5i
Y9CBfSZKd1+W0HXb9HkuxlQUVZUfo+po1uUpbI8EwrpWxjLuwtXEl9+hjJ65zbKj
dgJG5GsjjClNvvkZnoA8m9sraSSujaLvX7pHUoT96CYwcPRi7/4yPcbX0PqrVd+s
VFlTMFAUHRXUE8yTJpil+n0qgVza57ZvVL9GfvG+9qdewXj4P+qFYgNGuZlW1O/9
OQ/aLxc7GRvr+Y6jJ1TbLqwcfFLxUo5a3PwbJVIaLnKSo5J4/sIqkuph/mqGQFPF
sj1xrRdUD1bbZOLLSnc1Bltz416kjaMgUxaIZst/RacQAC25reNfStiAdx+vE1iJ
yHQBoF9Qc9XBTm8YNXAV4CSG+2vQRglzmKWB/qZdUE1NUdQRI46e5upfUXkF1XDx
gKJK0RNOuehD19avgRO/PDCOzJ5y77YvEZRVfznE3ZQqshQRjFAIvTnjgZvYQHgH
m15v9z6f0RhujdLdJsZfTvGPgTNcfXaqBkVBzzZhZZW2YnacQx7u5O4dP5oSMvHV
CrBT1txWgjNJCbI/u4IhWaJN+CspKnN2O9UY++wH2r+/Lp2mrB+kgiVfoQV7SNOF
yjJ8MvGa8SfskHG+6QXZ886Ylx5ueDxlhZB4buoz82LaKstfFKsymbANklmTWva2
V/vzw0mt4EAfxwl9Tj7PH929B2dvcXtnJnLaf92o+HUhyxrQ5cBSZTuuIQZUrN4n
QUnCGI537z3/S4LdomQc0+ECVWmEkn+v5IvKUDeNRWDWxsHuPORjFLyrDKI5Ohbs
e/bMy93E1XozEbnnbIeEEsPbKExDx+mggu0kC94LWuzyUrQvVC/OSZo66maiBmhe
2jJnd46rOU01UHM3loYjXlpU1HJxokJX8YkyXq+KKe4lFkzdbkc1bZ8An9kVegJZ
2+dyd5Acq0pXN0VfZqZkilCUfdfiFO3492GbfQvgX814enfVd5c12duS00z2y0qL
8zQZegSu2bOVBK6rttP7jzdviPe4o/IXUR7RwfkU01brDaGdPyrs04QEqQQC2nCt
oFVCiwVJmOp3PdIYQzlsaJ+PywPN9dtzqAlGuRDmfYirHspbxfHEIy5FyiYFoMFK
A052/JPq06zGfO6np1U0kKijpvMAABINcm86YvhF+Jpa4/UBH+q3W/1BN4at95oh
92BXTUtmnW3j4GnmWhEDUpy1ZvEIVRM3XTtwel+4LP39YVTR6S3y7rbSXuwIYyUd
SFyAYoune204f2YWeb0LGOJV4jzFLhQf9KbzIoWVUUDBS/be3UFpypkpg8kzR0TH
MXunmxePFSPTF437Giiof5BsYW0il5H9JEe3cjQ0FV0nGFxwgHahmpxaqS7FQNbJ
wDEzov8AEpMPRecVEdJoXmAMxPSAnFl0WBDevLSLttcY/Tu4eyluTyXHtwYEmNO/
AL4gDxy9zyAlmXQ3Hca0tV9dC9GBQmdUaqAnm/SeHWnoeBcYwV82OlVR18L4vTyS
bkKQIOfUBjdkn7gucza6T1VDZ2YRgkw+QTgZed2XdKJvKESQKfszp0VByUvqVJFU
RMWGaFFPEkYPDm5e5aNPZldwRSLcVXHe8IvOR+eFuRA69XCm8oYHU2P2RwS+PWSu
JisY8JuT2TqR4gqIkI9DyuB7Ttxj31zb4+me9tkccBhHX8q1PQLz37JDx//mQGYh
5vnAIWfJhd2hxogv8gWvlnP2g7mw1qVhZih4kiAcgkeOWRyft41mz/qcE10Zc4jV
/2Rio+uJuqcnn0TYgnxb2NFUsSXXt8NVr90TkeuOHETtvOeQfTP6JXzupQ9wr9RP
skR5K7VdLNAvLmRX/8aHP8WqbIaf2Hox3PepWlp8cfwe+a0eScvlCg96SxAQj7V7
2RzIU/T8sJD01FaROixwk8LaystD+lSMLfcBeXWPWZDAElndiJZc1HnHHVFtjWKD
Zju4VJcB5WCnrlFIsZUfkNcCHURCE8cNWlTqPUwW81Rx5+ih6ZUI49Ac2pI5hkG+
jUfYxshtkRp2X4GEwRbsMZAtPlhgkGPUk0PwC0hKQReZIsG0jvGw1cd0cU9PDHrI
a8Davn3KREYMh6PfV9SaTSP6ppPhYC7Rg2ZIpmbs5HKA40bxcE1ZP7xZF1LObvnR
jijOXwsd0BzvYfklA0s4J4j7RvvNQhGpFd+lGsqHxbG2XtNevlxnaIq4lCNxSznJ
LTnHpVg/jRwdwbok9lS3Y+Re2KdMYn0IqWqEy6ZLKW7hEqBqoNLBW0f5nOAiEAJR
L3dWg/vPUKSSmGuzEQ26OAa8jnG+BKteRgsfAz3dNr4QT+UJSkHYp1q5UalN2NaM
onyLLreRRu2mR7iugEUrkkqGM5l4OPdUGXlYhbO8QCVENAIlwYfuMBcPZAh30aDG
V58bi/u4aeFs4ms2J93+CKDbt6Lj50ttPiP6qb6UyWKTbRzNJ8mVAhMlez1f8+11
dMvgrp4alWcRF+e/3CVeaLIgfxasW2J43UxGS6pNQJvRqqOyW+Ikoli/fH5muETs
6Mb7vvIKw9bfD4yRA0M6u3Bfsp577D1S6QoQtsWuZ8tJQf1OlKGfWeMztwl4n0Jd
bm/tepTyzi3dMNCOMJnNx7WdEp22jl9vZwDRdCHILFxbGN7Hh2KGqgTsDb4493TK
SNY3KgcQ8yRfgqf3PoGsnhHZlfVJRzARPWLMdPuyzV03VvkSYeEQw4zFbhHxf9l8
JIXnTBSh0kDcAaCBpMBSdpagw8/IqRGag7HfzMEZpTcLmjDqFuo90uVKKrOKmqHO
vj/i5Jo4TdgDAYFGf/vD0xg3kT3GcOz7qtzzdDPU1zib9u7tvFOrZcxEZ+77CKSS
2QPHpGCfkS4VCnu3YoCg/QmgHM6PVHZYerzxkwZ5jbqQeWuzZJFf5SFhC3oUdYBT
UusbcVkulVWftmo3XLq0JT1ViOY8xP2QI19aaWhOy3+0FyrSfRPpw4YIYP5jMDpq
ZfF/WB2UzMUhS/r8pyv4q+YcsQq6kqZepywgAVi+aFizuLod8y7PUeXLki5rUAk/
nqksq6DePsbU6P6C/mZm0DTvKAt1dlfGdmyTjPAJiew1GkNCOtuYAUsVQCrZgNqg
K1FkNwKuhL5eKjUE+r6ksMrG6GZPnfQIXXkQ1ck3xlty69XU38ctUFt4vrujTA39
tj92zqkpnynjOxKpOAYVDBXDq0CO5V1+tPUYqP0A72rWDb1grAK3vnLDdGnK6nRJ
wv/zWLp5dURGZFHwYwq2NM3UfC7Fldhqvr4D/4GOC1Fv1IGdIhBSFNODQSd8oUO8
ejsm6lyjF2vNs0gWQYKn1FdjyZg6y5nSlR3LaCjPox1P5pVXG7NRdCORrIN4pPAj
xguBunlPks2uV5jHFdT/oKf79fM3+ZgUqFDkoCBGDDdnx54rLn5nZ81PfdZE1mIk
GkSt7VVdifAZxRk7EllUdLDwAFtHDA1ItHEdPEyzoYcO6/OpJfFm5PdHatGvmJlD
3Qp9MVxvYCWflyn1JAXTUct6/fjSUg0uXTrc76ZJpwfz9IRliE1ZpoW815t9NPMi
8LsUmE1WpowVafKGH0wcCSe+u96OtC+bCzxreIf2/fMzBesjvg+L8aoWuc/gdnTp
bIrkIbVgEZO0psmA6cbwsCvyYQDELRXPpHoHJ4GYSkCmWlwJ3ba/2TM1fpO7xxbp
XLzmgMVdGI89wUDN2bpCeoomYnEg/jaC63V5zxSifBkOcqLmA0JCj4jRPGXWUylV
Y6BOfesdhc3xonSGmyxrZZ+iq0qBCdcFQrYKkdEId0lo6WeYcHp7OR8Zdvp9g1Lv
DxHEkZwXIAraKVbgnW5xGwQtqb0i/xXKPLRnLbdNfIzbvm2JLt14VJ4RSsoiXkJz
chCkxMX7zMK8dIQ/zDwLWIm9ZjccirY+A88Qb+2UUrza8BU2g/g1rN8vw3jfzFWW
ptu/glVuiPFbk/kpUJ6i5Ob/JbKfDKcllG3kdmvxP1McU+25IXsOw5TlhIhUslvS
Y4njnMVyD2rKZF36mtQaw6zATMfI5t7C50dFb6NpFwFLm7Imvtnw2HSdsd+hhOba
8jd/XRZ1t0fIWmnzjyMyNmjhDp7xHuYdDe1+zOb3HIYOC7VDD7ZktQ/wzP29BGJo
XbD61tdzdYFFt71zLE/nbbbuhIAK1oa52JqTNHtxEREgLX09/LE9ANYCj0eqlOz6
hJCHP3DO1iH+t82tP3k1qN0exoCIZGPAvaJXjNWfRYsiHjI8g9IkzYRsZm/3TZqO
v3OTZJlcIJAfYIIKNJBXscHazQ1qXpSY20FrbMxlixUaLeh2RvJkOhPETE+hy12K
LqZTcWhhm0qrQR11OyWItGan/F/TpoATSZ1k9seOvMqQABfxXBvDRbaRZ/8ZBZJZ
VmYrsuqsKu5MhVfSrWb7+ehxIy95gHnQVO0FRg2NEeEnBdpqMfTPQu28CGoRShv2
G2fAXAXd+z98PnFSITPrGtSGaSaj5F3M1deMl1v11WZieJ07Nf8CBLjwcbvoQcIM
BF9CuFUu0NdbKynaU8+5sU0LjM+5mQ/5Wqxyr8CxaTeCSOJMUvbBpV4+fDCxzHnR
USSU2c6DTER4jIHEQxRaxFTKj7CpQFpxmlDXsqkMM5VyeU2v5L3vsfN9dpSWcYs+
LirUm8Nps6xsWvzQwEEPizXTsTBCU75jfk5hE44I6qRcWgPuHkJdi4GTToh9pGtZ
HJj3K75HtdwYtdqmM9Wz3Z2baDRbwxuPo0Dk9fz/zTcNSxbLn9R4mmFvQl5JwgwN
npq53b5IXmmk7+Fn55E07TXYkKGGyUPO9XS3DcOR90GXfkZffbgsYB18X3uJUGB5
knyIL2Tt2t1KS1NtEp4nV4+yg0ln46Zzo/+dKg5vwgXr5z6mhrzOldrmUMDK11lM
lJQZPurj9vyCJWR+Z1tAz/dHD4OVv/Ziu2iKqlYR0565EqddzkC+0pLpJwlZP430
hGCHo06H1XyTLHTHjjUBxyFrMJ3+lHSxTsTjwca2u6CrWTqk61AhKicr0kbDKm32
TqYT07lJdP5bcrV64W9rPLOEsWw+IzI9RVUpzO0mtVqB5EOGWtV6haBE1RPd+P1T
GjCOjUUW00IifaLTvWsb+Fx5J4HbcW88JtKEMPygtOvYtrELvDWyiCP+KSa+mVLM
QO5Wf6PW00CL4KJRU0K3/HCj2TYj86fAoOCBucLakqVKGYHfXoRigQxHbCI03Mp5
aId0s+Ffw2DoeN/yxWnAyoJqMJa6aS+vbmJdBBHa678K66x6dMQAiAU7fmawHDsf
D+diKCkmOJwKlWPlVPYAHGBrrd/EvK45FasNrDzyMbWJvgFzbf3HdhvbKtQTnNPm
RSq7pS2lxDYrO1VPpQ3IvuJeZfy4fCHDMn5j+QV3chdFGF3GJbP4uIItqvSlEbx7
n+vl77cIXyc+GNNQ3TnOoP9iQhrVqCIg2jroKuw+QeeXvuxNTpH9w9vpEubRWae7
nCjSF472mZByNwLoKiyuKpzB9hmbzNxV3X8MkKF+Ap8q7BX+MQaYBSF5tpxUurWB
q8csj3FC3rUnkHW20lirku0bw0UaLhYVRKl+qBFK1+N1qu+XXOF4M90gG3wVO2US
J8D9gPlwTb8ZJxfL+0gCLd70p8EvoaqTo4r3WYMXz1x1uA+74bNvksXNCynD4f/V
X2nYFQDISaV1lbmSRt39uHC9W0YhPNcYa32q/8v0vToruhkKjp0Tq2kWDeDz7DxC
Y5rgHP3jQgl5qBDyOWcZFB4Tr05Vn4zQTinLZcDwWpK1r7JBZwNkAOo8rNBMgAsr
ggcBarU9GipoChWTwVSdl3JljhvY2lvhu18y9GS1tr5Plj6YEVB1KerQqsZlorYC
Rl77PYet8rRQICJGC0mQfP6+hawNzNtnMxC+8BsVWRBuCbeosQtemzpKrc42WpBP
gkHEsCwez2euNn/ZkM8CA0/gTVvGSOd1u8lVJA71Ll9hFcTgZPyLaT+SBFHjjzBR
VQTzOPBAmgUAv8euvZj7w4EFgPDb/g7M71rzrkLjeO7cUxiQNFzTJmDrEdBwLlSL
xYIfZ+OVDXkMmMm8yASJUwTsc/UVqWIpOmyq7HBHN5rUtpSrxP7+t1YtIEN1Ua0t
Qvstn89wbqAh0UkhG171zzhxH4e2yY6FWpZkhTCBTcLaNZ1hWkxQtx9iKCpGm+mp
eav+UqWiRomU2ndttEhEfkyyYufFlrXUrvBiKXYWTlayuriQLIIIq49NfcY1V6ye
p9CQYgOGYwAxqFvU1VNKtoESKYIPSbd33MT8RR7kWBEH72RtfHh9oTDgXjwnIy1h
Bxn/+/eTIJQZCkLEfQXfCRWyXOONwVmFIbS6LQR6XmqMQycD9/KXyICRLrNtPrsw
+DdRn0R5i8K4/v9eD/1KE9iOMAgEdMjoBrLbf6z3OE2Zr4pLdQEnLxii6iPO3sXP
IwGoRcsbGvcbpe8Uofdp06ICjgHS8dN9HuzodmxEQoXZTTvreW6RH5J7iHs+bN0s
OcqwEtwLgltA5C0klNz8rmfk13TWqfgxXT0R3bXTss9/YGO9UAneH0e/UBspFGhP
ExUyuIjkk61JyO7De0vTdGW2vkDnmVlP5OmG1JTSU7BdgLu+v6rnBaNSt9mpF98e
b8k5yguBlH1XQmrbXg0k0Wie2Pn/ezMQ32krdcJgLVDr4cnby/6JdjQLylV6eEjO
C8EuSDffSVBpL1emJxIoF6ovbZj+16aECUf1/bm+dFyhPcecbUdk+hPcWwm3+ZxN
65o21xGYm9ckrxP1oPiA23p/uj2FySKayWLPlEpIpsHq92tr99MqZslB8VrLF8lR
Gx1kncpAKRshbJflKIw9q//Xp5nyExLlCAW1o3/sGQqiibj07hWTVRBmJ/jB/YP8
bNlyb/jTxNfZbzO0hw78zCR8kqCSIAbtlL2Ogp80JIt494I12lE1PnCvvyCARV/5
lpvIuV0Satb/IpaFhX/uGCHOPOrCphTXiFVRAN2qqNpyir3MFhfaYxPrnTy9swja
JKY5jSG2Y2pnRnxIkYGB7hT6gqno2cpuOfARrg80HfwgOUJxn3AHjP3n6Y29Ku5x
111SrAVbo+6AWr3TVtKj22jXlXGwFTPP07MDfHUU2WLzNrwF092RpU9k/aSGjCJV
Cg4AVMr2Wa6SuNYw+2kVPftgy5KJEEkcEdQFFWomQ6tHn9Z3Zuq0ESvLLEeeOp+B
ryx797DaGJm3xNRI/1DJ0nX+Iiwb0pJR8IQRNJDkZSYJKKIygWwGsZBdjZCoq5Ga
5BcMQADJV7rup7Giqzae5Ji+LrdSFFKADlt07VDGd+JSpQQ593FZ2uggR6rdwOVs
NCm+GqKezKznKl6Zi7WgEXpnHd0+txIXsWG8Y/NPRvUa0+lSOu2F4gnmDn0/vgy1
RUhG210WA6NaqknM4v3hsGKl+WOrJqCKiCWjKSIwB+DA3OF4QJ+LkQnA6iaofnd4
j61JBAyxgahfrpaSYaKrKPApWMD80iSYbkNaY8bFRCZya6m9KZJ3vxPaDWxi6EZa
lOI5xcBpuBPRzeZI3kwW+hvzB0isCde4lf8kcJ6wS7lkemoTGdSCz797oxk9diR2
zd+P6ICCUCpFhw7qbd0jk1JvT7vArs3tPmGlujxaUBPuN8V1hOx5RVLgNOQVeeId
jxhkmfoz6q0oOzO1Y8i8SQ+AGfoI05i3t/37aP3KSUnW1MxS5a9swm3weIMd4Ebu
iif33nSFsksKoWYbE3QgMen5tI8gnlBEdtfhpJtUqU0O69ZjOt8XkJmnbaqeQAOh
+HxhZ4FjYbGqMaNHOy2KrGtKrXrOb3HWDJ/PRZzbd8ll76igN8QFlQpXsAo4Y9zj
DnQEqGvCH7C/ygiNQViUTbp/5sUu1/h5RXjJemu0CxfuY9TGacXhgRIJanDeEgRP
/6AIa0EMwAKbHmcWPp926Utqo6CrVYpW4zRKYRO5RyvPYnB777qk6R7NJSGc1YLP
H6hrbRoOvv0jWfK5nGWxAL0/g0bWe2q0uneQP8cpkp+uD6jB5pXu2TeF8Y+aG93f
NbQpcJ7DsL1y+dLJwtrxRP68OqEPkACfli0YiDIaJn9ZmSEw84ZYEkOT9ut8zuXM
HaCARUbhBcphGlU9d5gF0PFiGX1g9KEjQJzKl0XPVpx50R45y/gujvLeX/znOB2R
oiBA5ur41LJEt+bL1SLre4vU/dCNGB4fSRmv56cxrMZG5K1kF0jC5K5JH1Z++os6
seJjok7ivOcm6CFUoCEEwchzvjppULga5kwyZjcveHDSLUj+Pgx9r7Ktbn/8DvOj
CdFu/1vFw1cgzRBrCMhFaJ6uB2uZM56hTxlr+wqr48C1tDW/0LkD/T2YmIYjSgGo
rbdgkW3viQ1P3C/3uWVtUM6QLWAFBQZGUmn/avvfKoFw1iUfK931l9B4zC5O4Fbf
hcBEtK1XL6C9FN4wVThNrqG55T9KQQAsX1h/MoF4Kv+WoVanxPjMYl/iMxQR5vq+
DcNtdR3nfKuhbgFtt6XtICvvKRspASFbMHR/paNaquLX6dx11Dw24sEXIOMPC+G0
KarVm5xbLrsMvX/CtJdR0HJaJqub60Q71A76GaLwTk08QB99fdy+KAffoYNSGX6S
Y7via91mrkRMLMt/he2Tq63nNS5OVT39qGp4WDbFE/FeY3bxSdAI08jdL0dqKtMc
j/9FVXVnV4f3tk1LAOInimRoNYO2QU1yEHZNbKnL311HbFtYWM+ooL9pvXwHTAho
l7EHPsCHX1W/iO0BFT0UNZ3cYirz+SaA2osUqaMoz+2sQG1UY/EXHZQ60QMweCdK
QWkpGkvNyJnsQGM+kNA0crO1wb3ktnJ4ECc5fsxCs3OirMomN4Woh+WLrsAw0H0y
1RGK276vVpwF2RlBjsTl+wtSv3f/h57mo4chm2mvT6tWmmfUJ0mnpIOjtORlhbY5
Ct4/esIzrYIgZ1+AngJEGJmondWTtjD1ESF5vQdsCAZhRvxJ0mToRc092BrCen3O
XKhAPFYMZ4STuS0bhMcaC2H6Mmkb6byR+b6fXQQOUtDyeX8KyNY98q/YYtA7HANg
3kN6IcjN7MrumhOnNNIfC7/n8NLrG1hGO3vybRlABOfH2zXkRgjvhVsCedfXpqJG
+T1bUwe9OPKgNLbNpkpyZMcOznf6Qi8g3fgIJF7YsD2YWF6UhMSX7iHHbUGiih4D
h5RToUPB73z1Z33Rg9GswwBpFjQNHKcRxBROIMCQMZBbXsw2TLvePkpjTDo505oC
EPM9Pn45Yde8l6lxjsKoGte9zMGvFNU2cXC7oZ5hripLy4+b2zwn9yMVrCci1tGk
EhuQ+4EUt2NaPitczUe7aPKB/ltlQKkhazrjvZo8zZ8AsoQX9kZ1cTplFMx7ArpJ
oHJ/92tCThlSy9zMBZoGe94OlPxQZ2tlMB0+dWVmduw+Tac9ITEIxbj/F2IeBCvq
4kygE5U+llFpbQ/zXKmVt+1MTGzQJH83Izvz+aAj46ZJbBcP/81lNzEi+BeLNw52
gnoSBgPfGpDWzDqTxFqKWow37YObjXQqhhokqOJRZED9deebyukZO4zBmInK7fGb
hzlp1T5qLLGN4DnFHBEl7u8z7RUk7xMADXScKgWdp5JjuQWp8A162lUqYwu1Mach
IuIgXem9bMy+BOmWKNl5hRky+XN/zl3mH6ga5SZPAjSxWUJqYHMQUc5pHduXGlMv
goCizfTwhtUGvmo3VOhzNn30JTlnFLPWvlmrzzkeZUiE8uJV/JD08H/hTY0idczR
9W3lAnNWOTpJupfkZrOsudFzPscnRGOkZ0pzTUj0n027lNibi/F+U5lByYLLjDb4
lpRhEMSPvJqNTQ8BulDLscvIMLQ5FdnyyhImlVu9XDZJ2LgphdYD6wX4cYlpaBT4
ohqQBOmyf4fsvnE1mDph7ICwnyS4gpVIjr3XLBVTCAJyVSgdrrCdCJKb7G7wHE57
4AYKYBTatnyJPHw9GNHD3SYrFRS2k+JnOyrQYTpD/xBwjUShkn4SCYenmAUXjfp4
yRMt0BhOjL73FmlwEkFTnVhA+gC7lV6WYEB8c4iYDPGLnCHj5R4375heHcDcDvoH
OmUSd9xaBVT1YcN7SCkReUK13ACKENYIJyeUfAy7jDnXA+BmXhFJV1MPuV0mVlcc
1MiiqQyN7dG3VPOEKicNw3+a01F/4sVdE5u3cj27SoGmAz/fmxssNvRKZ9J30ala
kMX6bkTOg3Qta5CLl4QZ0lulFvkQAv9hlCElR6JPs4aXNoHss8KPti1yZ21nKHKJ
6DtXNGU+pUxTqr3Dy+yGyStndoweB6HkjmTaG79ZCQETwSgQhaOHO37sHz3vN6/G
N3wnmWRkVDNeMAM6C+awwu9Hofp+5NzHRga+kzNGsJL7IlX1rryXA1tDaPrbxfIc
o1DbLoC6TUpJwqp8EIHv2kdAzgSyY8jacDHAxvvHD5gUvo0VFKyxidRZ0dm+97Ux
rjY35+54kr9qTq61e8F+MfFR+c/yRq1BzvXk1WgrYeqkQucHuoHs5LPDQp4rGC6I
GgDZADWiuz1Fn+qCfR8MNJ+TqQ3+c060T00ilCGFO3Xu0/npMLshIlL8t9O3brHN
XVg5zfw9z7R0eQmWCHM4lwpuea85X4sMusJNz2q10BKKwA47g1RsChsbn89FTtcM
ubvwSL3vVB7XX1DdJeAi1QKs7TIOdcz6SKOKQffl0LdbUF9dO3QWEUBJWThiockv
6pktWXu/HtMverF3XGvnsiEO6O55DGzemFcyExYXqHno/+JNEKplgMdgFMYGESgm
JyCJmEgj5NtSFUhTsTvf8ZA/LKOAlEzFC4u5EibCuO5BmbkYNFfg04DznoPRlwNe
9nqWDGC1l0nPCu4bIOYDBvlXaZX9KpW36DfAwhsC/cP1LhXU8hKc/6ZG+AnbujLQ
fFwJdcaddtMQbJofc/RmqEJRURV2MTGBKrDmpPcVQh+dJKLOXzzjG+zLXQgMju6z
7W0GRqtNbO+QHMmTKgzSR+25TzgZmbYxW88/aE38vqpabGzbY7MBlDGP/AEKkiHH
Ht4p2wCS3XsiocBKPv9rmSoqissdsHGnxYyAabYm+sep+mSVrpz8EQ9Vvf5tjMEt
4dtzi2fo4sJbRHy9x99uQVUDG+x+Q4MpTgWkC0sqn2gUEes4xmUKNEJsCNvEM0Wz
I3bTr8bGa+edAuUmp9t5EFpcFIzpgsKrSR0gRW2s+HS6h7mrvCo8s4GogVpPGT+I
2+UQzenCRAsq+Z1b6VP6XuYxgpefwOb04K+Qmc0Vw7R6PbdAcFylk8TYEtLrKx9t
6Dg+kE6KwhlmzEuIDU9MA/DiRaKbgQmadgP6V4XA4h3bHpB8DCI6pjQf34bKNDD/
RKzNXt+YE0QdtpR0DX8LmPAAvT5CMKyjvfVCJcGDRtUvJrUCaH4pXYemQk0kPx3k
JZutauysUxZ0nL8QYnORAzKAeEXU6y5GVXIYR4imRLd29XdyJ7OCqXZygE7/TrZN
RhyjJDXZYjBpMPOKQI06d8QQqKlzZAAJF16scj2kwufYwppKFRmMuW7GEJymwmWF
fhD0ZFeZKBoSdNY1ozReASGMIvaFJtWTxqvxA5muXSttSwM+Kkswhgtqh5amZzr6
cGIC9VVvl5cQE+Gc7Jw3tL5NEI8VYKHv08jXHEQ1nTQKKht+l4+ZkQqUXmmYti18
WFMOoHCLidO8DQPC26PVYseTMj3tobdCgzw4pQwMtmJAvjBaTqyzoc3uA9BfLDkm
hHdV8V/88Tk1mDetT+idW6+KnPkNuKSZbAWKlsw56MsM5hjUhvhS14qwLqUBIVKx
qAUf2jSYAfGwakVQpiiB9kfLw8KE8mZ38SGX+S7Gqk4nfZ3yN/Y+N1zm6PEahDiD
trStk0rR3bIRy3P6xmqHTVmMQ4Z9BMYbBGOOC5cvCkw8pahRAChqsXaO+w/Oh0fe
cNkk7wffyCpVLB3CcfZcIKR1b2fhJSv5YoqhF1hjF0arLsEyLBSX9yQAYfyk5Kui
JqZPRIGwdtPMr/HMcI1CWWad889zwpTpswxag3H7gZ7Fhd495z1P/SMKG3e4xI/j
BSn2kvPvBFW5JSds2icsxFi7KH3+m8mPai7h4bBSSqq7I54EglrXSZVq1KBoxMl5
shnBapCyuGj0RmyQ8xFSKi0q1zgclc3Gy30LBv0Ol9oOtMsqMlB1aPDc4w0/hShv
lETJoTdXcuX3SoJbf5PXemt8tfO/BI3aBzArOGpfDBylvgQu2Wb/O9pOtspPBo0b
1bULsMivZZj8GfQ1x4D+BLh86epXqGCPcwt26QFYX+aLVIHwWGkcoDYb11H/XXWD
T+ET7cNvnpEAab2B47lLBJIxEqGV7VdegdyFnVk0qcYL8cHmARsM7fo1dzhdRqnl
FFAceazDpZOPobxOxQc3LuUd9fg+N3ImDy1epO24O6MM4WG7BdNNbbm3dPUB21Wy
AI2svtqvEashK4cb/UGRuixhIIbFynSzoaPW2KUIDs5L/ERxTarxghjyovNuQ6rq
aaAgiMhJMC3ZaTQA+FBPxoADUkT+sM6B3VJbr2+YAuC6Rp+VvkZp/t1EYgTVuEWC
L6cE7Iqn0yFA7oHE1FANvCJxRlV45MHsL+WGHUp3DhLaNof4yYFJnzHIhi8HiGKD
o+AMttVwHH9QTHaWhAFG29s+tNLnUk5ROniGxPHL0QVyRbMJ5YkiOD9QXsFylxKU
8mZ9vjY67KO67CQxf7k5rVtTYGG8bN8fPOy6rOMBSjmkpSRs9orrSz+nTZ/ESS7M
EifCEp4Y+aB8SZ5Fr1LpOtVlUTdDhdBWSo/4K4q4D42mKfI0MWfgzOm+BkwVFMUa
xyid05QM9zuvMqtWSGAJvlXPM5HMAqThTCxB29HkeiYo78UGDJo7n/2fW1fYrukq
rJvnGokYIFgQEECyuaECCxWBLPrX4D6CkqxrpZeC+VXbGrrI5Yjcx53WenKgybo5
GcEfstKxld1lzPxSHObNTzeXf7dYah4NGbADGysKstS0lKtvEsqt02IpGahLVF4N
pN2pyBwUpYZZJ3Dy12U9yxmjrlCBQ5vr8AambRC2sbD/UQE/9kQcHSoZW3gAyK5R
56PmeS2jS7SEIvJjdIAYb9le+ovupWQY/S/sjbfDBgjqwSwP0AJCgj9hmGzWqpbV
xv+Sj0pH1hbuD0pYWRtmo4mZOWpnTPtdrT0vp+RTclX/ll8Z/XInQnUsktTmviO2
GWMxzAbnI5tYWoX9JqiDVh4XDhtRTA+rZNB34GjXupq8ZPgI8I5pc/dBeFSZKYrX
GgxHy9ZsHyGiB/Oq4Fo3sPfyMAbtYF2J1AL3wCnXfGjtSx9keRnCXJyoEmLeI3Zj
X/wckHz1vQfOJHgPTW5D6r76O0FDRFAmrqDIPdyGy7cWjuzq5FKEuAuG6OMeoviO
vIdg7PAkEPttcqybWjBHglXZvUY6I56aTejrc4c1MfF283PPOfWxYky4XOa+hB/j
bPnQ+ohnCwagYMxML/WX/UTd8BKaxFDAbiH2EEvQgbUc9BsgyaThKKrTyuQ7B30A
OmYEFr7O8HVhvkxI9L8PXAnCu9iC5f9aBoMcNgcbtXany+vCWCdEkOb+ogMRdVMi
Qg92ZfIZJ5EHE348lo3TX8vRDu2EBZlaRAjq8SXSw06l6ZelExnfDKfjDtf+u9BR
+8zZEPRTBH5c1VUXAqA+r9G5Ia4Itbbr24SpPY+ziw83odhQ37fqlT904H+oJv5w
PTGMZVn84r3JSXMt42MWhcryRqE5Qi+5o7nBzcmRudmg53jfTSLgLNVYNvpk/Kfm
DU3B5OtO9z+qrVRk/nywASk/aVktL7Al3h7+hMna5Zvx/MfTvmJCj1V2xWRsGnZV
h/f8aRapKBH3oD0z02ibMtcjiGW3rWOuRhcYOFMFnP4FeelD7SazyYKjtYgjeWGd
kozsauNUB+l6PAXa4JGbKofjAnBjU/i9LCxU8q9lRBUEcVbU6cnR36xrAmHL5HxB
s50J3v9jfBfiz1OEEK6oj39XR9qfv5hoEvVD5sc5661OIRBcwMRo6xbvUqRuFcgS
d0A97NWU4TlyhQFj5TRRLR07u7DedJYK3/14psDH0cJQHzrzCIM4jPL7fw3lXT/V
nPdNVBMMg+bGvEQkhRGPyW1YlWkRKPa20n0FdGbxq4/Q2Pk6PHBL1EB+mhKvglMC
8ninFtt4cKIKdrTxYqcewA9yfOImlFcxgyJQj9R0DMqzWx+kAqexgfuJW0zIk6c6
ZK0Sqr7tAbF7Qg2enrsUbK2DbElkzGnhEM+0GdO5paEmcKfN1WqLrVS/ZVbVsYZz
PVmClH9s5emtiaXGfq1ntceg8B4OSGIsB42QfGBTIoLrGTWALODUyiAX4CVQuy50
yD8y1Bpb5zaQluHyT/g3QGuNOewDy+iG46rxp/yBaT0iSInwrtFP7BJU5y8GLNI3
Wc6+XphBKnuEoAe4zmXYdj9FwqmApgcnQUJjQx1TLYQtS+M+WdAIRnDjNozrGOgc
oMe9iuvkmJi6t0OvTbZXvx9jgOg9++8Qmlzg7rUI08DWJtrampH2WSOq4qeGFBge
lu1rCQq+HlZtxkWcNa4qPCGfvylJpWNUiVptmfXevITJJ7ZILFK7wD1hYHNWR+rL
sltcw4i1SwvgbK6jTbGhJF7TN6OEqF+WW9tBVTSokl4ptBWs4sVwHeJcp9WhHrZ0
dqJ5y4dF9vzJqEQqcnxACH5j3JmncDhT3av4hMHp7M3fR89Ss7ugyiYqI3+6nQPe
HfKTKyz5zzIWMqD5iwo9gMUgR7zNCkJgplQInIjqIZVTgHfEY4yQl+2y+1bq3kOf
NB5zDU2AwqtOGc4m4A77UNqEPjCK35CeDYMlLsDXfG+7alw/X6xvreqs0Esd4ZXL
Kf+AHOX3B4kN44/yHZFGZsCtL/w49z/4X8Q7sccYdaqZbGO14r+ikolAFuPZsrIT
HOKfArdcpTZNrA2DSqm79pgWAHo+LM3jbzp3NwWhqKK519W7uB5i+ir1F8PJqRdn
ddtE50+HJr0HdqZDYGlZLv/KDLcwkY4yKIzphNKPxHBMgISqht4Y+aJI/LPjyjW4
LJRaO44j0fTmpr8mYbo49csWebE9/AvdnzVRXnrG64DUhZTFU1RZWdtzrhS4ubfu
1slPqAUHZmOw9W6q/2OdU3IinL85ZdcX8DcgCRSw6v92GVJqfNX8VZg9XKXld+Fo
RDmGrea/wc1pYXoPvjQ/yLXrU3ugdoggGFbMtXGZLv0RmEG51TJ2UCY6CO1IvmFB
H6pRq5QYwYA20XZXP5HJFbbF8XzSCrrDcz+cB25UFdrjmESoqZjLH73vqQTpZtSj
8FtIcryWK7SyTBCIDutpGQFWwz8jBoy/yRHYCQD+4un8dxpRvtfxBKmqITmty15j
+c7wCAyOFTJzWjW58GGJptcCsAlo6PF3nsYqi8atzFuNZATsWtKQO2eX0CSUJmuU
PNXyCfHDWyZzV3sGCquEJhxdy93DKnIToq4SGjtqdnIms0ASJEdfTUuKyS8Z/Et5
rKuQkax8V+jjXXUzdiiIKhQ/ZSu0kGgncouM19XoI0tgrVl9a3VJTK6Vpa/3pE4r
W9dogUGlx9vqkDzVtUoqhpc4lg+H9jc6Te+Bxb0sn3CpQbaTVY2XYlHBauZPaOai
Y9zmd0khf+yTg0b2kbgojVDnVpmI0KRRuG9dGEDHpZgPAGdICDWk6m7EO6OqCAF0
OQn1zJqV9L3uDF592Kz3ZAhIeYwtvxblL6nXR/W6rCXPUBXrBtvcBAB+nJITcaqU
cP1X2l5fzhtqGaqoAtaT+S6Ics0jiafJNME6BHldDS7gkIt5+9vvbpSLqyvfjtar
sJPELiZ/J1VEUtjU5mwQI318rXS0YnyWUf3YV4YZgJC9DNR/Ii5yf+bekrCbUH0A
sAUhs7D9OwAVlPMzXGrGTLUMCi9/JiwNFATBPmaOOY+qhu0JzMb0foIhFIKyYiou
0WNWNOVQyMpzd2oMnONGMohKV8EpsrONL1FIVYn90vZGqA8AV+R6+nZ0fkpW53wq
6OQQ0mjzPzNfwe95KT9gmtH+0FZljMA/UeqiTWL9awRtlRGILJW2ozRQZ1TqBQZv
D8ADOS0VthE7FwfSzdjhdSDcnJ6qkR018RdxU5dBe3CfDDP2NoE3OECUG0kNjNff
BD6dB+WdS2VXPkzH8n943ol8RwE0TzVuckhehOEHn3AGWb38yAiZHQp4HBgcVISz
gMFMkZhwocM4xHI+WEtP89oVbHSIjukXn9Q5oeMza8LirvO7GiheRcs25LfNdDaf
kzAtbmbzyID25Vulyb8HMoPKI9Vm3IrrRT4JIR4LN0lElbDQ6L+UYU14P15GWW2q
W5Mr5+UY61Gxihg09H4dlphhIzYhOODffcZy38N6YSI21fKsq5k7LJEyQJimikx9
/1SStxXUejoW5GijkfILwnhpjxanXBaQ9D+PUZOIFYqNqosoexRWsks62L8BLRGZ
IaaxyEF7+R+j/+XBe1HdG0B/uaD5dX/6EjL0sb6R8YZITZjtuLFWOUafBQS6xwTl
U1fdFwOHHsQbhyqkpLCDwWzhPsK7D4gNyPkJMfJ14bNZQzBAkQTBW/PkCvYQp6eR
0w+4TLjEpvRg+rtGsIuF0DkfM2D/4Nwo8gFiv1xGNitfYxMU115lyUSBY7Uw/7/0
cVHs85KVRM4js6WNjv/AmQa7vLLZcvKZZ05QC5f3e0GxMTOt8K6HCp2141AzfwZD
Hw8IrGKtqdxVUvrxtPICvrHVRAD2tF8CJ/ai98f+jqH9W/egQv/seohbjot6Jz9Y
23WXw9fShPZaueleVdI0P6t6MGq32YByPkazGNbGot48MivB840UFR7f7QHVBkEy
UdXbODocXkdOBP0ONNanALNK9dRBcuR1V2zOv00q5ldEKikIOgNFdZLD2LSS08U8
/JBR12rE1R4FADuvzEiO5DCrHCNk0kzWDo9wdEN7lFEybNrljI6YpvkBBeMHRM45
P6eVWE/0DE3c2xfVJr8rX1A/PMiqE/scou/iv40c0imS5VWNs3+bT4MuWes+Im+3
6axt7o0KzumNS8kllFMbqZ4PDic9RLOHvjrUls2+bkoy1SZYwNWcaWesueol4Bdh
AhyF0Z2g67F6a94XgAfP9JlOjwgySgbj55V26872xCr4TbwwYN8JylnqenEyD0fv
aozSXtmbrG6jnFHF5O4Z/Cr7KLswV62i/ksFOfU6xHUrXff5c30Gsl5F4IVesWt0
jqeO05IkOX4XE1qyCYgHMDsZOFBvYV5F9Y3xPopnHAeHXhtImYC2hfOrG2heSBUu
Hwr0PRpkxpbr5UBOWxSRtnVjusTrjA+WnvmwTA1d8i+Yg5waBabnFav6RR+AHV8X
l7r5tqSrWCOPt6JsRY8byNwU55sXechBIbCVMzylhrJbvaFHArIvaop2LFhWIuAN
6AnUldVvvvmAjJI9MwdxPHwBrSc7hPzFnq3LhY7TmgFGee80BogcfPJ01HksAF8G
YtEiGHV0BE3y6Zf+huhmCvua8ngQbJsvMKBW5B4OqFWfHXR+imAWShkeaoKPjno0
+SNRH1WL7mDaQleWrAL7rL3RV5nIBlR7CDZWRxKnZYwrm7VKHKfLtfe3vIoHMhtG
3+bRUurZvt+bYhCGbDVRTnmSX6AGA3mDle0jHdiUWFODo9fMxwxT91rHDjhTOMwj
ODir+tImpdloi21h5VCUTQdy4bLfexgly53MQbrJuaxfog2hYs7QgjR4fUQ0cYD8
29Zf+X6zcUI0iO2VIP8AJcHxV33jvy0500pLoCDfL9fRAHXjsTF3jjASlEaVutQm
BFdLqkweg/HCNfs6uDwG7DVVINFOzq/xyCHYZIqn9xSkOmLkc6tl26+20xk2BAcJ
5wSbPTqPSKkM0BdMmH/jDfnqtpt4yEntzIZrIg1/GE+p7Ab+9QiwZ4a6756g0Q9f
VatYIpHzOQhg35T8o4db8hqI/ipy/1cfbSJ+H6lzH5wT1hOijtYRuJtIIUSBPXs7
LSFZTtwPaSm+QPMVtExhA4UK0UgISPwwsOroIjS/AA1GiZNvpLfSbzUZgRb4DmGz
zx5nZYr1S7HePKU0GZRoCFCHti9MV+xOR5XexOJy5kfBJYgby4W4z2fgDYiHgMXw
tWM+1cVAJUH0XCv3Z2CkgZZWS/Gkg5QMaPX9uSA/Y+safoYfkufIEWrgt5bs1dv0
cHMA42t+01ZESsMyV3RdvNOmzJMqrtfJMAJ3khyZyW8VPJk7geYzlFcfAl8+Fnyn
lBVYjWDSnXbkdqpc+JO8f1cJHB8UHsWSxKqTqiTy4mnJk4uMmX/1DUxrMke4HaQ1
ERMsYatWSbvWt5wQyTt6ALkE6Yf+4BP+73AloHODmqARSK+0nXqQopJtNAE5WHOi
pqTf1Omug+Pyo6d652YVMyk4FwCrJjgbRrWOffIwU/Gby3D3bKXXW3sY29Kov5LW
pRjD+Nbmot0pt3oMaruua+jywOU8wyBg6UFU0sYcXFgn3NQucOCEoImKYrNY8S83
XEo1o36fwhGL2LKOduzk4v4OpsTiS3EoK7MtJngXTb8ct6Mykok+2cstvckun1WP
UrzFQjjcDGu6dHWORH5LtmbcbjDHJqZrxWb8JGS7VfxB7Zt8iCCEFm0n0F/ICjNP
9mV/PpNBpl8lZympYvxlbu/SleGVTw59mtig0hzlcRqBiJtIW4dMeVofN1tb4Dx5
J2pauVURQmn4Tob+0mF0WxGyxbqRdkYSMeleZt0aDegEplm1J+4IOzv1SkcDwgDc
Nkh8EOhj1qlVcxk/hShKOUI5DHBLNisXPBAwX8Gor0xpiZs93dtZIlrHn+GddCKt
zH2KOYSi2lUAm+W2myY0B6T3fJjUh/hx65qhW4eLpNZfHQw2wYTqNF0x63q43jyk
I1ae5aTwGfiQoaY2XQrx6p3z/0Kek9m+om068LV1HMRar+sNVxoBjBntEMBAZ7i/
BHamm8NrsOJ6YI5vuormnTxWDJV5Gx5lXiHEZZBbkYKNshLLFuF0nWSNysvC5JUz
e/rxtNXttv7x0vTE657+XRkt/2dpFffmOUs9NT8RChbwBZyOpg4ruScj9ksvH1m5
/tseQbrAXexOKqc6ZIW3/zCqN5Ii/Z/p0kJyEDwz4rqCTGeQKCa6kicSXu/ePc7x
MctwdRDUyBa8H5L31xDN5YAdPUI/G7vXBJm3waCmn8K9mr3WziuJJxIK54zdrSHw
d/OagXOdUxmCG4QeAnOC2BXC1sENpj8xU7zWJWjF55n+WCq310OXYbgpuHqNSKxV
RsLon76f+Ru9fdspm5uPejrqnhE/OfztbV5cs1BIEb0XyJ4sfZMVQTgcyx52IHKB
jcxW2HsyZKdFzTOuvu/Zy6zLduufnnHU95FuURJVv8wog36ezH8SN/43HsfLpl56
lmVqXFJEetA4DbHRX9YpyNw98gVcSfW6gtGmcfkpJ06McAmTGby45LDgBpPtD48u
NvUQPrxbdyW03M5QKP0Qtal5TtJdvJlGSIv0xRK8bJsueh930SNeIwYWa4YzymPa
+qoTti7+Y814CC0pEVlQUICs9kZHR1D/fIJDfD+pDPf0XY8L/VjQrZoL7TyZMQD6
ekPJPlkO5o6cL37nJLrlPlG/TuYfx06QZ544mDbn0C6JK0PUSSxKk8p08BabYg6I
7fEcoe/M6zR5S3t86YAQR7FLkzJe1GaoHUITiSDx7zi5/T0DlGq69mHnTfSaVub9
1xmXAttpXjBHH1NCCUcE0Jacaks/cZxbL+7vR88t922ZI0APc1Pf7mma0jsZ0P63
9IQO8kLD5wmixdfzKa3gAGPvvz7yfEhm7xbZCa6FhaneJiAWcDUGRXdxkEkXr6Z0
SF9X4/4nKHGeqcR7t+O3QGEGCpv4MSGw97CEp5VGUX1Ti7S1YNQIYgy6ZF6TSbrr
EBIu8HrHab4LTe/2kZ2smtdRoYxGGbMiQ6a8/eS9XcmWJRc57CUoo3JPPT+4LwU6
cgPE3yx+/UsnEi910FBETxbbF6zMFSUGA4xAEgD0+iJiVztBYUHBWyKCFDzuQyV3
18wOu4QrjPxljwmsxt4zVeEtOAgjZPkLTHtSH8hTD98aTkCd/ZADGpb0eR5rXmry
7DMEjsk6KhLvmDDj7QBB3koGrmh2RxLGH8Z0+aatiAIX62gxZEpp0zjj8CcoVd5w
idrIrP8tzveeSrv4LU3W7Havc0Eks4gQynpxiXJKsQNUXTfs7+aLqQIVLZbXWaIH
nNb/iiYJ/mNCj7NcVQ2pnub4bcmx//W1xvF/xdxYeGLq+GWHG8dE3evS1EnWeunn
UBeAVfhALcT/6g070UxSZbfPtt4IW6FnzBiuEfG29UmCBnAGGoWpC/J98MVZ0ymW
M2jq9lfYWcwqkwBAgARlaQATGt1EaCOM2lPKDSvywuMzO2KkAMgtR676HgmUtMfT
Y4OC2HtacLzEAId1pvJbIU5vVlCtKvvmAxlnSw3jSkXRRAOJLq3wix/rVojGeX6z
z5n3IJ+czUlTGDjXdLiKFFHFCmcc+M6bURZ2Te93k/vu9qSycX0X5g8BHkZZ81bt
qU0llkAmDpEUbiyifP1aYZnTVW8S1MPHedNSc/9MGvdG1gvPPCX8doibBhRtjp/5
rcxHyU1uNr4MHlzmADWEg655yIjvaSTfyD+jSwtQG8PuifPu4ab5U0NqKiLy5nKN
E1KgFg9Ft0+oE2LGiTEv5zymPWYi5wFw2N8A3hRV8H//LUzcMUwcg6ZLu6tAy8L9
vQnTJG8Bh3HZmc2fQslYqixr6utfL0CMiOc6gdHNuXtaEi8kQQY/wkmElpYzcFzb
3Yk10iNTxRvVB4Nq3lXUFB3FeyZT+LMAyw8cC4FISk0eLAN2A1xKQGdeutGgKCdE
Rji9TfveiyisHOszOE6OdSJDC1XytUN9foptbjxW87woGYCL39DrgKl+x9ksBP1D
CAxI6cKyRcjk/Rf8brZCMxUf/1zI6RDEJAigDseJHCBv+YCDNsMEuIF6sSGje6N4
b+YF5nBedRgr2rZmYBE5Fi8RRGAWj/UcGXtFxjOX6tq4FMrR0XQmgapbIHwdFOTK
99HRbhBuxmN0dR6+xU4Q8IEd8AKYhiDNUnEJmeiLZstwwFX6fJlq27krM/fD9sxj
pLv2iPltyVqrzaBBHLZqlMxYPnqIVGnrtyc18+Ta9zVILpyCI6ezMLwTI+Q1oK4N
npduYr3ZbJNGEVFZftgITo5ii404C08AiHX4iqBJuvcbCDr0bxYQHmtSpmtgs22A
rwRWPcEjdiWmiNZXFUtNRGOq88ahc2B5kWhdQeCH6PCQvo7Z36zhuxxwn+L1HMof
v/veZhkKSKEUAV/iM8e0HZJ6kbF+JNuxJFVMI1g5RT0cmwWa+crHuDTrEJPHNK6+
oIYdx5UGKP8t/DT3Qh6AylnWxEciRBpT2Y4SYcItL0I0gY8wbaeTSvlvDWvK2Hn8
oHIgSsLvTBjG1Bt8D2GN7gFIt1XynMkmjnhXT/1aQYlNT2TCtcBu5sppW7JliN0G
qDgQbtYqgDaaFAve5sVeGhuFZwZsPNPYMx+e366Ov+gaCpZKfQAtKpKdyjzAxgvN
t7RUo5sNq5vRV9qX3V+4Yxdu0lN4ZY6lPxp1ABPeAR4a+4hMMC3QHwvTnNx11JUY
cgVIdIK18rQBDARmCmKySctRDmuNcL1pXzoqPofXGFt9GKrNB77Is7azAXdjoU1J
eO9UDvuUs0g/ZaTqOeRMA5JM+lAs7w5hDNtFy4JVhY4Edpl/svr7ExPuTJOr3TSM
XTN0PKiFHTui4RQi1VQU23pYyuYYcD0zNtcQt612G47SYI5bQgT7H+GQ+4I6gBlq
Qy1u3fjjOjWfoQs/DGfWp35PTTRF31Ihzvrp8EUWoe0xfeCKYV85GhNkcQyUybef
7n9Lu2yf/gJjZmhlNCmXGMN9lQnpRTwQEN369PjLsAWcybVmeBFzTEkcA4vBBtmk
FVZLQjToTI5XvttLnf+ztnL+eHhvAlPKuQ7ocDtyB1Z2TXg3WZjGiMaVVrRHVF5T
lBsxvJqLE+uAtVV7KhrTh0l9lIiBGu7o7OxnYxY7mYjYKvzgrIi5Bs0RZf7ktz9U
sl0ZhkYBG7d4QCZ8HcNAjexq5RgFtglKQVjfw+tNT4fprut3VZgiQKwHFEjyQMkY
SzBFc2Qij7tk8mrTtoZcA45cK/ntutCiaVSJ5gv5GxV2Zr+WDOIVKEaxOUs13rIT
jtvVREx0lktDGEvs9/AbM3Ydj6sKLoD7vwVOVXY1dL9ipMsFCRXSo052FnJdSClJ
4ywGO7Fo57wZZQeyd614a/vdRGn0PLbmkYptAl0YmakKL3xsNzheyaRCt6LNH3YX
FWFdmAu4r6Nx6nVjzmKOZcVWgxvtua1JxXfT7mNmDNMCv9ProXBCDyxEdUczuxpA
Bt0ZaF3nXLhXgTk28o6yf8jID0u2P2JPUFfmral7+Y/kmb6uM+AUy47R2ZimM0ZE
PYcuVZDhWg7YHOvNVZTZYTkiZYOuvaI/cZWZ7IWSGBuXzSMWsu4qf0/qxmWAuUOk
ht5p05gZxA6rHbAGZ0mZ0EWEYWGjuYckVtqKzWW8UGA3kkpTjnfEOjqg0GQgMGcZ
FSzhWG20HjmqruM5KT92FCc5MtoxTIk/PzUuu2GOmW6/6fMeA21APtKt9sYwsXWf
AcqwicO4PMTfTQW6LvzvlqMVvI5CxN7OS1LHwigiLt+m1paa9uGdUUecbMHxzlfq
7BHruTIuWqwMP7kfLJ+T49ZK9SQBL+1kaRnd8bosOBGZ64h0lqkwOluogWDtqE4S
X6NVlz5uk18cJpOKBTABI5t+ql3xIwj/4o6H/kG8hlOYrZcQyl9EjQSCvxGU8D3L
Fl6qy4iocNK8uUEKPqdHdRCQhh7b15vCJ/LmXkxQzUpNsVxfXBa0GQeXi13Eb55H
ICoL0avjBh+p04xKn+y5VPCXAASMCY//6W8D16X3QDmq+nMJoSh63p9EXicgq3za
IBBrTVTaB1VIRuCPETvXxZnTygKSNd7MsSqbZsoT56KABUddFNWE1wtE884RNKrG
iBK7JgrKRNc41cV9cl1rwDWFEwA2JxuZzXlaQ0I1HZ1yG7w8gXhAqV/ysY/y77gQ
v9+z/WYGA8cuGJuaEIx9ttXdZuLnmsihAhCwdOGcTe23Y4BfVBQwGSZEgWjJKbCc
ydp+ihQuANTYv65SR5Em+d/dx1Zll/TdGPDgfahyyEdr8DAAeVII/Q2lcWc8ATaJ
jVcVYKuk+Z4PFXLftYK/W0iZ3Bf2C9lnqPLJSeGyia3HvuILHIizRO901LkHrE1n
8S1enLQg7BkIr1J/B/jUXppsT4cBqsOBh485eDYmvRYN2sGauM1DNj/xYGyhedG3
n4m4f6C2/XoVyCpaYEYywFaT+Y3vRKbU6fS21WQW5s5l0i9pSjCIICZUlzDDflyZ
70VMcQIHR6lNQvpZf2wOgyyimv+dOayKScvofzvE9SkXTk6jpN1oyLbcMZxXq207
HLdaO1SdA8LBKBp5IYE89NSHzM4o0gAqbLvS5j9ww7g4ZK/PjpgyPLuJUs+nJYQ2
GbZHJPAzG5PwcDgd9/L6bTTI2LujSM1+0Lg4pZrMulf7r9tZw6JAeaQurkgc0WmK
MxShR58MV6M3mkJTjadcqHyvarxgIp48HiJebsfncsZAXpA+NNn78u+3Tk9zML3X
boyGxXcT90MuwbvHtDLrejs5fAp0wExcQxP3wSbOeEp5bp9BM/z0/9c2j8SRiKFw
LZ7gR8+tkUWg9VQOPZ3dNUuXWVc+YKymXswrbIAoS8cRhfs+UpagfiG4CE6+GCTj
v/o8UnUYzdRnw4gZ1WGxgMQmDJUpCV8xmioW5ewtLApXo/TdOVOEPUQUBIKmPf2t
8vM0VfABfY8xf2ZVohkqdObdtKjBiwrlikaYelqpSAl23/V1sZDCAQBvlSs4vDqr
Xf3lgJ3GXjkyzgAi2ECa4FdaoLUQRiXZN0aDUchaPX7PdKYJXbBw54SNJ0CKL3yN
6gcLvCdsFXyXHvCUHvcNnRvIXoY4yUsIVRUVS5unadEj/P+6JPV/knySMwVvKeog
ONJ4JRLhY4eZQ2Hi7V6v5G7we0bNg6DAurparr1dcdjk07mzrzWKntGDwikbKR/d
7ZKGbJ3r66DmTEepmaDoLW6FDl2bkcoqAxWXxAF/MapGADOHD77TKmRedlhp6UXm
GHksV3Yqm58tY2jWQpzwli9aWmHE3/M8LR1vT3FZo7gHuPpDMQev6gnkPoPXqIN3
ZR/i5UDU3pTVav9bp8uNrygeYsRLqpvupcQ28wkH7BnL2Ahdj1b/nM4ml9qgXH1j
ytwLUo8OGTTyAaR5/cdbme538gP8XAopwxBiix1fI1UrOYprqHsnwShvOtVf57kt
q7+OD4ewFFlQVR4xRIO0FdRbHe28d6AGIcjyoC0b8HbWnopgE6vVg3OyUcMS5Xh3
+l7eE79ktPoT6IVSBpWds5VRBvJBMUlm5h3bXYtryA7MZH/bjSJV1+TqXeOFt3Um
+UoDsoya6UIlxr4ItLf9PyuSsP1fru6Hcxu6nPSBjaq7EiVl5Yw1G2pxxbe24NkP
So+uBcqK6vfOS6PAcdoD5trYslYcIYNxsAYq1tJdKbr+bpL85D9tEqJiHQy8cQOV
if7R2vZ1Ayas2b0wZFgdGTJ/+2ak+IXLXe24I6K097h8Kia1JPjFWNACSNVJDkf6
DvsTLqLaXpyxgHlVnmv+2TvO/BI5tCstLzqkzXdeqCl1+POJ5GUxh/0Lj58rTuTY
hlvRqNmt9YvGlKaL2LMTPeoD5M+wE/J5wt+A0t6EGMpsQQ8bzwDynYaEr4MYrPQy
ob5XlBkFxfL0sE9T3QK6YlnLFkj3yd/9p0fXZYTG6scIsvwkWVyYdQcjrsGDDRsS
Tsdjrmy1VQIVW2b6OAzsb7BsTZdAmprT/MBJjzCoanQu1SzLluuu2kmCOeXOaCeO
olSW3Q92aDLjUpn8JyJtM5RZgXW+1jdO/LgvSLmTv3hUQtm4OdpITAJHa/SB92Xk
5sh7H8tUOs1PLiV6KGxITSaFGuzhVTaWRuS062ZI26exKzNndSu8G7n57oM0/Tww
ir5IhPGd8+pM2XDxO8h+1TT53zDhvONuqIa1fI9QSIZ6h3bqVSV9URtUllKfMtfO
z2xQYUWtaiMNwheW+LwDVCVDjIqUS62J9xD2DwSwRtyrvlIkBGnKAD6Bia855R1c
rldbXIskJYXrAwbIzSWN1FHuXPqXD3db8urtI5Uv58bZFTWEZ3zCDOfDoK80XLxf
Xd+l/e71aIsiNBIER3lvDXMayfOvLQs7jdhQIrGzv9ywdxe+2evkKn/82CGwKyDe
q6aZsnDM86E35osAl0UxNgapk7FLcM9tW/lrv24uiWUX0bmZLccMOcHfmG/FNsdI
2DeVZvocU1MWvIEssLlwj6//e4RTli+GRTs9NkAyIyAUTFI1MxTgivNkCexLt+DN
3PZITTDsW+S7MFKuzoyZpiUR6jAtTT71cRTwrKIsrRUI6EQV2m9jw/yMYa14eZFs
0qbP83ECqpqnShmeAzJRJttcV+EZOX0vHl4duKWvedF6qU91zg3zErJysIJL3QIe
PoVEK3LOevmAa6g4OshgOxcpv3OAcOK7f2A4jAiOCUXDcFSANQlMAox+SJyp/yK5
32Bti+fSPa9iTVqPtPykvjQxr0tneCpuAmmMPiLkFRnfbXv2lE0cjuSKEN8FBxyl
ZFih7SagYS5sHljmC7khXoUWdfX729qYf0aXzHVx+TBEjM1qP3lLK3IVu9/nkIYR
J14Necn+sKIF3NrYrHBojMmfxUA+7lY2AXFW1ZDeW8NTbBvWWo6J81XwbXJX3WEc
nRrQjmmQvvEdzLFyKggsBEg/FzW/W8Fa+gcZFIfqgwavSRHmuuF3k3aUwqKB4y9l
nPlt8fbXuogUxpYb54U4raf78EKZ1KfDDvF/Wvg171Bz2fSEl3Z+9h3kyQJvzXa4
bW0CUxpaTPAk2rfrY/gbkxvK4tsqWxFNVkOKYZ/Ja4f5Oe2Sh3ABcEOUqIhnuolB
bOmiwagTC9vO51V1wD75l41aq88kAIt5xJbPSw6EuXLbCDPqAgGmHkNnRcBE8FW6
CCubleyNQd0eIgQ7vlf50amlLghTscnssv5UWLDF8qW4ryx/JRanuNtiBcXLcNXM
i9VjkTKSvTOSAU00gUN14+KmCafrRhFICrWiCqFjUOA1T7FVQ48ye241TFxUXoxK
1FkwXTFuDfNJIthKtVVHf6gJf6HUTNudI15+IjOwVhKn8sCVHfUN6Ulcf9D8S1R4
s8BthoK+9y9NUmh60D3YofcCGGVo/v8qyoVdqxC0Qo1ooBE7NjtHjyT1JXuseWVk
OpUQ9sxygtcpazDCzvmcIr7jbWV4TJCcvJpIRb1oUx2uhOFFaeHuGo+lNVZa5oS/
uH//5y9lGNR398H1cS2nlI8iFYR+5piq7ajFPVBpC2mH27/5nHawyewa/9BLNUeN
j4kwPNT1EaRqZHI+YTVoUEMEjrOd80J3dFiJ2YaOHKymDwJBoNOmuAFZkzEXL8SW
EJTWXXcRCyX1BqSuWBbabu0iPDvr4R5kJesnJfSqL3ixmw+RMkwvVllQaSOnPT3H
TfWzXkmaMq0LOk0u8XWS33S1EUfT+eMJz/UAONkwlqRyJcDBR1sSpH9H1D4rJ71P
8s8wibjAB7lxSRyocsyxPIjty/WGGP7/i2QhDJoK20bCNph8fvSRZoVU+VQfmvhh
Zr3aefRGkga2iow9FBRcPflOU31Jy+LSVB+rRy6TjoV1wUVPJfwiqzKEhjQOGHIG
uMlwFXavJzB/WtheGvQgr0Tp7EbdwL6sBsrcl46wSW4r4UOyxdk+ZcDqJVNkuhCC
TIOPV/Mqi5r31tQnU6IbIErZOpobx+VrhUNi4YUDJA/I0rVEOeoER3UHnBev812I
U41W4yUeAxYWVo12DtXKuk+vPIlcV64kXqFWrSYet95cp/4T06Dfq10k8yKIPpnN
BKdp8u62U0OjhJZi15YbSUnS6iH9NHpfncQXo7l8Q5KlPMKMAJKx7QgC+2nN+VmT
XOkFs7366Mrqp/YYJgJnzapS9mMEI8/AwAvL5GwAphy3r4pIUB/RZVY6fLb5xHFb
myMoVb7pS6TUWEaRNrp/pgZSOV14WInfd6XWn4q354uK1bH3eJ2IdTFqYBl06ad7
IETJ6g7m1XivBPG16RfHYgQbAkxW5Wwuq2ll/U6MBHv5EuTTJ5No7dwQnkxc5XmD
N97z5Ag6OiiHn6eQ06yeP/ESKqSYVdnJZCBGXEX8rm9YkkYCZ5bThCfZpYwWhluW
uC46bM75Ss+J+v/twYQAEuWEC5Kh8j/a/MeUBW9MDZgKkH9gguTrAe/XBXA15Fcg
DZBgRu+esF2OnoT40AFn2XsS1SnnJ/wRWz/z02XPJJjHzvccgo28951a3g0/Nu7C
N2KQ9ocLxvMZcrJQTs/5by5wJoZXo2WCq7GQ2s2TIute1zjaaXcmRn/YmA71WyNB
YxTI5pNb1J6XVRwMJNndr0lQ88lR+o127CvUzs62ShcAndoS5Tm0Q+hbdTnVyJMJ
+FsC2khpnfrHgYaNM0cKU1cpcAnzNkTVFTInZ6C/i4iGYY09bjpBXeFP/jQsuIYp
R2B5h4twsdaajXWmW399wlj1QbCD8Jb/3EQZCXhh5c+DaP3Q47ue+7hXf79lVipi
jSENUzpC1en8eNnLT9KLjbka5+7ZR0/9u5Ua0aTKje0n8TBpy5Rf2vIsmztxkEce
Yty43pM3zKrv0AKt76u6fRiXPT3kO+/PnrEBGhJYVBtSzhP9S9wNAJ0wZvvIRSrF
4thou7Xxb16odPTLJ2Jb2Ucb58U90pFjbzDsOvrl0RpsmcFZfpvWRknUdAuvQRrQ
99L/da2Y9rxvYHonAxYxYDJyYietHaijk9+rFTLv8y01MR4h5HeCnPU9b38eNDE+
LHJQ5RNpMOneZ9cUCLYdYEAamOYVz8u9WXjqh37xR8WgBao3S2L+zq+wb4Ai7QrC
bmmwGfKeCTIwZB7lzixA91wO7k2TPYW48Z/awUD+myjWcBi5XalZlzDOba2L6d6h
1bYJnwknjb31ka47499Pj5ybALGIqYrpPm47Q2x7re3Zryq/nu2hjkQSyZ2m+nFU
m98hs2pgJeAH4vC/f+KdhsvQ7hU21pemHsX59dvJvaunKz9D7am3kcxgVupYyipW
YUARLfYz2WhYEliq8ZttNxHGKtjeKwWx4xyCObf8xSmdWvIL6LSDsYAUM82cr0Zh
m5RPPkiN23zJcreiv96y/wK8KQ+Mqhb1pUuvMoabAGuaMD4uUwRWcgeLZQ7Da4IA
mtrahyfJ64da7f/G6VBM9SeiJEWYecqHFyGLAmg0ec6SsBI2w6u4LbAaA+ByqkMQ
N0/wb37MwP6uEJYUNz1Se6cjDAE4O/1OxA6NUCixwRco8jKj4ILP1tn1Gx2tYjCT
Ku/UOj3UxFZpdYZudtnTqTWem1RMz7/+9fVH+aJXwyUDqM8P+FyfSUnzbQrxJOLJ
LGimUe1HctDDGO4XHyJvWdA2ip4W1DyxzFAaeQ9OyT8lhHnNVt5xHK3w4J/bvjDA
evosRkB//fouYLtfbo4mMDHLBl2NekTlE6MVVRKlBAgu6naw7TdgCnAlGSOfWx71
mJ48bFjNgFD0lhx54uem4H1LjHXEb0XScjwmztJp6s3VmQBzXx4JrplPwdB4p79A
bk8yACC/LXv5cg0FDvUvJc5wiBdmjlgrFNB2WC7pxl+6QOfjqw8qA7s50eSF4OkP
e4bBOOiw87LQBcA3cZuERyJREgZ3cuupxYymB7KsUN4hL00yOLhicjcUkHmlJoaZ
Iq+/MR0iwuJCewPZLzqB7HqDTdBaWkBq5rBhqDoUO5P1z+kYfshuN0VYIi4+wB2i
XAMJ+c0YVInu61j6F+qEs5G8M4R5kx2kGqj75EYMJ32sSwwLpBy6+6yIQx0EXTK1
CjpejOVhNFAvHW25P3ws+2FO+78WidwkghPmjq52GfskjYEuQaPqZJMLtO2RUjPi
ksYdNj+xfWulKDeg7KGMqANT1+ax4fWdgOQ7CSd0DIaYfffDmdGje7PiINKGPIen
cvFB1K/3mAqYwKAEfvWd6EU7TOQjq2yHG5LjSW4Lj/vjQUtMIaX/1TEsMNDOCqqc
OEAf0f+BaDxZjTTX1ie+gHWi3zypN0plsbyraedovs+/wG4biEjPEmWuyCSo+x+l
u2UxMBAMBodoHIaXlgULMV2mlwOZPkoZtQi67PJEVCXCOymvYRgzIqRbbPVALFZ4
MFOguFIeRhmzrf3MR/r12h9h7Ro/3hGZTCnm3wr7ma7lnnFVn7Q1RoZyumtWWzFW
I4lH+Q6aHtBPxKjmrrCk2zWvG5dIv/RCXLRV0RAgWFx5VmhowuO2y9vu/KxOAnza
ny6loloyDiF2SFvYufanUl/rAHw+dqakOV6gJPtsjXjg0n07+HRUCm7AWcAoExJ3
PdJWmYjjXuwv4/M14VyE3KCjWRnlKLwjPtAZ8IajU5+oGBG89BoSSDnz0sWh43It
6bR2oP4RdvdvXkVAu9TNT0bVRvEVQy0HoVz4MnPK8xZRUckEXxwxVqWT7hlEhPRt
LEYwGTYwvnCNV1EuZE/QPdRgVX3AdEySeJ+Oyu2xuKk/91+fE3EJWPAyzGJwIzr8
sc6Wq622v7OZJPrdE0i0XN/uWqwo5iR41rr9fcrnzQUy6NIwv2NQ3NHGe9Xdh0OO
FUO0V7fSK/OtbwDBjM/0XomyOrJDc9OOqv5vVuRkilKHhIwc7c3CeYn/WvGUi9mM
TYrGJnprQAy5SfpeAlaV63Pv5kmKMjbfsVn7GAU9Qo4CIV7bur2tChqrXIUET6Vj
81Prq0/rHOPZjUIlsIMjRUfKXdSc/Jk1ZCFP74xVFU338/YZ8JrdTPdAYIPenF/H
wjWQyBqKs/vN+WZD76iTv4BWX31WNU83Xv50kGN5LBb4nzulW9wyD17TL98PjKTS
Qd2P3ZQpulklZWjKBij5cefTzDIocm7usC21I98yYnKAWqgs/A92N4MOSBrETsRi
tiA+x261uPI/BevUPposk28h/B99y7+IsvXSY235YGDs2suHa5c56OK/LeuZUdOp
ah/um+jR7HiWXDaltlm3koZyDRJmvJOnPh4szo0OysaigS7XnfDZ1BF9ZOasEMrg
oik0aR5QV0JLq3Yc/7VQZFgPX8iHFVZQhC/QA2CF4PhcLERtWQGfJZtQPN28Wmqm
/LaumYSj/ngX+UYA1i9nSSSWIOCx6ucXFu01IKP+hZ5SGbMI4NrkaGb3PEKtQsvz
9NG1qYZfx7PCFO0sIrcPpRRuJwMn1HSnSOEI2sK20cW19DfgttG5BtDsZGIz/mq5
Re7T8hUZpQlEm7RJH8QGyhsenHVK7wIx4vM9aKrSiJcao2AdH2hgsyZ4B9JR/jfO
K4pi8w9530za3VkpYrqvUbZZwDIzX6yvPFnzqspS6D4Nbh0UvIrf0HeeFx82VCHQ
lH5Rn45QfGw9cf0GorHKrNHNGSG8awyms1/grTmXm1xPYRAWDMMtj3OKzjtjLiCp
ao0rx/XO4Uc62q3T+eWeuzWpYDHnqEdSwZV52+ygU8tcTAQZQ+U/lzQRx6bW5xAB
BjF1I2bvth7+Q5lXxGfBxi1ZBO5F5yMdDTF01MxyMiqOLoF4XrbkyMOxksR9CR9R
JbsQAQDB7Ua8JgS5mM0QhaD34cW0pdxADgkxsdhRbeWjYRn/Bm1MfN0WHO6xwBAO
diHsXeKQ2Y8CN+fuHNfhwJANQOEvEgCIf8mDONiTz27OXvOgtEQRfeAT1xoV5aEX
HQzQtP510gDABxRdItLowEZcAJdQ/Qk2aS53IF4qrZ1YjrFpWg7pRJM2cAkfN5U9
fSRRr04FCOT+39ow+BNbkB6Jxk6csFwEjBUYf9w/R4KA6K0ifQJDaze88fcnA09n
B2AlHVgDXaYQR1f7B3AoAp7yqpqGLfpM+mNQOE6FOXkb/inwMylF4eCZO7ZQOfQt
s12kch+yWMJ8qnAxnhNdDGz35mwx5EDvVwmHeO8ocs7p+MFakoDqc8OLO2j/j+gk
xaeNjgj3xrDBTMTgSJCn9rtot7VV3LIcul934s226t9r/dhS9fK0G7HQy5bonTzM
Xl43lQP+gMb07G6f+2lGe3x7t0naTGqWf0xi6FPE3aJWktA/Pj2z+u8goN/pevY5
k/ghCvjNWqjf5Xi2Bv0/Kn3+eOfMKc5Y5B5PEZ/GB8Tz8x2n1n/8Pf51AxwG3Fvn
nGA17QSpLy0ln59J2yb33lbWX0kbjLezxZ/wpaH6ccbsULR5xrc365oOicxpla9w
2I1CgmiLgFmny/4GX4K6pmAVfumGLwGJVUdEBJK2BTQ7+CM5NbkZTit0ThTk3otA
/YjFrx4WpuRvte9wTU7f+wnhk8T3jSh0rmeACLRC8K5r9Zeq/eao9QhCu7DtR5rB
63UodIWZ+COgCAQuvIay2l52xDj+he/19Hp2BgmFbNAYeop99NKzSFZrtAzmAUU7
UzRrK7KsIXyymboxUhU8GrrzmpvK/Ke0fnyLbI0cLNLAwJZnQNUOXnG3MLu0ynlC
nQ5MJfpSUd1zf+lQRIVW9Onua8uw28mInkCliP68+6Da5ek2va6FPxJkT73PzeGp
A7xziXnv/klIr7e7T+G+YelwmBavPqVsVFOt+3qsMT747fwHbN0M6AHoHFzQO+Ly
32brBwCkGWczRiI2EWk/DEgL1ehCIhju+++UxqFK8AXLuFYMRDM+gtZ3R+B2CmNB
XhxCtOs3ew7vH1ktBu7AMnwaVQwvz70D5L8Ofod9b40C7GBqurCc4msgxOXAvJiT
uFjQ7x1XIwgPREALVRLE76CpagRkjIR5gMMuRZjpJxAuP55KlrVw/oOB2jZfda5b
FoTkcWlOTO7MGuYHdK11uLrI/uij3tKQioqgtMn1qjgrcEQAAQQskKmG6MfJysQj
a7qy8uu2/Sy9N7B58R/3BN13KwDJLWp4ryVjuIHqqmyvFhPM/nzd2ZN89WABWZPo
6o+F4eTcwOImd8HJdzgnmfmMMNwVawumKfO2EFjoT340cXYOlzT2ds2KgTZeIQ/w
hVxDUTJKqqAZh89PO6F0NaEXml09PruN1j4jwdXLjSGflT8sQh+O9usS1r6RGDw2
wQDiPMHaO2+lY6T+/PSKXMmsOvHVfX+sW/bXEHY1mVKy8/uQJX/0+l900b2ohW+5
Nx+ewGf2H2IdXXrhTIpbfLH4uQHxVYnteDyfyl9QvVHhFJopJSYDrX1UDhLVWegD
NmCjxRi+N5MlxXFaTb8cGt2yki757msVUNai+MmH0TxHmpyHBIdOsvNCSOoRT7af
3a/i05L6UG2Fnx4tTeBN+2w1mO3nc27HlvohNwjCSpjgg3KwrfsBc8XgDBxgklKN
FPJZJVfM5bb93SBgIF3c4xLcI6nKsRQFVRmCbs5pMrqiKwSA2ZyO9Hc831RS5FtC
LvGqO+EKfOrK1NNw9IMJW4vQYaBJNW8qjL+ocns/2Go7fbB7lLjvg8rl1e4LWrwW
WH6KfgJjqValcVZ4kEUIwgXAHQ2ABpN4WIl6HO+u0SIgRKoGLbi7vg6t1X1VuapA
tGMXIytY0hyvvhQaLy9yiRrgM3ddRtk8vo1o1OYOY8E0Ez3auRbQgigyy9BWF1br
ERjvGaqTEfxSVoO0kmECrZsL3hq/BpZr+23YWHW//ptlfvfrKrEbf+8y1rN8Q5al
LAPVL3/yV75b01oedGzUs8VDUHIs37mfnKGsQAfCLeCoKxi3Q/S9vRhVy7t1jGBK
bBUkcgKrC4yI+5NSet7VXl7MBFNBYSB94GCOYYxrD9H1CIvQqddNXx4M/NOSZOIv
sps0Ilw85qQb4vybeMx4WB49/1D2ehFB3mC0ib0HEsFQd++DudSNmX6nfzvFH+qW
ZNEPO2jRUD+z0C66TSsiXLqHRS/kvjXoH9dKU7Pyk8UuSc9M3zFJs2YCEmlu3wUZ
MZqs9jLCxIJyBKSMV79+J6aC2Xc6Hct60CIb4fGTa3ksebTvqHgcseDHsefX1LaS
3Po3h8rSxSPUio+eQvnEYBgdyZe+G9aJhEXxGXnP0Vyu0EKy6jPNTkFNRpeOooCg
eaNsq1hXAyXgfqAhKChLZFh9f8W2eYzfhyvBi5D2X7T6qQt4gEPxp8C0w+mRtg6g
3Gr5NDEcCjCzbc7xsQ9JhlDGimBIkqMHDe957dAN+XF5e5rhusou4KlHb3myuWsp
Hz6EiCpjD2bgPqbbPcIIdkR9XA3FmomIThoFJX3bTqz8gUSIx94NJvjwuDGE970V
Wl2tXQqVXvLiJPnQXzJqd42SPt3bhOY8M8kIgy1gTRA5lywmWouSRLlrHzGMSBE4
gmUImmNODDrMJnjCYT+8m+YYMR2+enwnwDPM94OveVqBqJoGYLwckeCEYEJJ/ke/
fBuq2AHzBTl8ew5VBOAlDEXWL0d+fq2sG1oCV1aaSPt+PLnCDDkcGO/1b3Lb8x/K
GJ1bJ6FBMYqDJVegvpBva6spg886K9yw8pdijtd08jonMBFu8x4ml29UQB+O4L7V
nn8xCgNGZEVYyyR1qUJo4GU7XA0I0KhFT3+XOiNOSiKS/FBMbF7h+RxQDdD1LEj8
YvZShy/02KOa1eEl25iBzy0DImGWN4CJMV2JNjxFUSxt/gYa94jqRVq4z+TF5/fe
aZsaJ5f5VmFocHXMT/ifV+ROzmFvy+z01v3tDS8lJfXhyCveSJJj40Bnx+jkqnqM
y8KlMC+sMQUXRINt5hqr9pczkp/9l2YlC3lu/BL+e8MYwRvUnvVkeiy1OzS611dl
wufPH0X2gLG72Iylj2GVN1FvxqfY6O9L9rTWhSZOIjeKJ1nC8rdpxVxDAyEvQMVO
jwdlil2tFXvE3ySrPpHtYpgbuAwpYjNmGQEg9W0RSj4DnioYAYPx6KZCbS22+owj
ugKdkdoMcxVGbE6y0ksE8ePPoX4JlSuZ534s625u7OrB8HmiylKn6BNOCJsSRdFm
+etq7rEAWx+CzxWNL57LBk23/mcrRqFyS0DqljsbBi8MxgoS5qGdRfB+0wcXwfAB
9nRTkXBfDX1v0acIOETqgFwhZ7UucMk/FBpq6W3uxyWIX5n+CLZP1g1vf/7BrqTl
qfI9qcwsDf23NZaWPX7EuD4xWPXQVPkYxKDa5OBqGrA8dcrWIaEpgFV/dApRHfPw
Bp+7EtBqACRYiULcZVh0s5hWoWQhdUQ6iaqYAYAzQFKObvytS+7luxA1RsNXdrDZ
KrbuV9H0p93wJl/VQLU0iG/Nq77HuITIl4KD71qyGaTPQ2Fj5H5sWzCCK0ofrtJr
rfT6IDv51Kf7wTjGktI2y/s0eWOHwsHY7xww0e647CaEnEJ2RqumJ2U8rmh3S0iA
/YHlTkHlLvfNEpm6cC0MzclLskJYXpJqQwZuRQypnAG22VLRvrAHqEUYSGGUQXsQ
z20ieeZHwpPNmy3SioIkgDmc3DTPzhe50QKvW4Uv4iscVjlkqe+9KrqJMeJaALFH
oKQm+WHi7OJidS7nC9nTbpPmYGJnq+y8Gpd/T8hFAjnzxBfFa9cGVMgWwW07rMMt
YIfAum1fvRnUhHvaKrIAInHzRdyL89bxeYBg5bva+ob5HfnTYgv28DXYWSYhpxNK
EIIuqFCpxSoNHblvRZ/GLp9kmX5dkY0c6afa5oTrr8euliGYFnMNW41XPIxUiqvj
dleCTLLP4yiAKVllR/0V1XXArMZfQszJcDWxggNOJNQcaDNkojlQF8WSCDW3s/jF
Qgz0eIBx6n2M64XRw7SKmaHO0MQzQ0TBl44HPxd/Zq9MBwFeYVuGKanwdXN3Pcz1
Fsazf7Vtevg966GYtn7NNuBwAuonPY2zdIsDnezUA1mUZl4XGDKLW1CFcTdm41Yt
+OBiGJX+2VPfRfCayngoDoJtZAC2Y2UQW8utwnbHYUehX56tKdbCqYHfOyhqXTu4
Wr0kysBklS25L7fZD8CPgTg0ZYJhP+2o9VlRWtxfXvLPWgbm5pB+rg570+KkKDBs
fi2E0OB8Hb0IYjHM8OaxFV536Bj7l6eC3fV3F6gunYE9st3SF8tOP8gAZEq5M2aL
1Bygvi88KXPR/fFLJs8Kmx3gpdZvAhy75QG/8lK0IanHTYmZeyEQ0l9Vt2NJsIKE
pJYIPAgGRN92ir4N9u9av+n4l/e3CaZQMrXaQyyT2laM4CkuzjoGEG+LTiOpPKb3
kE+vToqEdu0MLXOCNjpzYS2q3CQqfZD28jexpZ21XKG2kGl+nYvNSKm14PrOZlxP
RRC444dcIzAx3SZE0FrwxYhXRZC5wDHeGUffvLFSQN8TBaTl5mVBbPpXeb7L/mnV
NUXHw3+qDUThz4Ljgx1txCogFvL08+jVKC787tJiEJLFzx46zb8T9TLYC0hNFesL
DZo8S3xOBU0zvag9H7aKzmPvMM993uIsPxVW9UG/AsLz2Gluo5/XiGSKsAkAsD4r
/wc6gfS+DoRGL5Q/ngldy408Vmo4sj5RMuna4pQ2ix9ftAYVR5WDCCyxR+reziau
qiDy29dPh+6U4joDEvGuf3eVbY7i+TkbQ2UEw2WW3j0OT4765ABVRCGIF0w4iZcQ
/uTJaBLBCnETqIWRYagLHQ/WACHFN4jqvBqUHDiA3zbtQQAtVQrBVHo2L/4U405Z
sPNCob7gVy7br78QdzLkNObtHqgmfTA1WV94Y8R1yDmZ9cq4SthGS3EMQ7ks7lOq
7560pevg2DC4FBhLAHFlDogyV2nGMwd/CA0MO7t/asnioVfJLcas3nUi2APBlg+E
TdLVwwkNwGgSdSGwC8xJTElfbON57IMSSOH4RFyoIwTIGlAnq81BstPGMFddFxVh
ekZumjSiG+osHs/KqGTBMZN26oupiUkoVQfBTnI+LdnMn+MIo9vH5uCioj/oLnez
E/GmnpURZ0vV3QXO9KFfy5jK+Sbv6I46WaGhqZbbBrOK0qyInKfvTYCb63JPdgop
Ki8uCyTC2LF60DPp9lELPcHJoFl84OT93+DOkrZ+VuBqjcYnF1j67ZGlfNteQU+J
eS44+2B7CiK5Yizf3CNJIE402HSSiEaSIKlxQGPRBt1jiVOFc37E5lPLZkxpNppH
EPPru/9XnjjK0G2fsvRVAilyl6K3cJqg4XKiFpYST/EBRLC9G8s9zOcnT7tQpkjJ
YdL716i3WOvOuh4ZKOlEzInzKYYrd+E06h4yDbBpwS8UMh+MaqPlnmLm//YA+1t2
NZZjma2FdCNCcRJKqQOPD2TMDq3HJe8C6EqUUMxripLKA9T+z2iOypSH7mw84qaf
OlZKGmtmdrTKgAAWaYNFJOKjmR/IqksLfDQD/0i66ViIbIJfLMp1Fx+FGjqFPRIN
6eTcjy+GelOja3lnpGyfl5Lv+4DYH4+z9nfZEmc/BNTvDtBWOhp83kbOUwJcSEb1
l070XxmWpGX7T/Gc8pmBr6HpnImtef162kHbpdKSW8xigh0YPCJOuT+QaR7B+WPH
PGaXoq4NFAKpPv3YecGO8Effd9DiEzfw9UAn6qyBIa7Nnw8U4MxRWU1VciF2Qg1G
8xv3duJbSM2pvH5fWiuzN62lSBW2brC5c02QCDZwnIbVCQHpmr1pQL6Gd5F4/pRO
M9GTnPmVm8GE6ala7GkindFD8vWi1jTLm84Dz/EopqD3tCjG+1GDEWys1TykrAuh
cyn0HUY4jqZWn4Q46flkgCQBLnX2uDIwmOuJ/rHMrybzXSgErtVWWtjA8++vp0c9
4RiEJMA/bi1ebtfw6Owd6WIfholu969GhEMfZp8bnu3pc+8hJpjOcouBoW98Bh/j
ovF0VsJ0HqdqUeso5NVtqcCr2Wxhnojtii/mUhlikecvg20NJhzU3RFestoBYblm
bw79XtrhEbAdfE4JPW0xGucdICyJ7CLKH7AIzAi5/TXDE6z6apXpFzFL+fWPCdHQ
01KRFPdLBpZdk/2FVs3FdP/yTfwCitArLeYqo/STnDygz54tzLvzbuWj1IhxNYNt
Pc0pc9zYahNS3zlzy2gU8ejMOzyF6XansdakEiVQDwUTQjQhdsx6lGAMzcg3k+//
V0DKMSQHAjg8TneJJ7U/KcAT/PDOqHxAI6Ik85FrH7/dFITLKdnOWQen3ApnU+pi
yAxPJ4jDKv2/Rt2O5S6z/dTziWoAkzdPNnXxf9ikLaIgZa0lNieZJUmOFQUPMjP6
EE6tZVQuonfU9mWcM5BlDB/g7DayDAUKNDZwGKxKrKT8moUs+6gzCid8kUl6kE4f
fpcWlPdaG2/M/YfePIl8U31upLzclsBNFO0M6IhS3xvD2RI9TV5E9/bkgYvd2hYp
/vq8ImJ+WmNfNtf9IUBZmAG7YRR0R/X/i0DsPPcGFUxLMedryflZoNlvOL1D7w8R
cmyoihhLpp0nqhQUAQIbYa8JPLaqwwwqXWGd3UqslYcRNR0Q3OEFuptymDY813bR
k5AhnMt9ay5GsOnyHGcJmzAQbyHQf3Y6IZTlsWqtLB1kzhFq9vxSJAMTzkRwD4DO
z0YtVFufTbzJjwL/HGHKj8oi4o2ZRGRKMgP+boPpLgMzZ4qi6+Y6fKL3AJ5jrezx
Gu5FPGozGiWAIpYOsacdJtZjYI5D+yBTLw2rKGLEjfm6FMQwyFP77aDdC5haVyPb
heYlQ8IkX0SqQu8ARzrSN03wE5pwTyQC5KP/xutPws0c8kY0muighDwcMVcCbLRW
cYHSpilPfA8aQF4s2etot842m/0RpML3aDlkW+btbFgGYUJ+lxqzX1ltZgnSD7V+
S7KQK9MIxwhDi5vXKwWFyrDnlyyzw2X0xtv9EEAWoXSLzwS2ZD0nEDgGmPQT+nP9
NFYekIAJLRuwwauaR20iWoIM0XLA6nv2kZ8Qc0Nd0s1ug7CFuZzDvwjvXsZPnMqy
J/bDkLOJ9qk7ZI0sjAEsJ8qHwnYhwWLyvETb0nOVXIDBKv9gPSo3N95jsdubDXBZ
62be4p9sKLc89z4GRHGhz8jSfi1wyf+tE84I17Rq1Q3UnSAy8O/LVdxVsfosBp0+
GNgWAcY316aGtxT3sUyrhNdXIfMUILazQBZakCLLssmpx0/l7jFEDIZSVhRsfd0Q
WvLiN4riBXRo6Pz/Lw0UqSgAISqsHhhr6AXjgLp94dAHZd4swLlMCnikJOw+3+3v
5k9Xc86EerozS8NBLpcRQeE8X4QJX+y28IGxsAY1fBe0l6vO8Y//vMM6cnuS9T1F
mH0gCjxUGZWknXCz62qQET7PEyHU5XE5rNtbk0IlTLY3QEXg9iyCedskY1J3wraw
XhhizjEwB2gtPwozzUdKI2MUETPQjxMq7KunvMO9XbF7YqESBgnMe0nxPEULGzhi
Vj90HMfxn7UZ3HavTMxULYPQu5HgGCNQWQMVrA1QbfsA7txVENiPbtiZkdtGhjMa
MLfhUhgIVFqdsdc4u1EEcF/QUByeUO7FgYMc3Eniff5DOiz+mTDM8BhHYJaKpFml
UlRwvNiVXLCTTesfGH77c++iM9AXS2rJT+ltPKkgvf++LSMzUEJhQKmdrPmi9kt7
0VXLh0tqbiKsosLs9IMDaXI6fdKVlibMIqhrWH1wSBgZIXjzeOLlnxNT/Q0EKdOj
Iqw/soFK4RjhxsxPVefyG7/hEoPY4DLAsPFzcf1YHNDou4NiK36v7ZhNJHfyA6F+
fzrUe2HjH/P6Q/vAJS9rKUWp/Yej6Rgd/tSCSsrJ0ikuuR9omZOPtOgoPH0vGe3h
51lTZH0heDX2gt+1frT1s30s/Ux3xUtFpqE0IimJeYlsA+bMf2u/11S22JSocVjF
jQg/TWf448BZ5f6NeYWIBdwa/q6kfJhx8MDgA2nGBv6rWUpzzHC3mJJSpyaAaJmx
NRBjvvGxasfIjgRZ9bW9zjuof80Yc+W3BugxYhBfRsAANFJyRUPxvpJ/BObHrFP+
QxbfnozqZgOZNCkhbYqXC/iQpVK5+wk4IBAHI2iQcFWb9dQjjEXGmI5t2L/lLYEO
piJjGm6f/OtA3u+rJU/5ZbFgAWEd0EBLCgdRwxDxDbmYBmnA9fCVXvuo1vBNNIY7
0UrA94OH4DmGzklgcjgw33SR3LYNGlqwl1J4pfb4IUIh3W0daemCS+p92GHkUY/W
avn9qT39JL6DpSS239Irf1KFg5zXIN/UKeoF0wov675luh+7HnuNaszA1Y9mXYhc
d3Jbqep/fUrMQl/wS3GKbdUfwmSU4J3FORz/Hit0dqnhb2/l960pEuTpa+1dg03u
f46TpdwFea3ud85aR7i27H5DRZmlKUq8wkO+QB1nDk5xbyPkYeT5BA7Y51J0OvtZ
UjjfqAqqh2i5j5d2juFpFdFlp9Ncmr5bVGqyPW5mJnrmKlsse4sYGKZ1Ip7Tmtgk
ZocY8FhrBzPCbMLBviWMfohF5W+UvhO9gBN/RORI4SpxEjxzPiur+6+EYdCPDLWK
2H242zF3eYRa3Ckv76wrkmMfVpQSPGoG7CbfDOrpNV9YsA0UheLIPi9jNH01Y4Gy
DdMM6UE3yi+hVj09hZnGRAvyPNG4MFOFv34QIwUk/EB9780HWI9VmS4Qtg6UUUW5
TJpjjE7QWYRxLXXa8J+9URci15SNtwEfka76vdHSVopTR8trxpN2KMaQP8hL8sxO
QxAZYTqrwZytmAPVuFu0AeCDgBtJGuwYlE/0+hxxkIuJCZ/yC0+YJT/k0W6UJs1X
wYaYaAKernzyhHrx1zqIlYuJuHZm2C8N3VpGvD67Fr052a0C7iPyvMu3qizVUEJG
Yh7Ga0QKgxBccsqQgbxDGBP7jibfAFhwZGzqdLFhx9iMrXB64gWINBrRtpilY7fT
+N0leExQQMFz/ZxTn+a36asrCgTm6RX8+F+2it1glTy9oWAaucYh5C3BT2530jAb
Mge7GKjBeiyP52fvUM1gXqEAIl5gY7Prr0x6Mge8Nh35cWOrUzbr+jOcdcTzz03J
Yv6hnFLrgfFKQuiY4gAeUXp7WrTFhyEGTFwjIAY/bPIZYa0/wcUUx0q7HOEUipMB
Uz6ExI7YUhtWGuEYXHcP7kEvKTHh1m3s5HH5oogxNtD7tOVcTSl0j4gj0dCet/yT
U3jIp+r/X0j6WufnAPNqPBBu1cFs+B+hlX9E7Cl1gj6z7edOZ0zSV2cK6GZc+vv8
0C03oBOZYTPUKQAAHoV6k7cWjqKQ01zrRIWOVP/6ZCm8ZSjbTGbwr93La+bYyY9l
ydOu7CwLX6Sb4a365Xxy51B812OrcqNB+dtqDu1brs4wstSrQFIfmGuTeM2J0ns7
CIZcDqM4tKGAcRy7B1jv/lCYrV7OumSXXflsJu3y8STr0CMw/txMxQoTeGEmT+nz
95viryt+HLeoMxZV7R6k4VWtPnBRZyva6jpzWnvcMOYy/CARkdSmsn3A7WDe1KAe
GtCX93oVaIecZqw232jfm2ZB2tqRJVSev+3U+5936B60uphGi/HRGzrUX2pwtNVQ
bqRxss5bT8HnHeNhEycXfsQNqjLP8y9EOCZPujYuaUm4O+bQyEKGwXRrO+MXTwoH
ysav1pj72TKOsPEk7KZ1tEa5E+aGCwJLPpace3T5TUI0Sp2uXs0Jm9rZZD4BmDQN
z7vWBhQnTNNT7SXOnUfMf2XC01R0oo9Li5czzrizuOGB/1+6D7VOpAf79BqCF3zT
T9augBHWhleeJpcWh0h/hGBIUxAwkFqni+7iUtS6FwJT4RLTIFVjc1RigDqMwPcn
YXBCaL4ffiDoL5NnvWxMDuWynLgPBIYZz0vVQK4DOzXbLmf561lA8FHT6uXLyWlx
27o+mG6Py/69Ay7fPjH3WwIi+BebVN1I1AcPQ3wRG5tODwbWGQAxj3GZUbcp7pTJ
aGvTdD+3IX883OjcQ4WJ/io/4QPiZEWXdE26tPr4+png+axTiayI2UtuBKseUam1
8wOiwsTMIi2MjiNAHWHAncwmIc9iIrkvDIw5I949GFUbiz9VGi2+D5996h+mTVMc
7NFK+GPuFhj+9RyFFyA5zmKawtT91S3RrL/TnZE7sP6ysrqmPlY07GZUMCJmXeOV
6m9A9XhjGJKboYVrJT9ewlxfBSlT6ANPFjPM5jjn0G6yQCUge8pPLsgssec6bPA0
EwlyHZGGovICza4rB6P30nO1zi+7hizC8hh5ydsxeHgDOQVlTOHo3BD784W/SI3Y
xmpbLKIkFWsy87kjwK0hfazta6Qlu3zXVOIB5usqS6pexibcZnQTHOmsdSYIKkwW
3o2Sx/5INGjs6KIKpNAWRzy1K45uQekWKDYUrLsuvlPEkJz9lvQnDH3NNYnSv/fE
w2fjFIyw8KPagsx1+9xW4y3dQ/oCIL3DXMHPaob9jLHq4L/ZNNZtYrO9+93F0pzm
pSnO8VccJsrRoOhqwm4Qhygmj+d+egCXEAD5W3qqH+MCxvjbtU3iJ6hIPLehWibm
sxyY6d41I8wlCRX974DbvmZlpRNNZCyR7oeu/um3idTSBAz/1OmMogjS2godyzfv
suiDopTF9tWOcMraWtUkRM0L5lSh7ZgaNCX8o0ctgDDIiRk3j1rB2eoZjOcEHDCW
WLGcG4ywh97uFI3yKzJTq48P/i+Y4LUbbpcmLj6YLyMr8IEyF6AbbNZpXcj3OFPD
SBBfiVUfwnr4+nJHSBP7UOhLKiqidz6U3j43iyn7xhuLUNtmtI+lYh4nNFSsHb8C
GXOgcAc66dKviXpDxJwRkWKg9VPToNyAXLbYE26tcq8ebc4NDpxo1A5qeiG2ctNI
UqtalVJy1Nc54iC5q9z36OELeeJyI5vmFineNYmFCFFw+Pk8QEHTOfcrp7PQI3fV
fVpoQG0Mhn2Qd6jbzvoce9eNwSGhvGoLAhIIDJEDmz3Kpk/YDvgyySEJLO24m6wJ
+QF+LnZD10dDIwm3dggtzOKMTlHEC+3Jc/P8oudaq1oq/QE5c8F3NNuMd5ANC+Yg
I+9aN3KhxJnkM43JfIRdpey9OqKc1gPOMEln/k790cGu4rYKgr7bfwxH+NQSax5Z
ei5mb1WSOsH4WYhHNrYgbEtcm2bClKMv+1uBDbjUZD5ggOcFSNcAzuz2T5Uxb6Rv
c6EenanGYvxywCuTNVXAb6BobbiDLkWyG/q5E+JZk/BnHXuKQH/Ykrl7AFH6UauR
H4zedIdv0b1CRZQh3v9U+CzhOhuMaU8UotAcgoZyfLF1YIvYYJk2+Y3rBAkJXtLY
Yhk3w4hnb2rlc7AEF7qmQ89gVCP/7DQFVISj6LnTWKYznF0UQKRTIelVNUWzSuso
qbCx18ujoFeR8BSuaF0q/IOmbYUl3J45ip8f1c7ToIrjV2R/3nRn0xzSDSw63LGX
/+ske2B9jQOLg789vuioNME5w9P8SOGjh9vRDDvilsOkMklNywe5sWAaVbsHP/mK
m4wTxQg1JqZG6GUEgEGFXCSkQDLMVKoyVBDnc+UnGCmd2X7B+xQjF2STQLx7U6qm
u2m/oiYwZKpJN+MEpB7CWYKcoyibuCiFEsfjR6Qf7tq9ouJ5ZaM7m8sHHuXG2f1H
jcPZ7I+SSbHjzwA64u9uxHEEeqx29CJYUYJr5ZjJj7cSIq3c1a53nIoop3muwvvF
kVcLOhYH+vzHNNQSGc/sByFx/qX6jGc1Uen+SIKk1vtxiTkTzpYERFcQ2aKJSJeB
tnVErkLZatdtvC01Yl/Nu2HsNrnDep2q7CLuxM4e6fmLdPB0oem92hTVOie21GRp
4PGZ7l4wjni/GqfjR234r+JFF6MMI4In2xaSxCrStqLWoG8mZcEHPeNp8GEv2S6t
Pm/ky+aHXjDjQ3Y77rVb6OnuNDIu2tE5YqqFOoGsUoT3Uu6+YVUFAIqXpa5dINK5
VOiOWQc6YROIma4RMbCRusvNHbuULuLhY8pmAWB2U/LJm4wdqRiKvXGiiuQ+1S4z
/T4Aq5zYQdHSqwxsuWSU5KMi0qkrwsJrQhQx/1BEKso1AoXqztbn2nL0rW58xyRr
V2vASRtj0rXFvwws5D5URy2GqK2rU5QwFVRHyEqIaIvS9HOiA+Fpiy/cJvwauexL
udv7tas7i3zxNoYnoSlXawqnE/FZhCkQuD9S+Ulxrcsni+qbegjNQTob6jPBkA4V
ibL6YYBH8qeMno8FFgjfQud1b2K52QmF1BCS/Zul3YbX+WQDlq7wI8JUZJa4885d
sSfJn1RUj0A92rKnC6/r2l5fq80j7cMZbkpgpRh/RRMibUQN/9wcKJAuxgJuX37v
hWtsdlPtEku43SV5LBy1fLlRUGJaFNuhUr+CyCr08Q3gBDgbkDdMBtGiLJABOUe8
5Y4XKuIcRh8ibSj2G5kCgoBVcqHbjCOMyaTU2WibqTtSBy1vmqqYJKJfN4pGaqhC
LbP5Hv7NXs7BVhW5kezdwldMPJ4kbOtIHrf7yDPCseNFgN/iDXBVY1lZ4GytHtRw
69j67rrX6S6tcxpmwWgXXyjrlijGd85hLO1f6ksPT+LEV0JO7PAPTqKH5tiMRkCk
evbmUs8Fjhek6PqIwrnMFnxflg19BX6p8ixM94rfzIA5DgJs0b/l20yS5b6ALRLy
f1RUai5n2L6/T7BnpD8237ifs51r40tXeFP4JDc/h4Mt+EmrxUmm+xcV7bQf4hZc
YSD7eEc9yEIQCgdEex/kXXfnWlEa8c4UN9ZJE7kBg1+jewnKCxDHGRoGhxikInSm
C/aArSFQl+qYvKLH1TvGvomtme9eQj2Yr9HzRZ0OfoQVK0KKEBka4IqRKpB4+2vq
fTHbm4zhuYeSLM2sb8MVUZD655IAHYovfdRUOXP6XzOwJzq5z7Tmm5IDRJQjKlmy
B05kys8Y3F8S4xYoY/bI5uy6X5Nv+QqvvKrgMPiMk6F+n8eFb7JjidriNU25ccrt
bfI22UDFJSR2vPISI6ZNCo4ENGF3CWrHoKB4dLtJix3uRvzpF/lZKurtdGVqtMn8
7Ay15TqPN0ARBobncrF9gnqOdQCtxT9NrXj1kcGDc6RcJNnoBO3L/8SL0kCclqOW
kzC87eU0PR14QqVFmDpMOddQbRsXWn7y3hL8ZTiRe+YvdkyWsSETupzXPC9RKYV/
RnFbtVIOhF0Y25CcL1mSDVj9E0PK+nyq5RpNJN0uwfWnw9ShbLEflKFmB5Uqdm71
lsge7b+PkJXdRuzm+u4oDZztywMOEC4loI4y5wR/0XvFMF4VdO0chHOxnZjFMsfE
6VD2gbNV2HsK3ejGg6IW2gy1WiIuWVWUOKpadgJ7GGqKZh4eUFiZot01Esu1gz5z
knOxymWFQjbiH0JGakCJ5+wfijFC3C5R6i//hfp+fO1COrI3k0dxVTno9iMiEhn9
o2rGRSQgX8GFPiTvrllNK/lsGewVnVnbQ+ePyKkzq7mweubgXnc2U7XtxoUMrB7u
VhuRqOVbINxYJT+ipGInidkAnpSN/5JZj2IInQbLr2EpF8YeQSXus79Zeu6gx1gp
DSf8eyCwEfdaBywbOUJMGYhVxO5/Vb7AWBEh6BzBXhfA/2wrW7o2wfllDPJYG+dn
9cTZohp/hjIdV+0R8GIcFyG5q/cSFzJ6jRMxs8HUmqKFITuWJGOPy/BnUbkQrPwy
Ows/s3kDVC+H52fr9sjXo/KtOeBpM6YKyZAMDnBvdH9eqcsOu8ctoHc1cISaC4Ks
rvn81F7V4iYMGHzV8PK3eLjx6ouZVe1Ep5G+/ShjNE2Yaaz036en9B9K0V6NtMva
haGfPWoG2d2CCLd90Rde0VNzQMiw4k13Kx9ds/ImTW/zPACtGq9Zmqkqdm2+jKWJ
brEbx734m0pdS2OYr6rfGmfqZ8AG4E0oxLjPbePeNOfAG+5h6RQB65AG4ArOoUw0
VC4TJ3FtTBm6uZ9lBdZrwumkYx5+yMAvwUeuKsYsF9PHF74Sg+emIULRy8iCZ2ZN
8Du6I0ygcSdpA1OWMGXs0UdWQTEER/Yc+QIZxR8kurQmfzLwaLaHqxmni0yroA/l
sT4Yi9eDONcnw7QUPqQEiWGhsN/ZGppV+FzaojrWXgWggVl+MQOnk42G6UtDRooo
CXSC0UhVuT79t96Z3lhFtdySEmIXz7wSK9J3pM8fo7Ytk7Et//kt9Z8nN5Y7dvAJ
u26suSvqVF/aFTesF/3gTJuXkO2dykS1FqP0U6YO/8bYmvTZXp01jYfjWVl1CWwW
74qJYMQ3wSUu+bAk3/q59COJdN8118CQ8HhvzNu2X9MypXHCW5yjjlAVdkbFXRmP
QBT+9YdbukBIMv2MQVx+8iuX6rdKzusjq3qKD0B136cgSYYAoXlLPvvwZWLmvLvd
P4aRI8T1mfuCc9YjLuvWQXMmFhvI8JMbJWl47UfKz2yDuCqNQRotMH+OUod/2TYX
IcwnzKIujWOrKV+MdQGPLuZed5TC3Ul8PPPrqEwuQS83cRMs+ObkxxNSI5P4fil4
u8Aj6WGin8IZiuFmMhlVffir6ftuUW0FsEND/DW93xdoC8zzpEzma/vJe8hpcbiU
o5hFIx+zcPgV4SAjiJCUc06wqnTUzpOhuU6UGnpXGTCKP5O43Fd8edK3E+98C5V6
k8ck3Fxx8lFCw+LrwQ2Z1S4Uykua5nXyl8L+wyJRUGwcEUuU1MrxPPravD+k59vp
QaJpMNNgG9j5yR3RXVzMpjUCM9dg3hP3Q/mWpw8Je75wU1YQnLqq9CbNi9kH2zaL
XE00Wh0wsTslfz/YOw7WEWZg16jiy6rJLegq5M07bkd9ijLDvi/C+lEMYsYw0DCQ
yQB+cdvvg+7A15f/Df+/cEcbhMZCG7eQMIFli/T1JQbUaSs08MDhMi63Y9NJh4Hv
i6x0vWWyzX4akdkLqy/aNGPd6qbAsAZpy+arHU4lT0TuapxLfVbGR1o8DsLWVCXH
AnsEEfCf8wwrpE8bMzHT2Rv0QuhDmufjYvKhkvPrYq5m/pCX/49NV9yEBfvu/ScE
JosIsrbUF+UENq4uIe7XeAYz+p8TcHcHHks57XW2KuDQL2mduSsfaovp1AAJ1IRa
FRMOvsB6dZ0MXqfVg4EjXQN6ojOkdjIYG7zXsRZ+ExwRuT6PDPX6n0G1NOuWrGz9
gNsKVvjhklF449L+EBUdKUmSIezXbQOhl3mqqcXbBBqT2dHUnH+dJDNQ63IHaRCd
q7JQ5yU/nTk6jMoHbisjVEDnVIcnYCvC/HMZ/5zNJjvbUlduIDbBYB8+cDq9JPdg
7a+H017YGuE37Q2av6N3QzzEaGVmsq7EqQUvzp44rre10A9EW5Gc5pLQP4rmFceM
5wL1KYjOI7X17cs/5qNtA0k/O4f43juHy6ipNwEaolmtUkmBOM6GxHUh5YpuRmg1
oxP3o3fLP7vUgvabAnlFnOC7Px7pHwR+naKlNCr/Ez56tsu9PZlsZeeIrq6SqoOV
GhvNIc3eG6i+DgyK7Y7xN8euwNaNmHUCWqJreGD3Jp5sE/Evo3lpOHh3avcL7o5h
VxOh+SYyEpqneKYD4aOyOAFYB+vYuRpQeIAIpjt6ziiEDeK3JdFHC3HIet/ePQE2
0eJ13p3YIvUPhx8DFhO/i8oER60UBt4eVk1vQuJnQz1zffvPLdfYvwiIYpE2QoF4
F1X3fijTM9CtC/rH/3erK5elEyJZCIysqHOhTot2jU+LHqNGgCyTo358ouTSgZ6j
u9yXSbmK5QcEqIDjlrMABjz5EhMa0XBvoOOQr1+M0tg+4qh8agWRa3HyzlSM72Mk
0oSIhRGmFDnsHkHWa+w390sDhCQNZissIKoioIWSzIa5WJbb4oxvSgFTy5cJqJdH
igp+Q6ZmO0/XkdsNSBGZ0X6w6YZKuvF5ZeXpsgTCDchgLn5qds9DIPQHQbqsvasL
APE9ijOBiJHEBBhzYVDmGMJb02HM8h3XxjMDFLvW+RbHOnhxJ5Rx+U8MK1GPVpNk
UWKWfktOPe4WEFaYozdpntZT/+8cAhLKfTkQVNGRkuq5vBQhe7+BxK4uMrDlQcuA
lgT05EGlKIMtE8Pvj/cfkS/UtzTupCNwSqomNYCqetw3pUK4HmQGItDQGXZiMC8A
6z/857Kj+hWQOxgHFZ7A8nkjfdMWQ5z7aMAiqXBf8As4b4GC/yLRY3ULkZECYRwh
+pNzuoKFmrVOEGxZ13MIbd9cv3tokA/+E91DylWw6I+TkrIQp5CGszFXnXhDpwlf
qIzDuThbjMMg4w0FO2u3sg3a2UOOeY3BWIoHbcE2aRV4XHTb44yqhDQgXt4cOj6u
kluNOQ7uehembrrZk1iygDryfAUBESCW0vBw2HzdNIz3SZb+cEY59klDSy2Abugw
4TABNlYlIg2kx7H92XFukyRLjPT1NqQzIHuGBDvSyp0cuJEvKDY8p/Joopgp3/jt
D825sHioE529eETjffw7tJMkTx+DWXUqvfUs3nw4MH9zLd30Oob4yQZwyUgGj5GO
EybMEA6EmeIAf777uCywQUXa3CNs6HCJ04dK7izBZ/E45S29UnPKQtFPc02XdLmd
EjfmC0hch2Jj5581d+FI+/naJV/f6dOyV2WvDulrJ12VV/oueHxZNLmJagzGVUl6
gOD9+nPKoy1ABQ3rBijFqqxdNBg/hlQb4tBTHd7wtmrbCSI3IOz+IO51GYMNnVqe
bFFWpWVrkV5CDMHoiQRCzQ8dAezZxL5auMAqxO3pvK1XoM8Sdl/ruckHCMb4hgqj
IaNeuAW2eHsBvB+Auy09eCkXREuxOEQo0PPB80FrSMIczmBbFaiS2Ke6P7du001p
Cha/Ur1aYfU7X1hLwyYFabBy2IH9NTu7K0BFKNrqTkvYQoGjuHfMATN0j6zBXUjB
sCqzUAUGSwDaJDvUthEp+nADqdvMgleDVozS8qYZ3O83CLqY9U5oZpjdf6lEXJqT
got+9j2F8Id99DjgHyIXPGlFLysZxA9KNqQUnjKP/eAjEZO4VWoFAFTmtVHuV7Yx
X/mT+B11LUBNnYurl0aVDRcbqCHO85zGS97+E0quvRnxP6PFaV5yiwaQdJRVQIaK
guyLyMgJXlL9ootVmUMa/V35aFSGjVRdaw9aGGSTQOryRe8ywdWzf3P61gHKk/WR
VYcwd8u4jljTSa3RjYm6K5C/LyClaMHk80bcyawgmpUFQjloI++I/DubB3plCvK/
O5VFEJW0rtFMySxRIUeOIr9eWrMjQscm5E4ooyCaixXO2USVdCPQCtm1ZpQmlI5c
/y/NHtvrnS0UF0Gq1Tboh7xAOdOCCbczQWjgF/iklt7LJobIRcBHFkwhpKdrwwBr
QW/oQwOul+Y10OXwWOD4HEQ1ATEPveQJHeAy39xcN8tkj/M1hMKZysutgrItu+ir
1SWKKgzd9EpHraMFBxyQDbdgM3/sPtey1qzvbUw0Kg1iPmyMVgY2zL0qqa/pYQYn
W/vvVl8oTUYIvMKY8eP5V0Y1bJoweKkX3UfDj+ZFTSZaAVF2gtjaiOONnYppSnLF
La+tMyNeJlBQO337hQw14aPazWZ4tIDu3Im5gbMBkhfDL9Fz6wMXGK4S97M5bhpa
BXX9CbVqWcGy9SP4iVG05UEFTSboRNqKXhZvKhEVJ5edThWh8snmr4BabMKB8um9
Kk3kvlbJgQUbiU7NVjDePvP0U6sa8ogMLHRBB7vCnSdBG49MSrhJMWqHYmC3Y2bP
vr3r/VfCmLftmuDowvCdYQXLCwFXAVqgTnQ0+57PCr0ipVp86BX7yHaJxb0fHK2r
8mJpIWjme+MnBJXj08y7yENf4aqFgXzndUrWROs+HZ2/dXOOXIbqoQ4uZlb0e6iG
AyY0DQMHXIWjB1lAmyRp0D4dXvZNEqLDVErkTrLhP15IC5fcDhKdBK5L3HMhY064
/hstrp2i5eyLM8ZdUAGo0AbTuRC4lXIIeGuJi8LuI33XfIzBDaZB7jkdFcLzLvZa
sYvHwaQ8vpFc2BWJeLBVB182LYPOQg+JSd64TwgWdhZZM0UnazTGpUyMu3jbtegT
GwR30KQ8y8KmJws5YOtVTMWLbkzb/sVPZBaAF06d8G3KOi/g5qWQ6Zwt0Bhd8ZRp
iEKb2fHkLf7FqPX7nFfA4APGJg5ha+I2RwIyCMr6TErwEvuX6otQTgC3tzo8B+gu
3qCBBzzoKpixncQvQs5q/Iw8V6dkwVXq0bLY8StPAX6XoZfLz8df//n+czyTnLtf
35x+6mDEmVPy68hMUC6X5CBXJponLwneWiOql7BJIspGNl+n75Z3LoZ/I6WYibae
qjFoUcZbIBMnC9XyWg6/cCd8SeFKQmpSrpcMb2HptraCzxzdC8Q/ltRyiBSU68V4
Js6J19scejnf5j/00CdjtPjjSFOvDA0piLuV2OJMooUcfgPS8B9kzB9vCQrpcEQd
pYFXIZcqIV0OLM2xPj0QE0Cod5D0FlS3dtsiRhKQgucKqlkW9glssNAex7XuazcA
fjYa9IevwPanw6FHQ/Dgt3MYsGfvPUHBr9AVT5IbGxT8Odo85wdhKwzUhvKsFFTg
OlSavVUfiU3LInZeRaYrw2Z1bHixo8BKEMNzzSejZugJusqB9LPwJsjiXoLA2djy
qMSEWOwI9XG6hPuEfFq7+lON1MJ5RYlpY1nButq8rG1OC+2C3HUaB9ZA6IAGdORv
/D1EFA45iesByFo6mFs2fP0nlMHSQ5/P+LnaFxvrqFubfhEUTE3KWCfrSSjhjLfj
e1j2c2kWjO8Pv0fKNr44Tjtulx88RRGpqe230vb8wwFg9y1Wz+bsqg9TTcyHixtd
gEHv6PF25rG+Y9AffFxor7bQKcwFVddVfLyScOniLczayYkIZ1Pw4G6d4QQHeQl9
3mU88rc0+p3wfDLAF7x18RaHp1vqCE7EjuLRJQb44QxbEC/VpSazMTcnWE6okMQi
trxQqYL9BLG5NBfdRtYJUtlxTa9nMBdWTg+go2g7mkmtmkxVqFt1a+rvW9x/1UxR
Uvt26HGmHNDyCW//pfau+uEPmbtboIKB5hShD7j/MgMIf6q4E97e2x514WQCLxKO
iGeIzpD/ECt2U7eJ7mxVG7X4IFHAxaXB+pn0+9+unXAjD3G3rVRCiJ/tKjFG6pHf
VQmB0o8yLCQQjNh3i9CzCFwbFsYLYOnKon0+aSAD4e+BfPw31DmKCpQpfUTPGCY1
DsgAnUGQwaCQd7gBuyidfNsQeUTK3ICOWmZFwKwsRtRdfC9SWzO0e6FZtlxcoNkf
ll77MCW71MT+DADiImKYafyNAnROZfbzOuPizaXOzCGyjv8RfBOVK8mhGtn3YtkW
FU67t9tr3ITeIC38JzjmbCh7ogN4GozpU1+FD+HvvEjtE7rphO9wwQ7YLaySIbfc
1iogEO/fRjFCnTUY+/IJONiQOWe0R5651b3JmQXWm3RJSEjs56kz/gPuoLNv1ysa
frK165XQVU9a3OAd1pOEs2Di5VY3WtD7sL5V3rjmLDEegRxWuiHMnobRsef+3PnF
gVGjPCLNkaR707ohQXP/RbDb+RxkFSVkr2zxpifNUGLpCjSTexRvfZgjG3Am8DnA
cN9QLdI2QzOjpxD27GstRamuGAIHTBAWEydCVY4h5Kd63dqLinz1eSuXs7FiDX0k
qDb6t2NSMMME+AjRYQYJJTk6D48+q3c7Vr2G6aYP2C+NVTmQAMD5KL2wbx0q4wv3
c4bnLPr0D6b0+cCmbEzzMNemKBxxiaDW4NaQj9ROExIs7DpBvF+UJPz4bRy07MHy
p8SWrauP3kz4Qjxyg+V5Xg8VPelo+hd8Vufhzp/3xDF/sdBmFfNrPQal7XVXRZh1
qOWwgrdjbzunu48AEDR8TBjRJOcpMqXnL0I6J8D2jXMUFyAHpfS3GVcYUMczJDxN
h6TTDoULa6HFZ5kOCFLItDPLHrNGcIteic1SKAMVXkDEva9syTsTu+IIo8jWrxb4
h8FVDmDdBwMOlxpLTAp604Tbb+eYY8JOtHNAl3spaKm1ZPtfOw2AHfNpNX7VLoJM
RTLlUPubwxxe0KCT+veXaazVYQftSfvLdW8rLsNJEgxC+Idrt3vOjLEFKJoGMnSJ
HDxjZqqUBfZEW7giTBB533Z7ehX2LiLsfsRcP1imMlLXWzcJQz5e9qM7NMDpmcHD
I+hkmlApsjUP+Lmk9tWfPDTln/eHnPmopTZz+1glpmcbhsPpmPVGgCchjuGDa0yZ
lEJi5RpUlhoUGRCd0Kgvan2R8YwWlH8N9YzS7XP7RM0iZAkackvwilVD37lcFhMp
g2nvw6Kb3MBgYJCkXRWhkIuXFhTUHYrKacGOmOzKtOM/hOA31hGufTkhFR4CeB3/
w8c3RgMAvflibHl/Jrpt7PVkkKFZZOI93uYLk1b8fylecAGmnIH5W0i5MkzS/fcu
CsR/ILRiEn0Wc3ygPeGqmIWRqiRcZNejyNd9i+BDYjlpXT3qJa84iOzS3oh1j4rm
NRrKZm1cS5oZILNqaSr7vKkDy+vrpJ95KbED89RBz4eGlFgNA0DeFSeHJl6+/z0f
Y5/Z2DSvayzEf8RYz6/10m1AyKhdZ5CvpE6xfcWUfEEk/GWCHtvpnrAgt9FYtI/N
BBHVGxPMI+mS3dU8MLOWgae3D/9Xm/QtubN9++V2IaUCSGm4R+C8uefP8d87ITR6
O8QLLTICS56CNSNZeQ4IcUHkbhgU6RLU4LUQARTDk4j3QMPSSZ3ytAEgrbvEpe+F
DrBhlroSsTfRKN3bNd9asNf1IQ0EFW+SPvXEkyZncb2zONjtdM+QREt8i2ZriY6O
4IIAY/DhRCYIziw6n4Z3lOpyDQkLNlhjY8n8tOSYZnju/3rQ4iU3AykwJO281Ehd
HMWYxFOcO8qO87f8xVdOsP6a8ouL9fJkUZ14EibAg/w69B3lSepV/XP4G8rvNa4c
VCGIo6ZZ7arJ4P8dtsWfrKx2FE5kJrr0iAumlLk4A2ajgOxKwfniArYn+KRL/k3n
1s5srOQce8tV23Lt++LI4eoVxy1qTpMQWpteNN317ECL87oLd6zbqQcEHiYQPkjr
XrWROu93SedG7IEnA/4ZNd/pE1rFDGpOAQXnEBXEx65vfKopKlt9gGzv/9VHt2tD
8gssTd3gLhEnP7rvoyPqBhohWOvhrBMz99/WQRl+VzMCZD9cCyEkRRp552TMeFxK
8/i1xj6UScvpgXam5uw92uUbtOl87rG0Pp9lw9yJ9wC2NF7P18sG7jXCHPWXGdwq
zHY/zYuGRvnETyQT941CLtDJ8gCIJsra8wu6hKxtZwpVkhUbaCrGVHVm+OQ9krJm
E1Wg05PhIxNkQeT2f0xA3RfZH2WHNV8m7RNBmdUTIVXEeqeuQTXHOgJsWzKLLvA4
XHeFikI7EoCmPwTZDIrt1pq/EeRvl5G4TBRLABpc8F22FKWXTUjRksX12XdW7omG
O33H9XUn0FpEhrQln5tgY2zz4HvMKdRp4yhFqOtCMCYAOjWx2GKsuxmN9+Gnh8TQ
aOGUDPqMTMtTqOL1FgWKs6GtEaKr/dOjCjfNbiS817hSzv8u7lilYeybuZVNgACT
nbI7iRJoqRxjJuwzqYN63pP4DjpcCm5+4H0kDyzSolWgm/06XynuWsjMlnqSmHtM
9kJSznRuwc+pQYkRcs6ep3x7rx1ge2d7iM40KUvutGhXuF6xGuIHYuyXZUJoMQLD
h2zkDbkwkobTvG+lTme9DJ0wIvDIphWJzHjc1H78GDwt5LYWEPpSHManaRLcjQzG
PBuB9Ghgjfb9voXDv3ndkO6zIBQ4w1TMn2gfWaOKQzz4jiYQsaAiHgFJdyMG5q4G
DSa2rXOS6jY5A8cuvtyuufCoTooEY+dAkXsNltPzj2JiZGzlVbT8EoU0mqg0D7C0
DEcI59PwdyvJX6Vx8hhnI/dmFGCQPVpeY+EWMvLI9unePVd9nhdABQwgbvOWA9Vq
ybkCEn22VJloV+SGctcE4JG7nKiYJp1Abh1JuJKsgUqUG5EJXtRU8Axsh2zHUhDC
zdbPdr55br4g4lDSKBE/90nfU0vQolU8m+rKHUmgKbEJxZD6i55Dy25s16QVdahK
Rn+aOfIYp8q5ZeKgQeqdz31GtYJvGW48NcwG665LT1PohgdEJvhTkMv0fAevGKO6
EGBa5NDERdisPaRJDiSZqb5ZwSpt/9XCTI4G65VtLzxcW5Yqc8HXwPpY/hIWgW0j
kANpq+Pt94/P0W3lqF9m4phZnDVgBI4AdFL5MxFJvwuocTZsauOALuZc+Pp9xgCH
5AFdOu8GNdEeA2fddjsgiJkrI/NF4xawocQgA9dtzzeAZgzw6iBImCk4vKXlwOMO
MKVI9VqxB2STstBMs0zP8f/rG/GoaYy51vWWRjkp8dCY14LC+Fkbist5u/g68dO1
3Uv2KhZCUQVYHcQiWXa88CmbFQGRZKJVHesTFgRusC23q6iVHsdrEgc5pAOdzkR+
rXmfXwv03DBO/6k+Aki4eIkggwog3d3hdP5C8ucM0dxmU1qD7gVflX4bjabDvSV+
9v7TMDc9TG6wUug0BqOtx9DUybQhqlvJzUZcGs0B5oxsv+keF0iJiwETJ7y6fwA8
LVnKmsj7RnKc82A+8q1BBy1N2zQnAwztAzkbxCDTfGs14YGdRT+Qj5t5lPTFyMQx
unRn5ZOL77rE1l+cVFKYNLiGXuG+dDM3XO9+iHVDGDEextJYRBP/R19oMuPLEWdP
NqtUi0tl5KD1IjqsfMbQs69aXOyJosJgFdS/L5LDrEJRGbpvl2jhtYPhM774LaRb
je9SJ25g992KNX8PsuywhWCikxYg9h2VdrBIDr1VAWCnFi2IaCDJrH7Z6p1sVyEK
/90ZH3TsGiPuQkLL7ofJbxDlMl13uzuV7B94MQ0eTiO/6sk9x8+wM2LYAQLZ7tcN
xnTmWBNxNJPSsOlcsFfmTK+J3GIRanUY1aPjssLC8CJ59xmaBVIeobKLRtvxNdpN
x7sIbTBBVGEwW/aeK7TD8bPM9zom/IZtlN8EvTqi86+7AGWSVF9WjhPiyk0zeqhs
U8N8tK9Ktp5vfPeOPBgH7p0OX4UP6I4sKuVUKEnZ/a4mDT8suGXy9sgTB4YOflzY
UosQjBt3SpikdBPzfQARwFK7MkzZJf9PA9f57HfhBJ+5vNIJFWbrl2dQ6VtQv4eG
JlkdKc6ckncwsAuHeMmhbYG+0ULQ2MZeXcPmHmL5TXDGYbHUu3NIEsy8TZzud0Jh
/85eH+w8gLWsFYU0JP4KX9+R5Is/N0hzXAIXox54kK/Oqvy6/TaVE0sIY18cvKRp
aURgM52ICPenwvbmmTN0leq2pxxcCtqWR4lvlJgUBA+rrry8ceVcM5kiqLZdQ5iF
jdhMOymoJknVEOb+JYAV9LRQ1xFwMBoChnhmQqpl4P0mPU2MZ0Fwnfsr3kwhBSpg
IfhnDdoNtpMCinn0/u5noDzF4bvSK1R4/amSb37tmhkc1AedGwqZRDksyQXDs4PU
Om8MUm526AqhFgJ6vMMQyoYitP4AhYf2Vs4gU7jVLUngWB/YKz/Xpmfu3NUuI8DQ
Yd51EDBs3f+W0CoZSz5rhst5YUrAa8jMl0ZX0CVJeUJsjAFBxqG8neHnEj0DEYS1
YQzjCiWiimd0eHuyhsuRkPIwGBeUQXsKIOABCZpcPTO+NKlcQGuPGd+U63fCveks
9GrIfX+lKfzIDQOSuE1ShRRbEXx5nIWu3ddkt0ZKKyX2uNL/mSg4CR7UppVwWWkF
8hwF8m0qoSwa+1bj3xX2VXLt5K+Eyr9DbPe/DyTdzChAs1H+GQkX1zy5I1dcBUd7
iTEHBzYamHHGa+dKkVJkKQKSBRczSh1wahi1a4r5mILnJdehPJhQLO34ExWP+1mm
eewybeVYBr4PP08sxHa4DWcMZGj2u+0MkZjO6hIVAQi6nNdDguix4SBZmISDn1q5
D09ahi/Gb0t3K+KhWvac+mOU8yDQfYFu05j0gep6IVoym/Kp4GFAdyTm6utmUkQD
U3/pummgUHYVQ53KUrPXNguzIvx06ehI/PaDte6wd5CtgtAaw1kci6G7hAbVQY/a
7QgA/BFQ5KlZ4IHRp25UX/qlaWWoylDxpA0Rx25XuszT5Lr21ZsmlLrF9/pGgm2R
BZHbefPwgzrEsjrNOutr2hm7ayvfTHXbPoGs+AjnXowe15KDTLtLpYhzhph0zUMa
lbgLLgrCLgtRPQ4xsaC9QI54cYwbF9IWYULQxVgQoZ/cMJGKkuw/I4gE0KXp2Li1
NzZTcu7vplXrGa3ACTn1CoIZDEVsE9/MZnRYGd2fUqRNIWA/lzGcxq68mmy5xR7F
lzqejZxruLs78e8e+du/AVuU00VxX4vbREiSKDxoncqdudJ+/N2XSwgG9PnyOW7s
2f4KzXnrKYlNbNZCVEJDVjFUIpiFXkJvfmZFkJz2ZjgjxLHpLYGt3lEVY5Qo+gxy
+JYQYJffpOwhFb6Y7NzEDlw10VM10YYF1mNgkMDw5EwiBaDXdAy/EDKx/XU7cguP
BlbRTXME8rCjsWWzgBUK2MTRKPfJZepBeD7Wbx1H9sxUaOgF+MUZnS2ReW6vwtob
aOnZso2pLZsFdCa0QGhEzBXPgvOPtvp7gJXPL4SQ0XLPONs4B3Py3IpErqxT6yU4
3xjc1PzfE8c/6VZW/lM4OY2EH2qJvPOc+WWu+wdJjTqpcHj/OIjtmU13nIvbFSP3
wtzExLo1Q3kYQBB0AgWQHSbbqm0ESdKDj/FUQA3vNrBWEwgtqcKftS7tgb/Adun7
nlxqfBYyVK9rMwMDfVxtclrAf80xOd6A1BwK6OmG5daVGjEY4cKXfPC//3v2ska7
nYm4k1cZpqx70555iZEMtE9PGQ1vQ4mppzBTeizkPWtI0GaiwDnIH+hWi2G19H7R
iG6ybnX1VnnHUHj+o6nVlswcR4UKkBBzqHiDHJMTrT1UAZQbJyKRv93qFTy5w7pK
zX6VJCZNkqbQMwxK6h69xoi74bJyjynsFTRi229McxGdN/Urwo3SYqJDYuibNeH/
hpYRNfPQMEkdFPA+Irs8Xox6ShRYfTkx8eBt3VmQuZei1Vr2KHaJugHoHvDM1O46
uIaDojY823DqdiRMmvwgs1u3dF/Bgtk+DQnPYFFdpgBWrz8MfAXFgD7SbSLyqZ3X
NKwIRNOwVeziuUl83Aev38zjGUpM3mkTr/F9ERjNF1Arih4dceHGSHXQXdMUsIDp
m9MX1UgAEH2kpYUEc5H6MdmBVZIpsMr0+5QMAGA1BfEicipBDZJ6pZPaKht+gYph
HtKR+bll3yYXvbJ4F0XM9bJzqkXi0L2abVeVXUjTvnEpw/fT7+9xhFQST0J07cwK
T6d7jRkEKq57RCkVkbtwtOFlXBEVftPUonKOQWAYehT8q1u4dRkUb4PRY2rE/6RG
67NHScOfZhajxtYve1VE7DtGVzKnsuukDYHT/G7ZqPgLpRpltsvF6AwfkiecE/yf
xu9nS+pvs8tN5B/HjbmihFRUmZNqtohPZvHSsNUsRuGeF30FZtPFx0s4A63HO5tz
dWv97rHFY7WyKHdhVPKJpmDs4S8QuGnJk8ycDQQlylXSq9y6cIW924OQ2a0/AM2w
LkjWFs/1gPl745r275aHwm0xO7ogDgo9d9Qs2Zh7j74NYpeUnu1ZiP/gqzd8eWzr
ixvVjCzcqltvvvrZkxyf3+tffxfIJLH7S3vXRKMNk1yQl+YUkgiC8eXuf8jPk7K3
KkyidVkS4flTL1nJEH44fbSysyHCssw2IkHqyKSM9f4b6TC/Pc0O+OaJKb3s12Q+
MC/y5BJuuYuBozEO1EuwRnruI7JW7LZbodi5EsbRJ1QO8i6Gr8hENgeHpHU9iC96
TvVqAJ6wdtkLJ0N1y+26fB9MHTcHchkaiTq0kEnGimMglEivuMkajtp0ZJfS40fq
Jj3tRD9Yk8T59eqg48JT1LpDeC2CoVoCeaH7VmZisPalxC7LB5MeZSilYAPBV6Q/
h/DSK2+dphOtgFFUkJKvXNODD6ZfrxHL7QdiZ1jlvSNgs0RlZiwvxFNfB12iRrdm
ee6Xzrxel8EOeIavvQEfM1SXp28HyLUq3If3gCKlcPNg+/hSD9/4MXaiDBrYVK85
vllj1EkMO1GoJIki9JvZDUD8zomXipVNDv9Le2U0VB69XNgAPxyKEZ+y5CoCKDwz
5HP7JxPA3ZlsvTKqF39trGWR7eOfpYw4enbDzyGQ4arOpdp+PFFNF+IeV4slq51F
VCR+0OyU90eSyM8415m2i0ATT9Q+TOiCAIJ6Rv36VzR/R5yly0b93O1ae7bp7cYx
ZocWOyvskU6AS8yz500VNtt+9kXS8FkCVgdavx9dkY9vwjCFSyPnF4ezp2Jn3NlF
yMKbMNgBaPJcXKQxou7VJvPezbOEjDAzi32vBLMM9gNqvJDmanhdCcnmeAPa+EoQ
J2cUJfAYiLiYvGAySyTuBfJyUhDjQN0EwaMOGEZTbjwjThlzesmIloFGd5lQElei
Ivwd3irtYjDiq2O/2zFTXvB7XTj7Vt/eW6+wJSxSMC1/04H67OhaU4smgIHVOaQq
xpnfZK3jDmDjhct0HfB3YyW956/LohniAkrBVl0fQyOB329M8oeankSCYSYHB46z
qn9rW1aErwz4WdpWTuJToxmDBTtvsw9ZSEQIqWgfUrsCFL2AXou/6mVUkcWj8Gfg
+0VtDGg0Vhu76NKLRhMAx3I8eI4Qz1pg2yxyBW3dGgL0B+4ZdOui+kg0EgTh7Qpl
VnSwOwi8ZObXOd4yMUWu3gXfcyey7LZTWx5T5dAGlOd/jFXTJkULgt8l4ACJ3Y6X
crJ1h4c7dIhzONSjh+vYNRtqkkqNtUdqvwz7Vbsl+bcWFqA8CdQ2jPBfg09GFVsQ
a1y+p+yt2ZRcwEzfTHZufipo6uVF3EibVaxea+bOzgyOITKO7QLCNoq/NYVQCm6N
l6VnTF5dxI6FUb9lPVf3VoW3lRGnGjzHZcxWNec5z27c8riqqjHEj3FY/3wyAoAk
dy6+QRE6ns1JAaFBl4JLu9Z9wyK/JH3FkK7fvHHUA02k/J5alUGTduhWs41i/5DL
T8yDWN8ZZvOSj8Y5Nd9LDkYgl56uXY9zGDQX267Mi8AQTsPL6fHgwFGo/c1r2//H
NsLUndEbDwP7q9YYwL/JOp8GxIM4vk0vBeuRpjpOcgesm7qrNxiXFGCHPt0hHM6h
C/+d/fVyBEitQjMbLUU/Q4P/5Jei28QWhu5CBeIfL4X9+xFiyE5I1SYN8CeGvIJp
5N3AmLjhEtiXQu48C+h9fnpd8wQ7VwJGyC2YPURUjlmli/SA5BLyteEsIjj/dRU8
KLsz6caRmg89TrcZLlVt/FSzh6zv3dGACzEHMqv35O53EhFN5OB//JPMEgs/PYTJ
kq01nGl+5zka0ib1IwSuYqB6EgAJwZxaeZE54IHphFp6jcHv6eHgBbGHriKW5vlp
VProBaSbw0Z/TDMXleZEmh7GtsP8lgDA8FRdI6Bao76MrPljSM249gwnmPsrybH7
9X4QUg+kregyp/w+sBxV8H43gVW6lvV8bFbJt89GHJzVssc3yjBw8NxhtfdfW/Gu
Wr7DqbJEMc+JrmvY4xCNijQwudVDWNwEnTdxJ7FfYGam/9g/dARvXBhgAorW/ONP
57PC1Cy+BCYjoztqO02fFbFxZKu7OttaFAL0dqBuFbb8cOWEe/UYzdYdNM/To+ye
7E7LqXpMEPKRr1dnwBjYJCMnKmNFTccuVwlYYhAoEbX5vZH77ILtkaPw2VBUiZpl
QA287ZnRiSYVxOnjC7iL8OGBmGutcUT1RNvuhBfHAHDt9A3xZ8FQs/ADwZlvNH2F
PFIp+eII99HZQDsV2RSmRwKFu2+feUp1ym55JfLeJkib6LW1DAp28B3lSj5I6fBZ
itLuF7uinGno9aYV0/vRYP2HS+9sTwt7DLKuvymDUCpw5AKeKW9gT2zlCiJKOCtA
oqRCkN1wvR92q7wAf/QuzfPhcjy/umEPqur6i1pzNjE/Mz3oD6YU/2q99PgxP9sY
a6Ldo9MP1/g7Emjg3g27150c3tz9aWIlYwNP8mXWPY3DRuzBdMz8bT72Y/IWxu3v
NnAy0A+AJouIJ678tYFcW6MRQ6OBjNN/Lvul1V4QimHmIdBH+e6qnlALj/Mo/tTj
/lvt/3FhEzNKRObGjSEliuUt6j6EvCoaeAn8NKc7Nx7709SmsD6o1SLfLcxlZC2L
7pbhP2RfRhzmgzNHNQHx5JusLB/ikH5r1B0RKpt8LA9yKs1QwkIZZ1h8AqR2+uwh
bVMvntdO1xyxhdaVUiTaIOANpjj98A61/b26q4JmgWMowoos0J8mykA1jDKSXJEh
3Nhv8Ubyu8a9/KhXxtKch7UjFGgep8vro6z8uVZrSbX8Se086m2c+ZlkGryPxiE6
6RbQTimjRWrpe09D9IdDBB27Fhq4/a9GaSnq9tfdpO/qKamtiLJ65hYdHg/PPiqe
XQh6TzCvtGQLOutuF6LBpPy23nrL03Zvg0ELj8jX+9PB0ZMdu+pGQLXaSAzyqHrr
gVrGOb5X+PSFKYMte86mLyKHTLssMtqfbRX/IDnGdTSs1XxdQH6iPABjEiuv2m77
96eHw6Vi6pgUAsjakPdzb3/FEIaztwcaybWf2nPLMEWV7Mra6GSBQZYmb0B7JqiS
irxlZNDRMQPHiuTD9VB6lzfKTzb0GzC585QHLNMDg1pTFkJG6JumKqbCejkjPD2Q
xaYqp927qTDi/xOtdFxmMk93+IeffO18SRVOAi6PdDs47GAA1+1xZWMn7WQ9ihD3
cArKVNKGSxrRVdSToOy4guxLvBgEsY/uvIJFgGqAbcAt4HqkaiP+eZy98+6vQb1x
wF8Ded3x+Nf5i+2Cr+1UAs9EHHrQcm96ST8wiQWevEEYZMwKTC3XeM9xGsUoTaub
/UbGmLfmDgGGFtkHAESjbK1mR28ip1SkstXJNxCc9cJ1rYqhInBGYVFp8YgkHYfB
adQ5erdxWmBiJxBarJGOZ7MrBQZqcQkwD0Fd6KPwqWEVC7AIdIPHISI2HtWkTStu
HocmxvKS9rCSNe5JgD+PYWUkAlMTHTZfrNI7BXHKYdIb171quxMLoTj1Io4Rug8s
4yEwMyXY5azpIGLkGLgvE9HoSZQdbqITZ4FrXbbsfMOg4ZkZoawBejSi+d/2RmP6
K1afden9BFwrUQlWg/O64RoJBsxbzvDDfbhdwNHcI3QbSH67i/PWSnxSMkw/zQw4
MMAJxEbSg71hjrB6hiLDDJ2lq2rsV4VqJV/uxrYtkVyZY+BudIPedQFZqqo7FHYr
Rh2EylOynEWb3XiG0eW+/fcVts73EE45Yuh2RvCbf4QIpG5iMEKJhSPmYFA0oV3/
W2o8OlthojH35nQM4KMFU/RlofG8VBgXhqajD42DzQHEyp+QQ/ydyhmcNuNs37sy
Yl3B4qcuq1GN/uH+N/9U9LPB5e9P0R77aI0sL2+6iNiRh2SVDsa4J/kMLNRCE5b1
z2LKu4m+HEF9dz9ZCWfLoJDzuQm+kebUfGpTEa+G5KIanor2P10fL0cJIfcZ9MRe
JxikkpibuMAFcV98jQKi0aOqAbrMoMn5qQzrwsZoGYlUkuCbEAFCFB4gKB0hU+TF
jYer8a4QeeKMc7AmNv2DTwWG9X2oBzeBNslUsvBZ/JA48e28ZzL/+NfypHQEiK49
1sJt6yQOEKNkPDT2dkxRCzPg3lnmoOYUgyev5DBBLY0UWcf2UzX8H6megrhjs4aY
YG3hMvIMeh66A12qeitidt4kgonyRQPECSk/JpwGGVrB5ME7MHhYdy+Zr6q/vlle
ySOKUNLC54iDPUWmt7Kype7yeZW2JLGu4PennoKbW56nM7otZajlYv2QeVN3rADx
1Bnyog2QTvQ7QoI95KKJv09UXXKY+eCNjRf0aVAkr+LRSPKtIWVYbqnZz/b9tLMB
zECdk4mkUOziUr0K+zdKAGP/cb2YkW+QOPosM6hMaLZvXq/qoKfUWMq5W7XvQfrl
1sVRWf7gYEzrcACrVsMJ0KCqwX1AbEMJp1L8HUa4lcCRDuuaFRiayEkBAZn/qktl
s0D3RlvvXP+bt94XwyF88ZpGbeswF6TPBxT0otwji1f3SFe01Raoq9HfAvEJC1s7
zK4DK21UCYkMi/fxBL0oGcHy8q4nZloCLMjkUvEIQGO1R7Won6H/keH7Jp8VDgYq
7la0ND/GXEiDj4NtNhzvhR5mUtH4j91MK1V09eDDXycOLMsbozGxl4U6hquxKHCd
IN0yFlQs1zvztVUSJbeg6lYWkzI44CncGfZjV76xpvI/VcliIGed8z5IDO4aQn91
xsPOfindEtL0XgS3xnKEyMrtza6KRCtEPZNzddgrYfQ+qinkLZsBaOSEfT6AQya4
VyokZ/uNXUUW9/oeiTjPpji96523y5R9C+kFwRlta80oJ0avPKvUFG5hsd3EmoM1
ZnzuQLcky4YRXvY9ZYhOI8nWho5lef27bB6Afq6prdBPGr6iAZ1mKCVCdV5KsBFa
Nx09Nm3+6NzboV5oOt9cMVlpNrL3FwS8ph6sno4838M+wpf8zVjJ+7mFr5AqGKT0
zNxWe/GJeCSsNYjL26tojfAg0naTIigogPMOobY3ngCBziQFj1V79jgk4TBfEy2p
IBaJPle9lBxbiNm4j9+a4f0X0t8BtSnsHnJ9wKwuIq7g3Z+12WF68OKgvM+Lyyvz
Ks47zuTRFNmjnhhR5MbKsIDKfDUrExwI3kH1Ge1FV0V2Udn6liFZSyDcQbakFTyz
1le8CLbSjLYrESv+g64Upp09pR59UcCJF9NPilZ1O7f9+w9kwh40Kqi8UT4kqBJA
5aT6Bj+gCCBboFxZ2OvkUwscrmScN73vJxKfS0+ZfhFV6XhWnpChTABQKrE+1bEX
0woDM+3VPjuW/S2ijZx24ujuwA2BAzKs5y3zBQ1PHcM7PnRbB9vxkkdupPG136o7
kHJwZVc1TWvo80u575+J5Nla9OOtCadO0PdfMTX7g4cWZfWC7NoURhZYMzgUd7TI
XS9NrfAstwNGGiVSANrHR1f+uuCt9fAGS69OpZgQBWDeJ2o7eblZtGibIStxh6fN
Qa0PhgHM5BZOZdMV0mbi2FDQzqvBYRwCBPrVJrHSmdLMSE0O31TCWKsKmIx1lA9d
PvOnF5DbVZ3yXnpowKB8XrRMoFhF5A/tQU1ZLhE3xbHfDNPMVTX9eca7LfXdQjJr
OGQoRkE+Tc5qSoZ5/fAm8WPEPA/bWhcaB+Ptnd6dqvRushjGxzZhBJq3AfMgZd5j
/9sVxe/6B6ShsGOuo53iku9MWf+QcCs3/W8iWetgQHEC4vBNGuQ/xzGtVlWUn/SI
nM491uVViKvefLb7SdhcB8qND6pM+zfURfg4b7zGLdp6QlQaIevcPQ0JgYX7NiH2
bNjAUS0+wXVbqjLNSa5G2wQujV608OB8G4otustDVbth9bFXB5yMAbKcjR0MMVtz
S/l7ZmQ8eFg+UBkpdIfUXO1uITRMEh4LD/lxV2HGxtjCVRhcGw3U9ijNGboL2HJs
eg5xoBqIrS22o5oPDbGbQ5KBYw6yIbfGOB9qki63sklYcOUy4uueiz1YKNwNBWTs
vMB2XD0piBFOFsyI6UP0Zr50jGKQG7KgOFQ1l9GDHnUr0c+pr7DtTvfgxxVXjg6b
V1ErH738+RmMMA7OxobnNNzv1xunW+JsGxh9Jctl9/PKghQ+ehoCwmOKUqdLq7vn
KB+aEjqSQUMoSmBRNegMPFB+RDmS5ueEIdhKCLqVcDG3GcuXM6RCx4465ot6IKdZ
EXPwgtLitg2LC787YcGLnfA0C+agI/UK5L5vUK9z8lKwqjjdWCrGndzpxJXSLkRD
W5K3Jnzivz+UYybUHJjEpBCDO14MMQ3lukFQK04IOGrnhL2sMWE1OHLTKewM0G0B
E/prj8nqw6nZFdhb1ECARAP54bOpfpfUf5MiXcd8QFECYXCCBXnerW5PzTAMqwkQ
7C/8nnV9HqaGklnhwZLRHGHRcknbSI+RS2tw4/AFXAzN93RNGhTobKMOyk8z0BAk
NNeytSv5eFaQC7xouW55uD/fF7SYw+fzgkuGmtH2wg+Lc0ESSIOCs13rUQVyN5YI
NGnMPoyVIjuMjqT2SbN3S4A5tzlXJz63KHfKgL1ucvwXVOlel3Yh2QxXcYdVJmsv
Oqg5u4Wj2RVxaF3ZJOtZVW+HFvt8Vz/v3m/GVweObaOoU1TE1eIL9yw6/KNhdJLL
qvFmPf2o2ILKmQkxkxGZau3lfG3lnC0/vF/f0LH+b2goRQxr+ngBx/UuKxthbZbV
h5lahQFMaX9HSWLeijAOPcLa9bvhqEub0KZHLvnOlWlfsMhUPJbWldHtk7XNgjog
ZqApVnUT1EYHsspIOVYeAOVY11dcUAMBAImGYUtC+X3WAONHqiXgk6K9UHaedjoU
SjIxJ7LhZ9alc+42TVovG33kLDpgPQasfzneElufy7euZA934pSQmoKF2EVT/twC
qtgSTGv3lanjyMHb/K1JeAm1yZ/JmuvaqGCgKucmPxdDihGSW5mYTSce3zJYcOP2
XJLJcbDrlfz5a0AhhhXi0NKusO8KIpTWuCcLP52KLXmCHy8igHZG5aZgmObOKjTv
9O6Mnz8oDMl8z5tehacq8MNLNF3tp+2HTC2lAwCXS4fkM06Kx6w2KMcC5kEWNZ7X
gRiaCTNsrjJG++KIYFWcF8H6o+NRQSurFYinC5GvqGOFvYOwhgs/8gBbbSbKfoOo
OuvV5n0arM3s6V9K+vR2Tz2kTzYP/P0GH9fEgN4KXYGskGot6f17upJ6KKiGtyYI
iw42BLmoWfM3LZ91bfqMySkmmY/A1jiJbRES2kSE8+xif6SKH2J79Y0etAVdpJJ1
kvi3MMnnwKNfgO8AuQfa1XM6Ag97BgtdHFtyPsphysT09hYK8GvGU3eWAFHWrDuQ
cKVIDDzECQlpES1Zj8WFJ0iZo6AADu8Di1PMX6XgYeJlB+eR5N46oFJHyESzGslV
DxD+djQlJtHK+cRj3EaFxrGbN7hZgrjUY3WuZORv0GOkzYMX/oNKnIvs7JzO0hwi
6KSsiXrKjQFbcPh/GFWOnKWhI2UgaXXjt9peoR+KK1a8bgKTnVqUiyMiGZVeawLR
msobV4AFqUdJoKjzh2xPyIo2iDiT7hLfuU1FK7wZiza3DPoY8ajOLW46KSftDTs3
DfDFKu281XJGV4maXyX3Oz7hPFWsijceMW2tDu+Lq1TPhEE2Usw24QFbiV6Mr8J4
enh5zGLX5i0kYfVp15MV070HM+EHlGSL56Z0wa7Dn55sZehF0BsHnznnz8dxBJDy
RNibdOByEKeoqZ00n0W0t1EJ/YTbsOB/+Km7l9gVByq9PdXYCJU2P3Sq7wWBNUao
LSCThDQ8J9KyoOAIL9jzJTyeTf3NeS+hk80aBTFy31rN9RrN8W7oUBm1ddsug3m7
7aAOVehqIPU1pZU1jG7RLaBAY1iRfx1C0iqZENa7VmdMy8AJontvXwbDxOGGzKuH
rJv3l0W9zcig49qCSpAqIB5CAk4IpoV6UN4ngcQZt7S8aNnaYAjCggA2rnv/WZzL
U4ip6J8FW4Ghu90fxGwVCiDByFW9nukZGtcoM68OZ9TN8tUV72X6XUVB41ENiYIC
vZLC2hQxNHt19K5U5iDziBlHq/osf7XdRUJgIUmRb+9zA6DCcQ6WcvJnI3INvI09
wxQecNdBuBvOJwxlm0Kbyy+L99QH0HFXzE5B9YQqnal9RoY7GjNjHglQ7nkTfMKT
H8F1RLlhezKgIehj7EsIttoIegYSguUGNSLwQlbwAP8/Ff2G/h/Ep1AZdcyP94W7
Q8Lfg+fSRgL9+8nN1tuDvBwNJIQ43Ba4ppUqTiNsbsPQ9R1RR1iiag4vG7k3n0ZB
ONbqN61TxyPbhj9rJaLMRbd0uIJ7duyXkISN7a9ixlqZNx/nyT9Cheum9iETPZ1W
xPWwWDzSeZp0xodD1q+2Qbh/D0zwDN317KC/zcX/uwTrN/Ob/ecu68ZwVxshJa3D
+HRNgDzL0Rucbgn4E/82ePhm0+s3jSd369+NdwBD0UMLCtned21Yib16YMU9mFS2
hu+KMEVbjGVK1rR12T4gnn1tFch4lQ17PY6ejETqS15bTRMfxsthCJswvkY8JIY4
yDpDyF/Xh7QPaSiCYDbTCh5lQqb73NelfRfRvVXaXUzkqowMenIDW7eW3DLZ3ftP
hJv0D/5coO75d0yreJ4x2DfecM4WAqPjipgIdO1TzTVN53QelDkfEfOsEYHOE1wf
MvhneL3oalgI8RSFMTb6oiGk5e8NlTTQtBC7LSAfBSKY/tzV1dRKfoMZaLqglBFH
R7FzfgOg70rfXKn6riY8iJ+bIl2+vDqe6qqGfdiEtWSjCTchwTWO7g70XVqItAWg
qeV3cub3nm4bSTvuNbv68yQBhHwuRdbFavBfq4lVHxkrYt1Vlzby8yo1fyijFQUj
yjb9v77GLYgFpIegZuOzSUtDSAtTAd9kNwNWalF7WxVu2vCCTRFQwA1qVRE+PN8O
h/LB3PwNmeRimseZIFX3X/obWyf11dwaDtuw/zysUKNsLkqBaECkXKqAxPgPQYqX
tqfZ9kCJnsJ8QNJBQequN7lcFCV4alKjI031zAu914Asim5LGuMj8GBupljkcenv
lSXftgTiGTTSM8mr2gP/5rALyy/mOjmdM5bRd9/yCC40+ECW6XAf8WSU5pLZMypn
uS+q0ylwb+Guha/p+zSd0TSBa6pF/FUsgRlk1/nK8dkx7rlPHP6inGmKhhJSLb8J
6dwypXav7kf1gx7J6svBy/nlJ5Np1q2zTCxHfh5f8K038cDIqon9OrxP5VnQVB5R
6veMPwQIiAng/5QlBuY549aH7krSX2RWWUv4NOUFNOABI2frX3NWP9XQXd7TntrL
w/V39ypRwDax06mt9ugwc9+huWGxJaOo9Np3TLUIsjCIuQmGBZwQxRoOT7PbjJM/
MEjGmSZgO6ZpDe7Y49ZqNvCZur0JjwLJLNgijNH4MVG1AenzAqyZ8IBvnnVkDpoY
kOOhSdyavytoDCd6CUoAqDqGUsz90cSmEctaDtNdQTd2UviROhvARLs/d4BoLKOQ
RUUV2ff8F3DJBPG7O8cmR9bY/FNXw4LYPX/+fvcrNPhh3Hbd3MjJtUOqehsoCqPe
ihplyYSMPEIeqvJ9Z4RI7JWsLQmgcTfuvpGB+a6aGlwDxMh9pR/kVYHVysvXWzgo
FeAPEzWdYoE1rlwavWI6hrqVoak6sTB4Vm0DmLaGgHlGN1n8rjLMN4ITkpINNcmt
7k1JqHWGH+bgAQJxzczWhJqoDeE/R+GdHKsDWHe+wGYZ7NMdBld0y+A57AecfoS6
FxZNkHHKiY14pua0YFzHQg2fOS4rPWHVayTDJcVrzgHDwGr5wx4G5mt7kk4gKpla
y5dqfd4JJ3j2/R8R+BHvM4ZmdNEmfQGDYcHu5+I8GZM6tx0UIDeVr1k4zqU44Nvi
3pg1uGi119Ku+d8BD+55VbIotb0qzi8JBzP7JwUvvohzToE8oSwqef9x94vLZV4f
ahjN73yQbKB6Z3jpTwvRQMnrLURb25PQBN07Fp1WpHgqjF1/5wJI54aduFQs0541
EAGjmKdh1lW+PF7xi16b0C9LdALC4mDJH+yjh2fOJuUxLd/q+ElpJxGqFNmMZS1f
ekF+/PcLXupbze4zZJgGSDxjJbBCmNu6PhErzL18jcqjvu4TYxTfUvngUOqmsRdw
j9MLag53cT1iO0nnpA3P4ZN5HKYVfyYFvCwk57x0PjJpWMoHWe0557iHCUy7Lk9Y
Fab5Um0kerJBh7kMu8163AohiugeAXwpBz7vqJSfX0/PKlCsjauyg2hzWWAlgWNU
rMyv1lH49WE3LUOBH2cLX1P6sZQoU9ZMEuY/dX+n+UR84kXK1WQaITOI9QA/4G/3
12XPKZ/oZQOQVjASWehwTkOGipcipMzuDR+71kVQG+Fuw7AIrdU5eHKorhUh0nPK
ecKws0vK4TzLGFneEskgJy6oJ6aj+HyXVT/2npamLil8MQPSPbU8RsXC3+4kh+9H
kzvbtNOJDqRtzxRBjAZnDhN1LRlkrYOCR68rO8NM0HybkUZV9Y8lz/eAnFT3zpU9
usvcsUYTjbfQUSPREbsoZ6HBNNaOCbLXZwhqv/MwaCc6fajwUdyd5BCNDCjVD7V1
999u7mNfhQiMNRrgQS3B7/NypJ84PSx6ozRFyVNZe0wDpGrbBsoyif9u6F7B1tz4
dedgfnnP9JnuyWnv1eIlK8M8Dqt7DnIVYZkyTxT/gskLAWyYwMYP+Wkyu3w+WgPR
NB+xIlmrsC/TXCzhJ0V2XWa331Z/rCGH1LAis/3PiqdSuNV9JogBkjeJDkBvF8Qf
qyzk9IoRxNuql+e73ZrWxDKhBUiX1KOfS2Eu3Myura/N2+53eaUy3vb3jm357tEz
XaGVIdoUiIL0HCqiyf7M4B30pL21FmSOHOsRik2V5jc4kqLiizTARDRptyp6hSnv
M5LDtK8gLMJb5jGMfy9ufwzGzmAiLapKXkRacDC50VPlfoIQdiyMBjA4127bahQw
jEQ9aomz2RyvZwI4dThT8GCF5btA8aGuBczfHFqIEJ1mvdXvAMfm7YckrXTTc5Sj
zR7Rb3hvyMZBbZzT9rnb3rxMTxcgREFsdRXNSSlQQl2KF/NuFF/qZ/iWSD+TRQH+
dYwosxKKj8pA6lL21246vgxsQRNiE7UqJjxzi7opuGRnR653iizNtTb8nnjxSEi8
mrymp4XLSd8cyy0qyuG/D5eLKGK21gkPHk8nBmYFFdJHn2srRsKdiEBB5y0R6S/Y
MdwSFLMLzHZj5VWPVrTLKXQro+66vzb6baw1F/02QjyV661qUfDZk0qzyejGVMmx
n3b+Wp6E4SMQF7cG9uZHuSgEtoNyWpepMKqPkrcqHQjDFM9scYgviF1F/pqRzV8K
/E9ErTyDQqS1M85u5QZwt/p5qq+h9RQdwUvArqXSQFc726EcelMRXk9hsgpEY7yy
LvCBlQyKNg9iveJJAZoIDbjacaEmGwiM+KpTJj0e8GZ4egqV8T33k4ExsNuRK0P2
TU7te+MxRmXq4RYh6wXEDhOmSX7LG5ZawJbtsQVE80eBgos/zrBnPcUjYNsv7TWo
t2YYk/NyCm664dqIaXuJwYCwEamxkvxIYSBwpqh43kVd4Fe7L1Lsfsp2TFhorjBx
RO5mOjtiNzgxRu27i0LV82vllLEtsbN6685rR8GutSCLHrONW5UaDskpBIrdSAlh
AdJHb2JuJnGmD2lFnw3q90qvfQRHnduC67GPSgYMAC5G21gdFXfvFBegEGDfXlWn
HZPKp7mPmX/LgwLcvo6qS3ITSy3e+CNpQQyEpiY3gtf97BRKzBH6DFAi7xKA/IUv
W6nEjdqrLeEye6LCxz9S3apzmiNMpWtHGOMZB0gN7TiWe/BRVKmUy6QBoEXNI+J3
+cEX1k4LbeVItYtrsoAOVrrI7YWxnBTKFIwPxlSsYrr6rmmsrl5JjaaV0uuiuUIv
SSfHIOOdDnbO61AEYaAxU4RA6Mp0Ii1wlFo6QCHVAAcubWWEU1AKSE1N0erxqhkG
w/fn5PleBh1qB1T10DlQwNTaXX3vKRzWZrpa14dEhxW9e9KlIyEcJncmVqYNnQtU
EauFpxZOkRF/kq1kSNmPtaxe4cli3HbkYopuOalJyQKX4Z4Fb9OWuTcyV9/fYvdY
mIGw1X6fmEZS1bwxGW11VKhPUcNxAkSkxlJRLPdjATex+nOW8Dkgei/O6DkC3O46
gaPAw2j39JhUXROvDEkkym7Hy/4fupVMPRnb2SAtUhS4bX8orFN1ewwTgTLLF0vH
wRkpnij4hHZtXWVVS9QRXL6tjbl6XhUbS3Z69VMd9GbCesRXW4fIN16vNFgoQyZT
fWvYc4djWIuZEJQ6TVtDS+2XgyuT7bNArTYePNVAJVp4WsBYtT18T3YQvq+6Tx5q
dG/mzBwmlZMys8OD3qIHk5Kc/DA9HNEHLNvThHYBOu9uTE7I+l3ZGYe1NUSMZ6ZV
7XbVlL5oQ0d60zXIKF69Q55Pq1lTbOgcjKR5Unat6hegwgHlEHnOgrhjj/x+wJGO
ODTigS/Kx//uwLMi/DIteAAZtsnFDpP81w8Hqz6/E2fgCKUbNO6yqGiqd1sY4W98
o1gsEuW73ndVgNZHH3CgMUTYPDufadUv/KFcJdR1AVQUvw69+tO+/2V4FJ56eRfz
Ba9BeMFmf3ZIVwyRoPxhn5qbi87yOoDvnCJsa4bWCgi1ymR9FO66+AQ9FycMDQUD
RiOZHC9hW1E9cQInCrMeaPbo3m5ilfBN+kgM1Fijpk8A2S/SN1BZNvnTdGijvYJJ
XzKabD6iYSeFBn4+P5zZ0zL9amercPaic7+q68C4wpGsCZoZ8w4LZ1Nb0H95WbZP
wfssZ4HvdRRr+EhWZyD3hWKoTYoACz+XdWjre9/AaORc+acXmK9W9xBhTg0s+FD1
k0xsDWFv3yA12peSXc4rv6mx8mVQDipaVrwEFA3dBI8t9WZx7SvU0rD6a3hNcCXW
suzycGzGKmM2NBhUZDpSOwon+aOBSbCYAaMXSTBVVgftKeSIYSYr1Nj8fgEoioq5
koYt8oX2UJrYOeBc41jPZIs7eVDGfYK5hkNg2pyR3WntXMGayQoqJt0Q8POmQEMC
Tt5NUhxd/KiiwRdqJfHqETObcd0XRG9vFkRonO546utx6c7r/rjfFaIq60AnKOSK
3sBG7jDZdQyJkDcmVbNHjLFFVp/zAUWZ0VAuGOVPLQv4g25zQncEZDpEgG/cYky/
zQhcoayZEt+aN8/GPmTavJYk1HuHVzrQZDG+4Dic5WV3+3qJXsKj6beN4sJMgOm+
grCGrIsmLL5ZvQuH7SdFG6SzS79SPqSQbXp1fUPHkHQX/NOx6io+/Oh5YS8NwI9b
g4xxm3i6KPH0/dVz1XUxfGKF+UEBTRjlEh/cPNF6ofRIU2kpWp6+SBW4gscuw1SB
nAeSDN9h27fcwc2dy0timZkskGdjroUGleACDyfbfh56qa0kS63k6arLVz2jsNQv
008sQUFEJpD70BXtDGs8r/rl8uybKSaCwU3wG5iNoarWDuYeT3DTaAY98eo9pa0V
r34QUjtkCMqaq+dJ7fqfs55ZgtY1ykVNo7jmI6WwfkIJcaM3zx60A2glvESZRkKE
b+wbKXeq0Rc7pLaO5Kths1EEFqBLasoBBCmtpmY9NSdjshOXt04+STXwDjgMqXRW
/DEitATGNK6mpqSv479TyotdieqIZjXwDHxSwB6zBzbpMN5ho5JVpqHxLd31OTu2
6cHhb+gXt2zKAakk9xTUauPYAw3DnIg8yg3QSjj3CGuvPrnhuvAjGWEOBiPQlBWV
ZZOiZozVylcXDpBAsxlVBEWuDPW1p8/vmeKQSsVf7CUdkO8xQnLeOoRNRGueOmJw
QRtqItg323FyEzmsOH2gre+XtRES6338A2YhlvJBMmmX1V1ObphSOIjYZxBjut12
5dZM5xyB4b+m1hcHO6UwKmeHt0m6aZZUEWUln5NhQDbo1QVzV8QoU3PsT8io+OyR
TvFvbP8ghjliwoiwOp8fnWCNwGnP7okoL79dpTDECTEdE0FUxh03FUZi/SuHWBgG
/c/MQjBgVJWYT8PlWMcR7y5abAMBslU8+YsO+MKHi7OIFuiXp64eiWGQXaoHXFit
EJC0B+E1u1UiCmNU4u7zuHnBNq+9sk3rlJdTuTNLn+jKFKzGsH1GFcczy0xtnqJd
n7NEtWkKi55fT4eFrAVsfOw/CyiqmQUHoYqgbFuQot25mZm8l0ERKGswBQNvjVUr
mweaQEzikc9fjmcDbiVnVSWu5HwhPSuWvvj6LCvFhmVBTbSfVfrHW0Qi93B0dfhi
Qu8CiXz3pr4OXe5MKNZ5YmrZ5OcrANOFBuuZGHqBx6HEShGucW0pm090wcgVOpLp
0uw9CbK6y/E5KMrfQ4usb7AwNdKUlJveTeo+pBJYe+gPFeiza/F9VIVEPkzu0niL
6F4LRqdDu38PPU0XJZsBBWjOarg46pAiJbQ7NZbuopd0SMALiyUU10pzGCCgq5mK
4i4SgIXn/qBaTeJ5e6LABBtTf3TxM3M5XeZSuenox0OofSyDUjQ4gAZFqbk+sEmT
+8StJqtWDsc2JEmz/ia3HlBY525x6mNNbfwu43FAsvg4Xyfk0jGZipMUGviGf71N
Ug4SFc++h0pk1QWamxvTYx21Bo1WLzeE36xc7aUmkL2B43DSJs+TEprl4kPNiECV
b4HYFsmaDdDqOiWzURcE6nedcQShvf9dkn6VWAxbNGFnKUiXMBum1AW3IEogYR+W
WxNFrUzBuzEluOjKaBzwVgjCm4PC8aFfHcsvrDg34L9Bhd81YqO2wk4iWuy3jaEh
V4ImP2NXuI5i8AqeFGT/3qeTdmNyZ57LLgnvnlq/53AIydR/e++D4AF8lTQZJaQD
kJl08GK8VGqfNqG07LJ06oAxsjYn73Tv4GrYAXdTmDR00W2UXYQt5B2a9PP8shDG
mihTm3wTzkwyNi28KYaytkz0NdpoPdoBQeAIvNFkSUMBjJv2QEhdWZ1OmO7kIVfr
u6823kyfOBM0/3wirsLGmp3WmB4+Jj43Jx/wUYZY+b/rTBM+gs3Fe2LEv4LXT97C
1EKGRGe2JSWaxXL09AZBLmcN9AJW6sZe+97/xKx4hsLPipiJgUnwtfTFaPsSeG/u
H3GzIprh9Y4F0sQRKa9tgCp63V4TmEJSfF8H87rQZ53lr93MqF/McNeZNBnHlVg9
AOLbHY64+DK20djO/ab8f00DEqmuI9ZMKtsuFHoKfNiZuNEvo8Bfho7u0XUSk+hP
G6UFImjUCPrGfM6NdDbwsA3jSk/Hs0VSjSuJOPLpXqhToFrRt6gs5uQwfZeN5Ji+
k0sv1yHzCjgcdwX5M7hWW3Z/R8IHwusAj6J9+IMfyE0coggf9NtviuHE3tzFyaFj
8DrioEvF1i6GbNm7HPfmKR+FkIjFjV/fzR50R21u9/WQsvCrOezI+lZq1mGqDsAP
5+r/8wQpTuIPDCXbzqiMW5QPzxXoiDcbXFy99sjDuiKsM+4I13QQKFWkXVafSQDk
k24+Ej+HiiBylbIFLYa3r7e+/VgZRfniC6/hqY4bBGAl7dDcr4r1ZmBcwm52Bxov
hVCPUcazgpz5LSAq4wjniAKGvLIJKC6h25IcOdYGKzAnmQKMIuWBO/VEbAHOlXZ+
G57KKHQlbiqVDXc+i9exjhnK4YszpBfNOoUdUbjPT0Bo9jmiaec6V1TMGRWR8+d0
txR3zScSCVUngHozph1ZtcXpjvbWEK7e6MGXaHXfD7OPxcggl4pE/z0vii7avlYg
P6PDPR79WZvZI3XjssA7vqeeGJ+gHqZmvqLmT6aU0tPTRtAERYcravoYOb/7++IP
arD/xcXDv24pT1tay5c0YHP0s5E8gOHu48A6CSTYvXB4O+wB8LobGUDsph9TsRql
jNLAu1JIFxGZhDRKR6N8Rlo4CLuzipCtAxkcTKSDLbFY/YDRtohiw/HO/hZFmxfp
/jbJfDT9lv2PPvnr+I+grGGKsCnfq2twvKTWKXyQKTYqh75GOZYH4PnkSV+yYkmQ
3H4DrIWgOQNTNtgia0vyScVG7wC6zBMYiei0fnwnSZJ3P9iQYsMS7KKbwGZD0UQg
6zvwdeSRnO3k6nZR3kLgKjcG074YumCdT6CLiYbgS1zbZFi9TIxucj1zqYdmQJYC
38bnas6VUC5ZwfBiH5AwlsaH9LGTycOKVGqyD3nJHUA4gvfYnnP6+VlK3BK7Nx0m
BzAvVZr2/cBhpkLl/2MtnsiRFQ98Q57q0P+QW1pN9LSDgWTr12b2oSKDVFCbOlRD
TAP30mGk9aRARbc2uDhLC8XF9QcGvdKpXxiQ1fynhKMCTEZXrCw/dM9mywYj4be7
vsSuLPANNgMCOMo9shwhrNTXkKjCtcm+oSeIudJze9/Fz0Dnlx1UmPhujFfuqXyD
v8IWoKPmAmwyhEPb43q+ZuvHwmwvd4uHlmff4WaJJVVBkqEgoRrdinozFXQ5iGMc
ofvwSezZX2xn6s8r5RW8lXDeUI/ZsqqHwPQKI7FR0aq9UxvzVH4vVJgjuoW9L+RC
KDaaVe8i0V0xGjWPeKxnqQ8a22YHECdrlRP6AwlfUTcNh7UbEWMHVb8GQk79UQbX
J4IZLMC02PT40h/Uiojtl92lnf4+A+CpkuDM3XNUuBbQjY6UxvMcXv8x6gA0JuCo
gvzAwHLHJ8sWVM69dyhHRnG6qRtFEDMGZjCSgz7X6A+yh7W76XgB563wEoMcOk/l
aKZOmDZl0GjXmARqMVNujI5R3o++7rn+P2oj602kqO3ohnl6GbqSQFMn32/A3Ah5
FeMecOrTqr/3DBMnrbRm6mPvGgaEdQYQnFQq/COAk8kK8ITEKIR11SVIVU6XqdPs
1pYxt7sx2StRzQ6DIF2ETdyMoT34v5mTQmpfabUsXm9D4arBXz3PYebnMIB0Fj0/
auZkus0uKmPbecxvIHl9uXEf6Dy2hvYpjsWx56BYDUGDlfT1EnD5BsWFVG/i21Fq
85VFi+8RrVpdwGTO8Lk8CdqyCZ9tnhdgj3gjX/NPcQMMhsMjvPwrZz0ag6TfongR
OiRknXaArNze3Kb17AOoeChsTDgZ/o26RiJxmXHOLbQHFRZjv7CzSEA6dXhpU9x1
j1ORsX/q1os5USC19gostMc16FxJ5G7khis0JX79Fkvud6UxuJnj7JLcm3F3n2EP
7qk9aJjH/6/c0NmbBi96bMU1yWvLPaHfPg0iTKP4Bb3a4A2LVNOr6SZ3VLISQC9H
VUIo59Y/CUXIYHH7/kPcKPaJe4JvYFHuVnRCqAiL2YCkZWNBW0zWfbpEP4b2rxJE
xEYLut1FoKINjKTWzL2EGu8Zcp1bsaY70k+uJa9MtoqEp/SrGcBbe8wW3tKAq0Ai
jelk9cUSezgJV2gIsVY8dyr2SqR5H2KdEeUF3U/xhWaSzcOthv2WnU4+sWyJUnXR
SpJwxORqFv1GY1u7NIZMoirq5h8dZZA75On9gui1F0l+nEGJO1hqDy+qr/mjwnlO
gV/zk7mq8kY8WzEwJl5rFg9Gp3Rm0zjXqNYFZPGw9a7OEIuHoKO3IkY2TbqzhqZm
r7B9aHEO3/yECcOlQUSSXHQ1rPW8LZoJkUn5+gJjZzEPCQa+9NX56n9TR3ZvlG+x
ee7EWhmnNtZUGO31tDSNPPkWfuOme+iJYIAAN/7upSx+o62TmHCaGBQ9WAPbxlrW
0QOk3kDjDAQiei1Bk6sp/AnF08NhzHMxZ+iNOF1xFyQRvez3igFHPMdWE5YA9gbg
pOjkkO3hGVoZgO8f0XOg3q5fDZXSFk9Kk9oTIApqny3OqIp1gcclaznD3Q5nfN1Z
2cIafzxxDlAfCUmo4eBfFCLrSmq+GnFwxqUJpZLh/1xaBmFPFwL4njHnrk42Y86D
r2RH/XsDnomhepr8oDFf2FoOrUze//Urrrb5kAivPhHDc/d4ehZoggh8wDBlYNWl
leTkq6RYup3Kb1SJ3aTFTofmoJHZ+VdqLKCx1clnpisQYfVmxnrBLT4rHxmHBBRf
ei4x8PLhIyImjdllC8nFuqKF4TNlBRteI8D0mPiJi1YSl1Pk7I76CWU14md/asvT
F/HYdZq96W8ATMsoIXpL5OpI+RQCaURv53Z2k0uLjgjpFPpTaMeTmEueOjmvJxOb
4yN0A+/A0NIJKFg1ovnOqDFydffqnVcO71YqRNdh61bD76CoNdAmtvC0wnJ0lUiu
R7nCr7nrTtCg6NQXYicadEfP2ovFd7UDSMoh9j+KGWrxWLUcGFf3ZvaEtJPgyK8E
72ao28ZOq7ty6FmCkqrIzDxqQ+8pVbKxk2FfpgmgSOw1p3KVjXLtWmQx9n6r9a7e
7yO8MbhwBJJJbndASS+blserfL1Eb9i08PsecQlySWmDLKtAaTmkrx+NHjOQ3B24
+ogIQGUF6zXJvEA5fCroGRY7YONZjWG4QmSkNsflf85WFXrad+nhTs+XKr64Genm
Z65crTQnF7/jb+xF1Foq760/QIHCJvNIpEUVpbsk1GuanLmfSXdEZv0BxLSHa5nk
fvzbcag3YCRK4gRQMXOpgocIEdEWHBLmYRHUj48p6BTxRUUkPWG6wx6kFPvvCeyR
YzY5vG4jVWcuV1J6JwJ/4XiT/qXf1wEhdFzfdeUgqIDjfKoYKAx+niuER8GU1ILr
rjNESrQ7pHe5keCQTeuXuxs5V2tUr5kqAwn1sYOeHtALQmWHN4+X2F63pDc5GVwy
l/uX4YQ/0b7XhW909qRoDacPqcC3FGDIl88t9LqrK9cENi8QWhdx4bB9TDMJ70mo
YckYGiWNus2rmIiJ29Y6ZXSAixv5QtbOVTZGmHDSLnKZngdmn43ejgTKGuY9GQFU
WTUFKtT5C04xiH2yEusVS/MVj0pw4NH/GRa5Uvc4O64vLJjFjSivyaE39uH3ecEb
MPwKl9UfZL0klC/SRXOQSRqLgO5ad2htBdBDfzqkVDPCrsaKenIJ4ylISHbxvVBC
EW/EhJCyAv8YopXPkHy466Gz2/GFRIrXEy4DhbsTlKW586TysR32K/ZFR3xSQFCQ
MQwP7eIWMSOrnFaykngH4pyenR4btAWMa3KEsJ8CBrq0I/bJPhW/raidvjOSYb7w
jTujJT59fyABPz/gOjdkOOcGngvKr2OF8XAHqfl75OKHGyWvb9p4o4FVZRTQBUvt
8SsKJISURX8HiUJXr0vs5sl3DE8MtxxBkmVNEyAOvh48LwvFEmI9szHl7sihd+g6
v3yKoAVyQMtkIbx0a10CgMZniDHxqlE9uVdCG0dgN0kgLDcRy3/s9NgVJEBI4+kY
+xtz4PNLrS1t0HucE41iBbjRqg23jFoyrPouNf2trQnO2cMkEhdfUejcOskVbnYu
or1Ph+Ubd3dZgpVlJ4POTsBAdVFF0LraylXb9Czi0F6Vod4DC+6TZPNgKV/HDQgO
MJ7bH+H8qExhINxgpjDTXZ/amqza01vAqFW1Xv3JXhpPmOd2A7iEc8U+1rLOwCFu
FwSsu9kJu4LL8ujCl+xm6bAKd6AzqQqrXWEl9GusgiRYNEJK4yYT4sAp6x5YKzTh
gW+rFsvAXOLZQA/A6Hnah28cRTZiLs+r7z8fyRmSbSxUHWDPuEWI5VG2L1nZxbGo
CSuvvnulo/q/8yiu/kaiE/R9CISz3re8Lv9QmCpKSSSfn4ua6RgxjRdnYuK69HuN
bi6bmGYPCsYWsH/YACLKcm/rZDmnF0wtWrLuECdBGtg4gUVdPBaCZRGcPAD6bMtp
Pgx9nHQcCSLLTVSYlBcNYSeqgIiS2FV2xur1jlvdqxBZiZcV7vYsR3G5oob4ffdX
/Md3iW0iAkdx7HC88LYjkNcttbHcHJfK7UCiOJQTsUBYlCcSKhPniAFiG6/b3KL1
WCzq5KmF4119j+HmpFQ9GxYEN5FpnT4nWc0xZd8zR8UBmQtEv8XtfYZbHj3I8Jmp
WYjnOBwVE7FT3hz/BlosPkt8GDBNXW+rSlYsQf+dPMViq09Fs0+Gzrd/zwLsi6AO
cZazugg4zKFb9eM73jC3WeZGkzH4B1oxY54fn/o/yrWQKTb2F/NyZQiEwxkItOpS
5aiy/xHXBXWdXrn74SZQ6o6yUoLhG7X+UaYst7NyQbRM1GYv1tTYucVczbL7dxeZ
yxMKqEZZqr3CYZPAHp4xhnIYhDumIA5l10Px6OkkS4Zbhpx5NT/gnSwrsQVWA0af
W4Bz1Tso2CYtI95Ux5tiWoc2sEzgJTAVDQLdOR1Qf4E1RVQAIWDhH/j6nDhp2NlH
7muBiQxmvADHrY4QeOGZ1EmcLP42ML83Xz0fdOI7qaX9mw97/toGZvqg4pAlgjPF
I1jsCypJjbpt/Q0+bRV0SDKZIxlWjVKyIfNCA0jQM/Tt30sF9h4mq3L3MSsr7KDS
c7vrqf/JksUEP1hWC7Mmdfl6YbIjqWEkatoW4aJJ2AeUZqh3eMJjEa+uX/IUBaag
TCWBdYiBwEyXEVdJVwKSiOnfzf2G2ncrf/iX1DGc5rAsFVH7r7VoXC8gTn9MDz3u
wb3HsIKaVwdRjPo2EzerefRanlp7tMgxA2KrQ9K7q274jTxSezS/lMW/YZclnrwi
W/kN36wWKqr3gTABLgLW1poeoViLHU5fSbpLSsSGlO1njt9yFiblZgRGJCLmS4GF
DFvtsPOb5ZW5P7pnb7pdAzl9p46rDyiCdY9KecXvC+2dhmAp0NpIn+sB4FtJiDCM
iLoKe+ZO+2veXIJIuOxrn4LqyvOCwqQhORocoyZC8F8/RyK71IC56r3m0Gsd84xO
dIBEfwibnS5BC4RMYvlOoou1Je1CEImCAEvGy6CgGuwqk6r5EoAW5QVIgvE+wSGe
X+qwj0qeha9TpLGPgt2WoJ8kDrBoOwcxDeyeP4t+eFLHrEaYzkuHueVrHP5iwgFs
c3DzvlSs1aJRGKu+a5fdOzEtY2oR63fGBhwJQ7/IHQIyZE8oPJ5WHz5qWCIqAuEP
LrsBU5LhK6Y881DZGTuN5TtEMfDZ7HiCpvA07UiMpODxeQA1IAIIfXcn9C6SOEdj
4SjDV0Yb/oWqjpcMFHbOsgBQE1daXytQ4W+X4RxkQ8yrdg94Y6yEw55dkHkUzZmh
Hk8USZUPY5xKFYjkxXgXlQJGOIraJzvwhe8J4ugK/FgFEpFl9IzHpDEXlvrxOg4w
SPIQmKAdzQOI3h9GBlpjOfTFlr7y79UPvH0qEiLFhHgQHJOxCKq5Jjk21iC6VFd1
hsrXUZVnvB8TpK9cjplbOgkjeqdTEYHqRSNMbyZ3DZJPviNLtHn6GFlAw4pPXkX3
DKdsRDfmDVvc994MQIkO/ZDwzwGvehdLENGodG61UNjjV0O5NxfEdQwF2rU4s/86
k/soG6Wmf0qGB3Moh4HIzlziXD1wl1Xd9PJy4wJKoivGGaIVsFipAgy5HkkNCxVn
lR2RDbfo4hL57beTpH/sRb5WWjySNXlF39S3sk0fDrSnQ0tjyIJ9qCbvztiUIhkH
DpaJHyAnzAZZ+RyWjwqyWc8ATgeasVdQ/k+QCkJtKXYL0wvlwhLqHlJmn+g9LcS/
sxnRCG2IqfrpylcCUCFXbroFRACJxW0Xpk/ZxMFK8X+59ghAHZiotTuO3sq9NYA/
1yqWQoCEa5SgW0rUuOBpRwJLTWUQt0+M7jwq1k16bkf2AH7W8ot5nuMjoaiNfAMv
kts0Y14LgepfHAkjKHM0tS5d+0Bs03BSIDIEaBJOMtSdVSDYTNam4n1ks1PpPa/K
IztWG2I2bKgyGVPh7fOaEqZfNF11iP+S/Ww/WSS1DlkF+7cm1JoQ5KQKax+7pBnj
kdjLaZh82NOzrAyDaRJSjhXMiqbLkGViYqhk/ub4F3VmSDIAeCaxsmkoQhtUcj9M
zELNDP4KDNy77bBeBXjvI1f1auiESPWpA7mNM40yca35Q7KpYxLJ2wDvdvbj2kwX
VeyQZJ/m80tUZOqRW9GLE5UsDoj1TCjMOFequhCzHEGVhVgtlsSNYB8aUEx23iHR
zcHfdXPb/ABMKfAtXV2rBHvxKg+elTZrpkfgTx8R+KRmstixOYLslTJLhRPIKCyP
BiBik6Wy+InYb5u+tpGARIoCv5aokO6npNiOzIYY0/L5mx6YLv9qzCZwmV2+l/xH
LeBFH4hu12dYSuxQLI8rCDVf7GV4Z2tfc91xYEWGQDJlCVyXuvfjHYI2d6vrVI5n
Rm9aL1Ia2rgOlum8zZ/NMgxtTzAUt7M2jQD5TKiGcmG81vcjtmx85Kwh7iyuwx64
tiPDiiJolAaW4wKc3DE1lCEwul+Pasx5ET1GPJxuWkSIGHvUkn2b2/4hINP0jrHS
HuKhFbw8mTLDOr/xGvviH01jXJ34ueYqSVgziqT3ys0sH4p2GU1CAzlhGYT6N7f7
KgwJybAFtofoSObLu1ycEDTr7hl2JjOgNPDtC6K0vhtkiK57jcjzk8v9Zluq/eVY
U1f6glsT7qsd8qInRGS6465ZDHMWcx6TF3QZjQiIzovaLdw6VOKzXF4GEgv7pv63
leboXroSgpMiKU5HTxe+x8d4J0cdE/r/IP/43RHHZk882oAWLjs17XgrtSEr2vTs
5zIgiW0JATimPD4LYNPPw3LpjDILmj72EIEkSKpmdh7wBWg/1ne1tz2NgUNgvpCC
+QZdMCXttX3gDij60bFP9A+oa2amdm1gJSFIlEFJ4FM1OWmy8TwZlJhLjSHtP/Yi
8NX2WMv+lRZ4LupeXSbWejte5fb8BxAcegk45ESRQhv3eHIWxGSGPORHchlWe7t7
Moo2esSGQKic0Bt0iowbqVn4trIaf9gNdejANAMXKSYVuqwwhuTYrVBv+0EIhI4+
WQv7GaUHjh9DPUxOid7itHlY6d9Qu6L+2plb8SeEuG4L1xSU8oVo4Pkk5ECoNXzy
Zb8SAQQG7h/CkwCFH7PbXDEhwiZapdM8FGQpp5bFk5u/mEjnodLH+v5ImxyuSMSy
SoDJU7no+7xZ+tBAbBCfzJnutRXYJbS0la3vUZWEce+v9o+6jNmlFY1JDVqtLyRV
eEuhjPE8ZhmOTxJaLhYbtuKjQqvsghzYqXWQ42u7IrH1Kb8cNdrdAXxwm5B7pg/M
pVQUOWCa/TalyDZBoEYu1rWHxS2/o/cd3rH8tLgA8hfRC0pehgh+gEEBAL9RmRXp
pvJnpFP/d/OlIvRBtC3o6g6uy7GcO9gQCiO4Wly8Pq7PTRPwp1xTEjfsi2jXO3Lc
ZluPdTXFZcdKHzQ6OZ/WPSSLSh9l5eylP45NggJZRJBgyCn7pm3qDmBvtAI/FSjm
jD5KPMVgqcRO5G85MH6PFb1EonCdIGaptgGvCOVgojitj2PM6pbDDnWY6VD8NUxT
r+WmwZLO20VOVp0IxLMjJzAdSGEoGUxFPAP8tvXqlOrBaNmWNVGUgk1bwIID63Tw
96a91Gu2V+k+mWbQqE53XobVYLfKM7s+yDyENFjtWX7++0hw8i3bqsOKld0VmO62
u7BaWoA2qX9fGiBF9pV2zh3I51Ovjd0OWpDke0bTWsEHYih4gqiXKB/uu5MoZRYb
tFslV/y6YIGqyBzqSPNU2e8O4TeyPQYXiZMv66PwojMcP97gwJafALn5OIvwV1GH
2jbWsgziVPdDZrH2VSsX3eSCjHU9SCYrDlsGOEnNPJ5pXluftmLOjsX1kkA3r3iB
LrtSSfktwQWjsYUHVJl7i6tTCjay2APhm1ujofYwWU/9TQ00vVY1a2QoZgQODFvH
OW6mVupC8M3raTr8ZRvaa8J9KFG+ts90VVAgd7VVidhJ0M3uq8CT+Xbj7mULWwzP
dHfOBNZ5VYlGvzm7jaK28cl6GO6rp4VvtcqWUIB47JCXk92fu4GjSRF4Dlfa8D67
YVPx08VpVe1mwx9X3Rt2pD90uZn+Vvtshzp/5QHTSK0HQ3rj5B0LcUE/6AZUfWuY
RSUQvWAGHYCjqImfAmeNkD+w8BSeB6Lws6m41O/N78cu34TMMrWK68lSIEyADdB8
3Fg61RJKoQ3ldYqF/3AjYZfPJ8SbfqELdg8a+N/i0rUNL6YFMjMqaDHrZR3QTgNo
Vh0Xm8jgePkVitJgGKAp2bXuJ1fKCV3+Mi7NNb2EyKU9/sFFarUwWmUM1obXVVFP
X9OyMC3IsKP47cJ7T9ipbj08M46/W8+lKyfqWJ4Ue1Ti9pH9Lli6kuiPm6PLH1VC
QfiXTd+o9TjcCc0jHeXojur7ZtxLDwLa3TihBVNZ29CZeSB2Npngr7gGvQF8wuHj
Bv3CE3UJHbf35PLxTYzGHaYnN0Tx3c1t/GChIl3VGDU3RPugESF0DkaVf/aDI1ke
KxR3Ikp+PMP0dq4inU2CU5/NkcG3gaiOagfBF+sN0YNpyOTIaZik7c6dFDKZPq7y
AhAOVId3y/F+q0LRJEKPprsZf7WSR4uvzu/yjsUS1vknG84cc+tQ8FcNJb+2kd7V
uLo94bv77lPCtMjMcrRz1OIdFzOS4k7yj8kOEE2duK+NE4VGFP82+0WBmocAwQni
1Ww0vcyIQbWGk2XuJbjqOXkOzBr+kI5Er8fsniVP47R1kJ6ViwARLnxNBE3Jz7C+
xD6qYcGI1v8htfGYIkfnDX1Z8SNWT7mD0bSdAMo8+c00zqfGyT9CA6QeqDLIFviY
M/eEcHVQ1mJlnCxwZ3v9w8HCz8uf8hhDbg23/vC0z2eDOPn6Lm1watO1kov65F7x
Fazhckfowd2b/m5OBAoJtZRBTVeaNmD2vLvA/Db/JePZMJH/jYcQWcolJv/0pFYQ
pGIPRDzjKv9Wgkf1vk7JsL05FJpyQlyhtBNOeUMxKdHAngbBLXkPC1fo6+y4UhbQ
2ZNMyTF5dncL8Edd/o6XGmmCMLPg9spoNlzrju4wZP6e23MBoLRAps+4WMkL5JwM
o0/K5JCGxfDlEeTqNSqjiMWZCFDLDfzmglo0PZizt2CDIOKXzHFwbA1cimFaASII
elJ6XA7bOuJS1hKBA3Dryq3tahzT86twLRVKyGpT5GS3E+lA7WN/bna0eQlUN8oX
E/VkeVSV609aOUAlpdYFePrCty7ZXVtdhyybJp31dKACAOCF9FMaREedbJhi/Qa2
xffviMyF1gXfv99E6eZPJpwWU70viNyEEAIVJc0Zmv3c7MnH3ghN7kWRshstWEsr
ZSgUHW8zXtIZMaAwdtOnxsSc8W1cA/M0FXneozLILA267Z6Z4DSGi6eOPAMIyP0C
/8d6E/+V/0NNTnz/OpvrS2jaccpWnFSDjCAOv+w/Xc3f+Wv3gGe6HRKYViBa6pH5
6Z+h4LTjjcGw1F+/zJGDaXvhouFkV9Ao+idjSZDijg6Vn7E6wmeUcKAYoXdxJpy2
OLbNUlNvTIhsjtBh9GgbRQFPhkGgA9+eXmUBs6fQAUeBPpO8RJnF+0yDoo3Y9z4a
2fmEx2Ihh3/kDeLrwUg/zraus+B8bCV66mKM0HmpYoGHUh6EA4BqsI9Rivj7LUDF
uFqbyScLtNB1jNyX0PUGNij3kNzcoAQh7tdboOFqjSRp7OJtsOA3xU46pFfyVrkt
I5s6H2PEM9g5ykhhFoh0/FD54CRgM1eAql5QUTJWqNzv0v0FeADa0RFUzgDTC/eO
REcWRZsx90P/qxQzo6CIKFLKZm9zOXyM0SIcXLje4SJdO9/5qT2nL8ZvukvTiNgl
6g76fwsB0z6o2tTgGkg8AgLMdQYDVP6IgVd4ovTZoCwN00IVW6DHKKKk59GSQRgg
ZiciULNlhtGrkNV2HhBIFLMnk0FN1y7ZRIzH1ivCQgSxkaKqr4c0UJ7GuGSYabZl
1kEbMIhU8uPhem6FMPwr/sQWXq64LBm/Mq3a7a9U9kbqpO3E/UG8hxdSyALQhXAh
FDb7oiqpRfY82BBtqeFfo1sgls2rLKNuiNQa4/eZiGOh3NcwuXcwcMxw9VT+34DO
Mj5UY6IbEUAtI1Ij2F0MHXBEnlKnP1ynwx54oC2Zjz7Ctrq770AnfHmJ03irip1B
E6jS0lys3o2JJQHQjfPQM1RhRfbVAPZGGIPciNF4AJgWuF6JeNmFk0D3ksnMgWtb
hQ8C1nOm7wnPmX1Z7ct5/iSBlxehOjAZfxCLyhjo3MDR/SdBC/wKsuIxnaTLo/mx
+OihRzVOU+07YiOez+bDMFiA1Vg79wzx1mFD7IFt2C8MT+Zjm3pDzG2Bu9H2ojV7
YNAyLMldzyRXPp303NDHZAY0IyeyHhqPRImvWwzIWoZ7e77tGqm90SpQA+3LneL0
ASGBKdP55gEC5LsL0USHS617cv30fee2ML0J8h38QKE01ZjbctCn4a3dwqW0bveX
UDiLzURQtMj6V8l3Yx7Te1fS9DKbZbzhhq1yXKBPjoaGN1+fbfyxfpCLtvC3LjXh
TfZRVlNjWm+x5/36QW306kyF2iV7yXUgdpoFvrYdOkuFllvccZy8zjRtm9Xy00B1
rC4D0Ly4onn0veF+LCA45PiZKqu7uOnyVwaw7a0FEd/bFMFzOe6ki67S1nLESR9W
2+VQpKaMGhasjA8qUT6Xygfb/LIAa0YE8/pz7vJWWRLeJE2Wc7YathzKJfNw3OGl
m5oAw/HdhYrxzoomAzGBLs9H7rUuGzu1+qo1q79v3AGnfEhbVNU7foT/xQ+x3ROG
fnCsZf2ag3jUekVo949/vtor6gSYOjF9k1EvJVhsRefqviOFEb0icCJ4t5CSwU5C
2sv35m+5CuqXJ/aVGRbgcvzv82dFyMH4e+6JmokPS9KXIwQAEJ1nGtF4AoUz2xxA
H3SX9yG3LW8Hq3tCoAy9Olk83HrVDo138WlbF8R5GL+DK6cDdHv389stbrmsQ4s5
o3/d9A0f0YKd5xKXjhi+yTkMHFK0vJPUgxkSUNU9vItw5ptZ7AzpQsosntRo4BUa
rfoT3sSEOM0jQIf6I4h6lvPxLpcwbeNumoEUdT+EfvDeHff2imbP4hwzGNIEPkeG
TmNiMCWAlGGQ+Srqeu31Pt16vMGFR13cnfN9f+DuDKKBODjT8CZVB0XOywe4Unxe
l2uhL3c9Hou+/9A0ZHEPReHH9pWEeZt+C2CGUlDto1ggs+pRnhfHDr0dkEeZNE6o
G4aLBkwpgq9n/MQD0NcpVqtAbDZ4LbktqmrpJTs3nJaScPaSuXlSpgYGP1LW7rTI
SE7YRfyQOqxNSmkofKdfiovcUAilgA430bruwlSIlufSdj1u/x4zyPdpi/ngajHh
XHa4ppIEa2COQbI9KQFOh/KkGURpOIAR9r5Ibdw4oyHgJBjD0deEtnHt5BLtGwC+
io7ntgmHyaXLndfJV5oxx8e1rMM0qJ2kC8OEgWG5pEFL94HXM/STBom9q9Vj7YFD
P7EzMiquY11had4HpkzwVdU0mVkCHUZ2fMVGaKvn5bYrwp1MjdlXCHmnxKyvFLD7
xGc88d4cs42vhWpONMG9ZBzfwHtcD0uKQNIMKC++o/N7P/XBvdaH5EbTWAk2araH
Ja1N3+1XaO+lyv5S0X/YwoGg3+FW0fY0JVfXGgWfJ4vvNZZOajxMb+goZwDjsiAj
T+RRc7ZVnzYjaX6iRxN1fexgmd1wKhRA4Eff6bQY4pEsJU9hNIu9oXGbk7MjJoXC
SpBQ1Z3u5AYE1Ad9XDOhPW75Mi65bg5/51m+MLJCXTisaHUZj+XAEhsYLJw8lR6H
zwWHgTRforKfErp/1r7ZxbBJj1RysI+mGwi8eYDYNcSL+swgWnDV7I1LZS39C9J4
DrRs1JNQTkpiVCSX6prOTHZN7R6TetEV4Ia+HtQbApFvdh0d07dYdqy1SrVA2xyW
a1YodM3vNP8NExVicodVXjm+EgrfnsVUgrP5kpKEDXrHCLFMTPxI3cmfzeRLphLb
Jmnlwp5msE8mSrOuF8tmo15pRu2JX98u37+YD6HakK0Sfe6ZuNuYmaCEIrU2AN6q
HHkxD32WAdb/T/3kkVrYt5cGVChbG/vrNrO8YiYUyzADeTQ0IvXQriBPy4A+XN1i
iPlZD/m3MCm2ex3BYd3Dwk4BMvs0Xmw60J9hhToTaOSjAg27igY29k4KcbtK7Eug
2TBKDHUbif7opIPsp9wSB5/Rs8EtyB6NJMeaLXHrHYdLoJhjal5Up5+PL2N5bZ6q
ymUG70bcFDlA/FNje+BUNVfC2bzXI59WYu4bWe/VEHZ0C+npvtXNjoQPCdf0j4o/
1lB9a0MfB0K8cKqjY48CsEye8/Cphwy+mIo/0d2jIVS+OUEKe56xFGK9ueqpDYQt
EFEDFINAMl8m6i2JTk5l+7aWS87rWXdCtgXOrn71V98Nb61P33LZBwQ98+fJ2nqq
PyXPuYHXuFhOdyrM5uDGG0CxBMxCpbgm799nGepWDmL/TZTeT91AkmJDe2JQyyCs
bzKCC90J9Z7AIM7BqAG+EbmUvfFhVxPTtyzXN2V46zW4W4+i5+6D3Gi0KUI1ln6O
t9ndzckg1O/stPntu+SZJfuadUK/Qgi1JpvJKge+leueoKhRjXJdp3+s/h0JmRjB
fCrXZGoY5i6dCcLw9QZPpGMwaFfzJsIKQd+gGmy3Y+fXts2ZDAF8X889VvGnh9Et
vok5KrrkGpsPKdoA/ALJSwH8Tx7VoE7joA7hCMw8Q/KKWHz4XxqTgfEk4YkQ5c/Z
Wf/sKC+XbRKjrjBrYhsH4eajXP2uW28ZU0ejSka0m8b3K9S3xqHxKZpaKVj1swoG
S29t151Tu+FGUha11T9tQcau5JrKXM0eejpBikjY8Pg92Wth0cxE9ek+wSZJK+U1
nVtWMRFxDYO77are+08SrjU+o5CEpjaFDHo1rojwWZbWEd01xSF3FIvBNxW/uhNu
MqWvjCFm2VXX4b8T1BeiUs2l1vaLy7e2tCpv0qFdBqYprfxJK5eSp+20KevsVfxc
IFKEL3V0LfTV1evTn55vyt5PlROtxK4tz/FzSNW+RwY3adopCZsk5CWj1zGy6XpE
ZBPOlQcqVsSFbHvoKr+BhkHgroHgwNRA533TINfw4PLWE3Lk/o8R8ofENzr8hIoI
ZpNLwHcauejOSdmHp1vvN7EqHcFPMgvNqdVLLtVBHidZ2AS+Mumn+hFRJF79cKf6
QIkHHIR3kg4LjufrTTzhc95yxuzcCvjIV0IV9PP++63E4dD9vcSQunAMor9sOoIe
GW4MABEVrUjARbefJhKJrZz13Nek+LRNgPUry2fCpiZSexiHEUoWeMUd2C4rmQt1
Q1JfeP333Lr0xA9ictuhpYPKVG0Hf+nf5aJwKDRKU85ixO4+PvpvHolei4hElqKB
WpJmUrjub6/NjA/OVIyjHIfcE7z4pIRVJz2LGdvLlXeVNglZdQaZ5F4mauPHQE9u
MdUhj2PAdbqw4KvLJfx5FkdaILLNFSp/zHxq3d9asqNmQZ66xzo/65RaoibafmdH
JxFHAgWyHOsXlG5P5qSWzxWA0lEZV+Qh5eTOtOaRRO6rwEFPEY5hvLdQNk3671Tf
avu9/rgNKr5XQuQC1v9KNd6d7ElPaWV05nLljJe6Tr2gQAoWhCpDJXI69iV7txLq
ZLmh3hIGVGeZBXUewycgspNotP4uuUnaRGtMUHgagVlKcy/BBgLtXgvkp6CAX4qx
KDFF9MOziOK3y8VOCpawSoD8Uqu7PTZeN0lcQCAWxP/K/OJATz24rKrIbfQ0ayyQ
PiUhxzDXw+FcvOx36E1JgVHoqKRFE3bYaaqHv4vG1dXoFsaAhSuOpwCJTVW7iQK6
vgB9Buh411Qx4HkEFYFC8KVz7rG6E/D6gghh9uV6QXSfM5P1eXeqFhVMh+BJAYWr
Wv1H9JwyFfNXir5WJ9vw9tOzSUUPsVe8Zy94yA/hDwXgMwdXx/L4NHCZDeeexSij
7S10TQe2v4T+cCKwLGlEG3hSTnEwy1jruyCJdamW58++rCxrol5I+HAZjkgRh5Eb
I3xc/B7IvtXugXmNwq20oVYc/okomdUH2pS8SUwrMhu+d+8C4TtzfVqarA1NNGoR
rc31ec4C5xYjwGvYMvgRceUynvnZLUiuspYnBsBTTdOFvYaeaW+I4+U69nAC6+DV
aNFzoVtcCoCMmfKS9/zJkh8RzA4bE1kyCkztrw+1JhahSrdMqS2a9i4odEjPyFUZ
oAYkqcDWvYjRFU1ZsuHj5Fu2PoQ2uOP6v0XTvUdvW2+F1+PkK4I2nxuaNKgiYsGN
w5zWqnGP0jiXvPcmBcjSS9e4a1moDkKRFfA/Ar4K4Gdz81nCfQA7iZYFosHEhzrn
VVdXA69PE3mUS9ockY3FAPyJ4tU2nm5fZujWcikIMzK7YXF/io3gYuaTWf/7Rxd8
2qgHs6ywnPoKPziJEcsqekIKvFrQEXokuJS70sFgSmUBchsEOToVX4+T2gWZfXyl
1yPesvJfL6aln2YNz8OGdPB+/UmwQyftZF0X7ZOr/OLabIFxS0WkOAibgTQep7/F
bC5KXfZQST+6Bb/KUZDT8DfxA//X2Q2o5mgBRQwMbjyiZWit35enMlRUO/yd7xTc
NUGpTwidKun6SJFgwpKHoqKFGt1O/clg1jtQSMTkNttO5p92eb+7Qm7MaE4rqyFt
U2poFpn1eeEyrk2OVafukpXC0H0sadQMRi3YxbMkcttXAtSfcG4OQ2C1XoVwQrLP
asPFfP+PmHyxsMAkQqruD/4coOcuwlA4DssTuYkmYU/EfzeiZ4Yi5rk6jBLcAhS2
POkZe5NSUMWHTmSwRAnvxHDJp9UeyME5FPVthTEjpJGPDoVqZnPvV9ovL/m3KZxj
BuV7lqS82Of3tJLGFge81D3BrG6C0/sQDEfv28zoFZFej2izJ08UcVifL/9dNdTm
ZJAa2cuSBSi/arUM5YhDN4RrTLFXh0BsuAI4ScxPl+MeBhH5KCGnROfp81Rf6l+J
uSquQ52zxKzN4GFbc9t/zzbXaA2kqgVv9UzSzYAHDStE7CniKbriwWJA5+4C9VF7
IrQlc/GeX4WyBFntG0OuLXYoiQ/dk4onRkYqo4Kb073302q8LUk+RR0oiXeZawqw
MyiGHjksAFQudCdqKpFI58C27QbaDAqwEvbZ8+CVxWk2zUX75hAP5V0b15OSVS7e
Dxj/4AH4Ped8noHrFxHzD3JPCEK+Mr768i+tVUbhzLYNTXX6qDMWBJTsgaIXgBxP
OxRg7nIreNq0HoGXOZKE/G95gtPuqVApsagVeC8+btuwfxoEcdXVqjv3ASCooGy8
vDk6xYNTBlCJIjxNxlfDdWJ0DUCf5FRAJiE1BS9v00SKOjr8gtfQvMUy0Hi4BXwc
np4sUBMJooSlY+Hr3mhr6dWuYXMWB5d3t1w9RXRPSmWqAkgZhzzVjIKfJ6eqs/nw
wDkkNJMKivo/cSF/6OUaHJStcDQSM4QB3cHqwg9YMaMNaWIVg6qPz4rKxbMuEKXY
jNV60oOBWMDXgoE4aYeak8++naUZqqvlCy9CJqXS9yR/2YvfTvaZrkjsIT7QFOjU
6JBCAwiAEjoAQrtHwVxDpM5ne84v9RM3LfePDtTADQkgLUeql0ouKQqricR6/Bml
0b0o/2jZNsCx/zGseP7Jzff10Q+bLFRjg3hPThHKDpbPaQZUJA+aiCKyg3bsqAsz
gnEQdsZYPhZJYJ3sXjOmhzxu7UZIUg9FmR3hwLtfLO2DjwtA1I3CIxSiZH3+BpKa
5mF/jSeWjmfgX7rWOdKltVifp+vV03tLDJbFWEPRD5LUyKBWrVU/1emV6omS9lUD
KfbXy7BKJ33cAB5OtEIXs7lldD2LWLdrkk/WUMqSUZIYkeknmP1V+CQCJPtEnC4n
C6hOehNhmvB8Tw0o8wLLZJnb9kifF6enHYYklBGwzkw/c41LYEFLjaGcErcJJK1H
aWDv6qlm1sibtikVLsEDKg2VpNa/ctaNssgBq4tJ5Hznhh/u+cS/yT51N8dmXI0I
UHNsufGhq0+ilrwJRUs6RqVmBWpxM9uvmAxnkpzNBz5DeC7/4ElKjqEi2NesNwHN
CghJPvOiico32kERHsc4SiOSaS2oTdPDtpoZGers4/g7ka2inRZLJX87U02M2oyH
xK6iM0JeuSyW+hA6R+wj/MZ74qGqri+2JUyuHscZJCkrxrc8SWIVcBxBjPXNIEDf
x/GN52ekh2TJq5Li2JG1s+XDBJdCziZdLGccTksFtVdMkTm1LnySaF1df5ItlL09
NH7tUb1eEw8J1L8ZcaI05oDAOamM/po88VNNK57vNsNpl0niJuLCq81tyLvXXedk
mk93ax4G11Lziv689I6E9cK9JwNnRWaLbg/wbdoJLsGauELp2YkUevbzJ0t68KT3
fAAicruktkctRMVW9zhHVU6RXsOCufBVOm+mxIv68KtDfBPU+4nUH9UQ8Ioe0KRC
ew5DbcMdx7wbkC8zYKnj3+P8R3M7yXzQHnjLNiQacUjrn5o/GXroGcR+kgjVl7rs
iL7AnJbUh7X6Ur1OlE4AI1OFtOSjofn9MrK4oF5VwHepTHl3+Hl4lF7QSn72gS+2
hwFERE6jF7LawFk3Y/Hb50kz6Du5+eywUFcdwhMgasWjEBOsnel4NipWDRj5ZvJc
4g9t8QobBVzWd5eX98/OlyVBTdqT9izZcKTAozwjf9C27TczH/JIp08PkPr5zuFv
ojuNFI/7g4aDPiruHHSqd2NTS0Do+A8X3uWdhYB3O1sfQlc5Yfjq6LtXLpaLiGpN
HL25HbvITS5O3+YzTmUOP474DuKc1sZuUjCIj7CIJm7b0Dr2H1GNGLQJPr+1bB4n
Bid4GgpJiPzR/DMAD1+z6Bv79F3Pdz++Jyfhvq6pm2UAFSSj0cN2SYaGQ6zk03RN
SKHQ287SXGL3/7sces6vBjCdVAJ6DobyAIImD70mLT2oJ6+5MviMJzFl7pE63Ga9
4TtFYHBrOe62Zx6FezV5tG1rc85OcmcrG+Dwp9xYCLalBAbnUZqigVGo1SRqN1AZ
eCdGfPBxma95o+b+q4EFVqzo8DQ8GRmstV0sfb3sDzWkO5jFu2csh9GLhw/mkWcO
TfMPat8whzy0Q3ruPa4tF6Xt0XQYvVlZXhCNqTSh211iSVAOotjh1VeLdUVL//AQ
2xoSPdGqQ0WRo/pYLoD8NH9Exr4pOJpy1DTtaIUDYb2f+8NF4GEKYsWdG9Iynhgp
U2YXnzNEkC8ppdlH/2r7minX9xmFJjc0c7Y4mgSKLBFxf/xzTi5Y8l65lbGiJpVr
vR7dQrDn9DenITzs/6XCiH1MLfxk7dQXb2wKEcPDy1K4C/NeLQ+mr7rKbZCEyUOl
RkKMxJ4qy7mMmdqok9A9e/hwS6zIa3xBdp5/4Zps+9lQWDvK78EbkjNVDhdX8WjB
rD4IM6d1OXMdZKlflehMBfwpPTZBO2B+A3Zyo1eTtu5mwfP86d1/hXpYm6cfVfv+
6/mQZPE2ZBKugQq7wm5RNW0IynfIKit7WIL+hNUzLO4PK4J3Z/TetRA81tyupCz2
DWui7ge+TJaaLRvo2tShHiXtC4A4WDxTw1vbAnn4VWPbyY0DjWlThiQZitlNBV8g
BhSVaL8V2yMVNTdDiizQ24Q35ItgydyY49v7jrW55Z75cFPISAkF/NbtpUh9mw6X
SvPo9Jn8gY84OLumJxUrXOi8PEparx4YwnZoHOYkMDcqZLPocArHPz3KQ0W37/al
kNNODqkbDdpZUppprK1EH6cooCvaDGYKkJliJAzsaEOHL1ygOhRBPgL9ePFYJQwx
ooEztVq1063CYN57r2jyAH6fBbJSK7pQNeLHOh3JTgWimc90qphdka9Q/7oA3ibw
7ZHUQHnckqkJj6pa58fJg3W92PTyuyJ/i9VwowqKRWbxig5/+jlIroX9uSAslPmO
SLlbuW2S1YT1wazZf9fHBuqzsGkcmY186UM3VEslXDT0ctLC8cOLrlwZje3Cv13r
dE+FcfMpFPN9u9UHEIRBnRVKJP4M8W80dt50b9byAkIJ8zm5jl9a79NzXSVIikRc
NdwoQQYut7fkCT4ebg8o3uF4dLZeP3BcrH0IbpgNoHjUk0MaiBb8bFRqBhPs/GfN
2yvsA7QslHDm11MRoBDaaAV1hzpSLMzgLxvTLMm27loUqOifcNB/w8X1yrOdzml5
9HnUQA8aouLWiQhwhsas6eRDtGAtwhdePwTFDWYOvJzy+H74i3jV+6FBQUurRVsJ
z06nzApOTEcdzx4vBj2S9Ua0vG+27MhgVHj29dQXszB37/jYj94ng/UL1Yvnd9NO
GQCDGBk3wtlE53ftW2I/2Z1kZtqcLlrayYVEV5dXYLkGQHiHnxmXjhIrXFcT26rY
MqgMHvF5p5PAgzApdBdIHSDiUfx5P+CuZRL9KiTSgx3FG36qf8mtz4te3CTeM39h
G8NJgqPErldj/M0NHasMWdEIJiY9N2IFkBWm2Rr0voZ0VXtfo+QatTjviOHlBQ6N
c4zkXXO0soj7g8IwGmRVHMzhPW2w1uZ6IBvL1U96khVUOnFebGKulSYLfcYFVaT9
X7pQwGA0fbNuSIRklwG6+ZNtAznKUifQNmrZG7KaUyhFiP1+96iitk7A9DIp7BTw
9mgqsvJ05PAqE5kb+FQ7pFznYnk3McTM7WLchUP1jocSj6PAHx2xTqZotomo9X0l
LjzVqog/TwHMKfW71wWbAMm2B5fPID/KnBTVNFqbLbtAKQfXVPH5KDvoZSmvK59j
6uvppTWJ9YDhn6z4fniikTecrAoAmMTvX6ge6MQa5FiaimHQimIoMXUCIJUevO7F
BZRBwkKXq5lpt0VP1CTAyfWgU+SzgHk/nlKLR8r+G5pkXebWnJ/GM+Oy4PwPvHAL
l+goj6v8w+Uw48PQC236NomRhWKeL1VekX6vm/vXo5i8Lfr8M4tnNIcFnEAlpJyL
9VWYF+NItTd5UHkQMCNbkMmr9IFepOM/ctutVkhVm/gRciQu0B+tQ99rKW2dgWbk
Zyf0nUmZyK6tjLJxsTZnOeRYooFlX3ji9HzliaMRMZEN6mwKW4u/6uLUt8+EOtXH
Zh9z0yRxZ6uNPcXBIkjzc+JdeiHBpjSO/Ez4Hjdyeq1TK6dLcMRqymdo+E8mSV/s
8FuNQmUX5FoHaIzjChJC2t1R7Koggvz7mzhgQqQt0VbflZq7FyyQF+cM1YIPCJ/M
QV5K7Jnjsmo+9tWFARPyPURVx/sqK9CTVeDubmbBorcv+OWsgwtHhyty2q4RcGJ5
lZDpd0SeKKw6rjapCP86tiFHjdQ/PTj0Zq55W7hoe21u/6UpOv4QhpC7yCeeiBSQ
tsl5W3YMyyuyZ+z0zJnuZ6UIGUxpH81qtJayETeiTG+G7Dmmkd66z+XZ/IqE1Gq4
215/xkWTxEiljZGfr+PDHhLzGhWMQyonba9/SbFl1dhbo0/KVTJoEXr+0fO6RoE6
kwV2bslE/E3gXwUM/bkV/3WoiqCuO34covmAPOAk4RESXEE1GRs4KTWU1EIeRwuk
lKK4kJ7kgHa/3BZSn1gP1FkLX83rNH5iCwQzm+lqQ0zCi4kOuYC8PlXgu9zgiyaF
Ub4RjzxZYGBogrYMGf7/UvHJZu8+0akS/gvulm27OBiLinEcwYqVBwYYDA493YJB
0t9qykNlfi8qNEaxvg4CJQ8VWNWgRsh7UgrYQ4I0SUBx1sqAOSYt0MlNnoedTpSJ
bpIFxPloP0zwRuAPJNtXMqWAM20A7VwYNTwMyLoIaGslL3Yb68zyKhD8gOxuw69r
hxlSw+V2UKUWQkdjxVNNSbkxfhF+6C2LLwi/1Z36FpxFZgKyAqmxcrCZIdfhJoz3
y6KMtcBizzi6dbnpmcgyS+KxPb5Cg4JixsI2qeF6091+celuSstNgGRr2FQkxtQH
43XJCY4tXVja3BnbVFIC+0JP1d4UUfovnfQm9VPiIX4yonrqnEkKIDYY7we8NKHk
V8mFzdk7vaapHhm8wIuOoYodwlI+7Zri85Ad0yAGejHlcYd2oL93GcUWbVjzplBt
i8s4LVpV8lrdG5iytbSeIvgkx2XcyDCpZByBpoGFehKXtxYAHndZvxWVkpoxN8Uh
yLUG6IGhM3Vj1CGAjIocAKMvwaq+kzYOXSrRgK0ZOCT4I5C7A4JWN7TVStoG3kWQ
rfhfNePqnauaRj6ZjgU2xRoJkt/l45hWbeT3IJ9ig8c/Jm88oL0bVyBt969N0ydV
b6wv7ZwjYhlhGKLIg7HTnp8biys3SkHD2jGagRg7ZgT3cfocbzZHwfNvobTxuTI+
VGeUR5jJnfSAQTtRlDBxpqOuGlbf6/ts5Gf2kdSBUgYK4nh3wjDWSthKa3GJjh++
jvOSPaapCh48IwHhXNI6p8QVxX5nCjdB2FaXzIy7/oMGlJxPWe1ugNVcWGd4d6/r
uwhkUiTFTMG04EAU7R2VVZA36Q02g8CYsFk8LA7Ru9iZ2jCcTuXBAsHoZ1gzwdD2
SUEOe4PSqmScSvPh0rCZBnPVxXOIT1UmHGmbvJ8PWD4o/0NY70BURlQrPIWi/Zpf
09FNv+r5wnxO2WSsvHzDp974M67cX5z0juicxlGRP2c+2r0jPiITEuWwfD6hzzXQ
sMofMmFWgcZUZSa3NovAnr4ZCpZejeNYAI2YBerWFweuoequscQpQm20Ssdh+WQM
jM16M4hENNiTP+RIWD+ymvJIvonjaizeLZ7t8gdrfMl5xfB2qmfFtaYS+W80RW/l
el2FlDXSXA7t7S/dgwMS9cbTTWAUU83Wo8OHebNGIdYA6xIcrOib92kePitjp0N/
Xeste5ncK3/SO8vvayapt+zUhQV6ux5CCTMPxWQi2MCZK0PGqixnG5/F+ZT3aQRI
4WHbaDxSZVgRjLaruRwRQ0NXQN+hGHMsHJZxQpuYNMN+/GX3mxQtM8qBNQIPLbDo
GlK5Om6qjp4Vv1C4u6gBIxXmQ5mWhV3OW6s14d2QeNY0hbIykcWdsQFBAAvdbyYa
8Ph+o+Ibk2oWjPswfvUp49AsgWSbfnb/6KCTmif621Kw+PCZ9Zw0jX/CQsNffa7M
cToFPzKVK6UCwbaU5b//cb8lsVOYhogssHLHR6utpTCSeOVjLwNre/9vpQuhYOM1
UkzN5luZZGI7NF4SirqKlkJfHGaGg3+t+pYWNWdSLBTkBD4P8+HkyB12Gp2WXqHz
N/FQBvFHd84IYOlfXokil7llEffK9IQR2VMhCtzNodo92l3VgBaOBMcc84pTIA8n
u9uGS5pfs/6bBpkuh9s7h9qO/L3Ljy0aGbpNx3zCiIdxRK1o1iq4V7saZdU38bIX
f/ceR6aKygAHkXapFxhAgIdwSiOxI6Lq1xc8wJjZfrUq4+4jjh3RJ8bksWLU/IRc
3rgZc/YorSO4isFEYqPBi9h1sipMvY+fumgoLxrcQG2m0XbdT2Z319IFoSXhCMT/
sG1S2RzsAm8CHGcrI+esXTygGO1/nAggZ8EvzU/h3ZdT+lKOrAtcPIh8RFnbSSGF
xMT1EwUXZgeE/ZkxC9nN0a3TCDRSkF+w7seBeYHW+CXnQn2gZncBJT3n6vKBUt60
9rd4TT6Vr9O5l/5sFAOxHTLoAATXG8VKTg+TOr1OwmB2hHbdbk2r6V5xjAVrpzCN
qRuubl0BYlqgdobnPG1wzctRCnJcfy8v8eJI8rWr/vBGBrZp0HUEoPTHH9jPynLo
i4HX+rF/emA5aqGUCPh4SuYZac2AZhZNb2ugR+fYXJeY8FMCvTAcajnrR9Wn2AeZ
KMLEY1KXDWo++VUucp0KqT9JFCuTIHmPg8O2t5omIs5D1ZNoQc7hrbX+//eTwSdw
tJFDSDgaScQ9a4SNVqFefcfKFwgpgHgLp0AUZRT7uqFdo2s0Nw5bW9udyDgD/D3q
FMQ4z/NXUL+hDw/cWicexRe959rkWNorNOQI8JrETHkUmkXf0qhUXWO+8Bi2SnAZ
TOyGkrUvxA/JywwrZe4gTvnq5GZ8nmk6oA1Kp0xjFeKHsxcsj+AF1pZIaBjXeys5
zlHwJgoPgc2c2hYcxhP5RMAdGBCR8tH2EXeNPNA/UrUyGpoaxeXYOYYhssC4eUZr
nnkw3Jo83Vk3kiL0twSuEo8ZxdknTp/RiZG6JRAtSAOFIMlkB2AxRdz8H0PrkLmT
9zxKOsQ07MXo4RZtjusoG/EOMIV6i0vAtyJPupjt/Rj3+dpS89qMz47RRt5ei+fc
+J9qoenDwjmfPDEPoaZP6+jVeeUHJxg0ftN/vD45cQX5AJ8T4sdo22Y4awxuMZcE
PhtobQYoM3LZ+EbkSs99M/O9hSkKuG18rpD4Xip+tACoohp/E/N6Lxm/ky2bv/ha
yBF3iGDvNp7q/jaBGrcXO/b1kS4QVlzEAAQN0r/B0gyj71SKY579bOyTt69NDEVU
97LVzA9Vl19ni8ytiY1j/1zR5oIR3EoIqJ7cH0j+efoalNFIYdoOCMVtqzbSq8Hg
t+J8qEcEJfV9UDBjqd93fsVqYsllgbFROwwT96GBo5X9x8rkoEH3wRJX5PzYo3jy
dgl09Wg1Hxf38Jp3UtlnBtp0Tdn0wxQMh9eyG0xSlL9xZWCRyngF2veet9z4jQFd
MDIh+miY+ibv3Pms9YK+CeBWu2l3agmnrsbgrZ1l98u1YvV5rwsQAFPO8o4EbL6h
NEPFnYnDz/3nZUPmzz9BlNKjNYFjsndAk6alVSlOtDVMAJzVmAgsNFDrjA+Wt6BU
oTMN7X8+8njloxrIgElIp0l+neeE6vuih6kst1e3E+Izz2ZwUvy0HC6Kzk5kBauJ
26vZJgrDAG9aJkfRhOYd667oydhgBNRbmMs34s222ONztzaTvHsOJWiPbmmi9C4S
VjyCWfFiT8RSBS4s2dzXb5YtcVKqc3Oqxnl+eq61qxYEzSNRhcWEamXkRWBAYMio
chSmxlbZHeGaoAyI9JddsJ4eVTsLD5ZY9U5qJnOk4Lwvr+u/uzIW1RykLz13LdN8
ZDtQJ6Ah/x3OEvlX8WubgKZmJgIapqiC657LZmyMmpDziMal4Afiwd61PiBTAnXO
4fDBpdGDvuWJ+jmvC8AcSdiD2NJuJCHXewPFpRaJ4S19pMgWi3qfu00mHgDtZxUR
lXf9VqDos6AVnl0fprxz9Ab4EL4DZjmZkZK5rhQRQFvXUL1lXSOZOqec/7HKrJ2y
AzdPc34/hzdPFMtUFwRrRmiWXzWsBn1fk4JOgCjmdCnp/xEMzzE2+gfvjwzsp55E
8EaXj8BYatGRJjYUUoxhYSPzHkMP4mLrB9Xlf61E/5ZbEpmKUS6YkYrKhUllFMPq
rJyTkKd3BYXkES5MW7Z6pXQn4behKf6+RneC8BIdhnYdKOILQay1Y9EMrM96J9KP
umhIJa6DzlZc4yzVU7q9Mp4oiUIDHg05mjE5iVWXCN+VTXxvlx758mgSnXWkBfeu
A5VikUiZtGMmHu+KZt3CsaJzDhDb/jEBM1jtQ2eoOaJa5chBeYaQNHOBH9Yr/56V
iCK642Cyssa8LLg8OJosMb366CqUCqnfEiSARGaAp18d9yQYQX1taIbBiVW/M7nk
6niUdaF++0mQ7dVlJABHPt1vnw1kJPHvvKiyiRO82Cvm3gY8trFtPZ8+nPck68JI
a617fYtskS2VwH7CmSspLkMjiXyWNr5dOscNnAsidbpGNodx5Ox/iFRwRPkaISWX
oCpOId1mUPN1nLPPR93sCEpmqCY0Tm7AR9YJRSOXjRQoOekH+rVjUkSAyUK9flkR
x5X+Xl6kpwhZgGsQRlz8VO8p4iH8OmS2Lud8/a7yui/3AOXnvSQHGNHgwhSGEzod
xZXQA1Kdhva2Ko/lpHaNSUlHyKEGSVohs4RW06lVMPftHD2/rZV98ivELvTuFtuz
WfKhoOCim3cjrLcMEITbCu4eFDuLjqS0ulRvbUnZJiWMlPFCjuo8p2RvZ94Kukk4
7Ff8wp1H9Ac5BKGN3m5CIukYj4CJ6NHf+aFLu1wCE9fhRNhQ6CrdHHt1xc93xHt8
7LbnX94lXDMTQ0liLqtTEFac9iN8/b5XWLf1j31se8PDlKU2Xj1O7le+qyKB1lGL
/ShCvxumP6X4O7VXF3+zkOpJzOXVyExWpBk+O3F03kFMkvMw77NsdIiTI+Sxn7uW
eJiAbv1ab7Drra/+x/G1zNrah3uNOQWz+wO4vj/jkxGBYCy0mTLkTgYpNE+tExDU
RbYC8PzS5jiDc6kKK45TlJa2nBQ9uUTd+aWJk2L5lHxXVHaZTW3cLylrB+nWfPve
Q+zQqIOvWTuM1KpLrPPW7s6vGLT8hHRc2y5Qo8ta0I4Cj08QgZipypanJklEoJ0O
ePsoWodVY43wS7PJRbH8q91+ufUSqDe3JNT0UvnVWRuAfnJZpTIc5wETTvaXmMXU
7BpL+Tr0Wk+HCzLsFJNGQtYwyzN0++j3TLRmV7OTB91YhvhE94Cxr3H1CR8+CUNa
xOw1H4l9gT641edc+Svb2aPAZErwjquUSKuzrgc4QY5LQmw0A308qGOomdvUl6Bn
CExwHjV45tf0BYcJ5NimAaqTupMZE4cP07bXDKbuJigEoToyTt7dprR4pfjSr/oa
iLWv6loOr4TstduhnqAT58uf5oAoFr6JNriOQNe2A987eTwN+LavP9iURU5de13u
R66ZnH0k+lZ9EX2vrJKm3r0yhN9H/p3Euw++rWt97RlvzXljWOA3D/LcmTh404IJ
OqTCPeQUpmU3fQ7DW+QJDHKCd2nLhHw4SJUD9QDBwFA+qKULQj4zyUoGKCIdNpoP
6zckv/YfjCyYPzm+KXnXILUZJcjJPdSYUwuGpOyljEB0bjJBUGOTN6qPPU3JCh/O
nDidmDpgvAV1d49674r4RaFbX/4LF1PKomej33bOJ0iGX6IbGcwsobo7EfPLi7+8
9saZoeFq8c/zZpnEesoUncm9njRZ4gq1KMFCV5A5lCZQUxQSZsU04iZNjNL40JWH
Nni7YB/JpPUtTrWheQ5Pf8MuuhomhA+9Dk+ee/QQUTXwxyLQdW2PDh1n0eFGlVDT
LMMHHu2SFjlke69blc9s4lkB26/P1H5yi/azSm0ECZpV6SgKLIZHddUqYlac5RMj
SGhdaCGtpC8hOx3WZnvPxrekboCJhfe6H3zMnfAPr7r17bwGN0hhCHKfVCE4USJM
VzmLiXP05J3t5e/Tx1MxTQzAxkyPdVYZdPJNzeCRmuwIPRACD0GohF8iE+pDElF0
GDRWyoXJzNjdjrwx9YLLc0PjcW8ZCywj+h6+IqpAk5bMGg14zeH/3rfVOq4xhppC
1SHt3WcmGIfymMoazpLiPhuoZHzOFmjuG9om+DftD6ujmc2FrsVE0g1vRuGtvmNL
eKDVJ7zWfIAq/zzfhxnXMSZ9ebMUHj3Mq0fNsisb4w/xzkqXNZbt/P7LDUQB3rO6
qY6cFLzMhz2XUGB9vV61SvaHptB/DwA3aspk/J/hVwhz0HyOLG8YhOAMe41ww3PQ
KNCjueiHcVs9Np7sb8fd84e6eMrF+QvCCwoe4Vp0Yun+3n9AHLlvZ4SuJxw+Oz6g
jn0jO3H7vEQ/RjOiGny9+CbmyTpclkwmWhSCHgAMrBIcjDgKWT7Fdq6uN4U46jFo
xP+/6ktEhw0IHeavpVUo5z6KLDjX8FDg3MhWVri6+KFjXbqD9z8j0HAT5udTkWST
V2/TdLQvwniNoOZQEVQYw1c35+aFOtA9wQB+3b023hPFG6xGCmB2S8FlhuiskIGg
cq0ztWEUEy4B2YF2/Tq+3oxVcfPCdEY8MgANS3YuCndYJ3nXJbyca1NzXlIQntUy
mhIXuTgA34HrBDfEf0eZXl8XJlwiFN905dppboDCpHMtBs31Z8cRqFAPr4pXQyA8
Fii7+4wYY4KKqdIAId/NU0Ie0ihd0QTKGsf/Wp+nxA2yZkGCSMUVE0nShpPMY9Ef
SYFAhaV6rslofKkTkiBd5FoMuxpLovENgX5jDtN6jfoogL6KbsrIYNzQAdbD1Uzl
r/vwjDwcd98v5x9c7CP8mz0XQuTkDXxZJ+gS4X1euRsT0qIjSixVYSjEXmzJspL5
C8OsgrnWjymDeQhzqbfBC02iMzLzqrM1znp4jI7EaK03ZwaM5FNerTE/5WJPJGqz
dPWEHQ86mWEHrJkxf9e+ipY5VQ/sCsP6/6OsjBgsJlP2FE6xCvyCHnAgJ/DQf7mZ
DdJ5bPPHrUsOnuTy2GzcEUoy8vT4gTvih7RQYFrTAcA/90ws12ukFm2qdqLQ/aRl
uAK7Xi841KVDrHg3lvlYbz/69QeW54BM2NOdHLV4O2FAflWsFF0wYpevQhx2DIyz
DJl55mp0FVHfq7rpWSKs9mTSmKWTyEYlUPbvWmQdTc0YPAcBbNydeuJG5MokdgcL
dm0vwgEoOJQlZDrStgbRrN1+k7uYrELuuk2Jt9V9YEiGDkBIKQM7ZwxC1bSm+mt5
E/WP/IjESGmpqXid9G92SuJwnKsXQ1tF5MxAmspZZyxrDgQ13Bsq4LL0DQChFR+x
VIltWNB3B3PufgXu01RRgxSP86dkd/fkqVqeB0X0+k8s/bAWFAVl+mk6tdNhvknz
GCRGoMMS2WmNL/pMu3tndiXLg+io3HrCapg0y9v6Qtmtu77UU/sr3Z7Da+L/Wiak
el6Lbo3Y6c+vGLbrfkn2N3K/nN2bvfeZMPyCoTfuvcaNp+HHdy8IdkNmM0bUbb7h
br39jP+lmjTw6b+d4iCzEXZ04AbTcm16zIdUFktPglxbLMyMPQ5fNGeJQAa6ud0L
HfmlIBhoInx2jbbq/omN/5yBEKfK118rHkVYjOE4tSPj8HfjMsI00IZuVWvMk6lA
/1UWHp40yy8+QS1fEUKaHYouZU8gM2zKh70Lt2YALNvY996KlgCaFc0DuVbkq5Ts
qOJ767W78MO2D7E63vyaaK9GuqVs7KzPKq6pS4uQM2f1AgIvtAhzbT94uRbE+x0l
6rv7IFnPZueoM1xSihEJQBv95utW63Qom6sc17nS4C19K1eHFFKVc/eUtXOqu3t1
hx3m3xZjNA/nwZcfH8NH+2MY7Vgs0C5b3ZNApOkarEQ3/xAX75/K7QvKGC8qqT9C
2qy2pLMRkNvB84of1EaL1PtRmvSsl7+wVK7gt/CMrdw9aOSWYEHs1KAUMo+c4OOC
I6z6bDVYxhjSqzZn43eq4fQoE8BMeEHR+fo6JfnyFgOsg6Kha7FOXldkjzTIlLUb
aVmtV1T2xFdUKsTCSsZaM9kEP0BNUz7w8iZMwQeuFzAt9pYEPw9dCPyEIk+LQpzi
260iw9SmPGzF6/u6X9P+UGK2U2JfBj4gLZ+Rwa/uQKL/Ca62QjVrpbexA20ysv+I
YtCB8zAJVTxqPAi9YIxItT8MLFEdH5Fq6ADa5Qz6mjLC6MRBdi5CZXg4Mft2gC88
xmD4+4d4MYvABOSlGTlZrTTO1JhvyAOTVdRR34w089ImPCorDhVB4a22Roa7LgNx
oxd6Y/2EfZnuxEmqZh+1L2hlZAuRdo2MsigDUpjx1G3w6PrBkeuyTfzs5V0s8wx+
vLYWRBsspq3Vtv69hmRR86tbgKSSY4+sS7S/zGM5lFf+kMIhN1iiljjJQIJeR4PS
DOwUxcAU/jKL8+ckJi5HnIHw2JC6bbB3cVGtJ6tS72jtjKUwrkwBBDDxQEA+i+PD
SBtGgD95+qPkxyGcnN1HzfbRyi+dJTrtw3o96yGiHK/QIi44MEkGp9sWHEVSmWHC
bmDhVOthBHt0Gdu9p+/LL6T7kVXnN+BLxmNu6RZsqrZRFqtVdxjn2sSvKA5oJxfP
ec5BsQMUCRvBzywB6SN6CGJW00/xhEQ2pJGwdzQzYQyafc7dpDDaJ8RDHMg0r+nT
232IxIyTbWj6vtZs1UqU0QvorY2aP+lCfIAFzs2s42R0nX157p8W26YD70tyxoez
tFv/70cQfidqQxHu9nOzXMeuDmVV7rUsvC4EJ2rU5MZB6X6n1yKcd/O2opWb/C++
dAJNd9UsSldD6vp8uzT6nLyMnVRgt65UE/YQj3d1hDAdGuFoq3KTBTrPFgzIB+Lw
pioZDcGBxLaxHaYWwz+ah8rsFXDuV4HK4ljaeoGxrfJUl6TwH38c3bE8TLKGERFw
4LHPrJPahno4rntKM6WdY/+KXtBhUINQP1g3/tj55CDUV4aMqi/KG2Lfo0sqFJIB
vx4Dq+VS5bC7fKVSSG0DdOXV+4UrO4HbQqXi7mvsNqB7W8vVNa8xmbV7ETayxz7R
hAI8Kj644pZSMDN1Gl3WYRSHkIykQ8HP81XnkuvfR20UtBOBphCYvadEkYTWjTnH
fnaspW3x0DGuyQQYxiFOGaSrImSNEbOu5kgT79WV2LiB+GWUstNKK78SarQl5rfY
yPJNADoP3tpl55BFD8R/a+LJStN2zb7JiTLBrR+OM47e7XeSlvUzaZwZLeHUjAeA
dSX0hnNbZ0nagjR7oV9Su5ABSB0NSJorO+EDoNZ/Bq0sYMAruE86aLOelEXuZIgD
eSIxZLiGNEwq3PAbrPxRl9QdEPtbkAqe1zi3Jk8JPDE67YWqiqzElOhm0uw7qZIM
JReJWzv4kFo0TEaK3RqbMKXnYsfYjlPZyvPz59GfWvyGfT9eJhdwrUPYBAwVZXhf
p2Ag2ADKi8wcWPA3OhhLIb0R+2tw9INK6LdZpdeU3Zu7AcHImZ2tfELroggfBWtT
qBAgEYhLd9ewnaA9ZlTEg256dmhzcJzqaPXJK3PN5HMvKbjwCbIGbvKsfNwIypUx
YXpYKi3Qse1Gr5EWqDvPGdE6EFNa/nI2qZIj8TxJAXnm/f/73lPqwmydWCggcYm6
U6B0U6JcEv1H1hB0I+e/+IdzcsiIF7oXCH1DZxOcsXj0odSsHfyF+XOxBo9oaJyd
awr9HAN05J1lEFn/0ibJa7W+FZyS25cJEcq04X9B3XrzwaF5hqmuWlHoxDc+KKaO
x5V3xzMqcNPrG2VBUGNSAZ+tW1caD9/Y33IckStHWGtgmmPiAuVbqs74r5qXrCLE
rL9fvBbP1DR+iBr+x3D6E0ylbyeXezt9xS1zqE46y7HqXPUtAML4P3TFQS7FERPy
wPkzxL5speiw3Cu3amWw/pSzIGMk/ns3lD0UZ53p6c6UlEQtuplGVsZ2gNiX3Zqp
1D9mX9grH80nmZtciZy/XBGd99gk7Qx5HfBt5DkNfjxPRS7Xo9bFPzvhFSfeCKmX
XCwHrmbRFhyrgt7sxVHA7hHWiLDJzDUVKP23VigmauSmJRVTDgty0xp3c0I9QuwC
nHVQY47mxE6cUyvLiNqtkEzquoxMUhHp3oW0/ZnyK3g0c+WVW9T1IIFPcq96XcSi
JDjTi69En23xDIFL0Zzx8EGfLOZ0OSd20ISZpb9m7PgGfuvtrnGgqt2+q8KwfKQX
1sdj7SjyzQBcLZTZScZDbVI6MVcoigrM3U53kZuYRRk0IfrngSmasOHLPYwsrHuR
E2mA30HJbZ/Typt8hoXt0+Hdpf6Ny1VzL8ehy5WMxyYop+n+Z1N6FgNzKllyhWPX
HTFpzw/0DnU/+dSNzeeZK1sN7tdyImJWOpKSYKZNog7IQnzbprq8gQv5nQ1z0ctR
jxJROPOzfc2W2Q2RJTwAOvulG65VosnAASm+/Z3PNWq+kxWPbgFnx7xGkR8siYuJ
Ubi6qrvA7kd2cXKsyuYZXoOEnecgi45pombV3MDxVOXGR0fOAKFMgyT/mURvgpCA
kR63PloVHsnfZYXAOV+kxjkXCtR06aTR05ejHtS/aL7X6y3NJqNfdfhKIFuerbu0
ir8voABb77EecHa9lPj8jC731dMueWIKdADAa+1qrHl5wF/Hca9hz7q27y2ceCR/
Z3R4+CBAEUj3OgmAMTMcTO71ebdyktuTUA2DAmJw+CpJP9bTwNInrapgF0GR58ey
zv0AqMb7rDePHTn6I0IuMew9avcCSsbhgxLff/d2u5Stbw18BL1U69UCyp2vU7HJ
6iTw29vK/enKP5vhcGr8oUBnyFI145Hif0LdqB3Qm6J7FHQnSx8jyZ60uWQQq3OO
primEDRlyfdYPphWQqQzOGZBvA3Jz3mBehKZTk6MHhkiPQiDR1lxJljw8t98/98b
AbJ3xxpiX66zr4EvZsWdKltPSq2xCzgPdgpVD8UM6/U/nsxOxRNNS3O8/F+NLmj0
sRfj+aBgYnAT5CfoMkp1UqaT/QuLncMo6E7oLVgtGUDhm6u/9u7Q8RaQzGHRakpv
DlC90U/JgfZSQiD477xxBXJV5XUw1ByLpWWl9kG+/9VowIaWjppUm66Ruld/ddCF
Dj1qYSRX+3go/cBi4um9tAvZE0kQmhMbUFyyG1lxFTeJ1oaCOaMkCWeQwqphWnP9
FPRTvYrH8NV5AfdDC3I+1+UByJFxpaSrdf1sPjFUGyE/vVhzXivZvJezg1o/LTIX
xvR+RNepTlCM/n1HO8lH331krBw6Zjse9XkWO/mqcpGS+45U02Gi2JIp5lHlCaaF
u5Q5wPnYmOiO4NJnvJUYuaJ5prGnIfljFS4srPQbkfXDyosOwB+WIq0zc4GZzIZT
KLETG27GXRd9SzP8LDF7bXrfMTYCDnaf2ZNlLXnZf04HJ67wV67S/ESWNAn34/zR
cuuJDq8RRSjfQUrcIwS9SSwiqU4byPpwxNcgPHRfi6Swi7Cy+EH+lXvUx1j04F+I
L6dn7gEhpmupmTkTwg9yivVYR8Ks2AXwu0eaAzi39+lFskyXkrdBjBnwT2eJbhDJ
NENt6LvE2/iiXzmRQHfPPY0j7PmU5FiBz2CPkDfztB4fZzc3uYrdjeIp4mtDshJ2
Yk81O2FRppUwE81nsgL+toCrl6NL3K06Y8mJmVkfOY8ENPKuFu/shB1ltgaU3Cuh
q4lVbblZfhCct1k5HabdxCRNd4HAwEmTKDcwUVkytawNc4rjSIguq4bR1ZqTUd6z
OGzV6xoIGb69nRi+QxFux7PFq0w0L1XeEPCVvxIVErdpK4IkUrtJmzFWXF1xNZj+
dNTrbKQlV58LAGp/dtk4CoZbfZTayFpl5ADW5DomcIwsYvf/vGWqs1mrvttVXW3D
QvJPevK1uPusft/cv8yIAn/sQtYU7+0S0trziuEtMfmQtqNDV7z932m50lVSt9YL
PfEJ/4HkAlKuk+QU3C8sEQUsluGge5DFI1PlC7tQnR10yCWaAtFYkqNGgyqd7N8l
FkwHLSj57DEYMMtGP4Z+aql80LcWcAuQxC12/DyJrlguGA2P16qelp1ErHezQfAP
HSTouwyPmD4d8Vvr0vxOXB62jtq4ZzMeaz2VGycyQn39x94zO6GGPIAPGgKJvOon
W9fvRqktvuVLwQHT6lS8LVV/vKkEk1zy01CsnSnv8vKX4kmvYL9YLsFpN8UZphnV
7c78Q8jraUP0l5G3h3gANE2t5GgkMLtMgVUk4QZSlFNetw+R4VsxcnTl6fHdlb7U
KVHZV2MN6mHxJEcAAKYLF4a8JUQVHHYsuP2i4rY/YRatQiDSSTyS/wlJ/R6DHKsC
9njcL/FBvzgBc/uWNsvWV7DnfRyyuA8vhaVykjrHmbzFS8V3kmQwDFTR05XpovXd
8sEOvwSNR94a4oKABSMjjfDP4rkNirs27Ti2QgGd19gAzuQhg1jGaHnfLOIrj8gH
q44v3q6cptpjTf1s8CJHXnfc4nh9syr2QOHVO0H9sMRf2SATCzNF02y169EfCTpp
ibjLkA+2SpYLZ/L6UFuyGvCwXOfYHcvhoXJA+bX0Gys+cvuv/S0WXox+Iev5uKCt
4pqN8ed6e5LVQ8Nk5C4YxPCIV9o+ZM/Go0MQ4cNqeQzgFpo9ZpNf1v7hEpgqa5hN
0O/QVcPwd5ySLtkJ8jA9IwXXp5Xtxuxw2NN3sqMKKvpEcIjpLpYCc7AC2ja3ukEE
4IG7MWcBQmWKhf2Zb4gYVS30vCmLZLqPETV1Zi9kxS6qDI/rQvOt7wNeIj9q1sCa
Pdu7/IXfZs7yZrylfF+DQosRgPlcTcvva5qQ2XvxQuMJHDsH1+E0rQR18Fkf8pij
skyhOYIWkfN8d5Yf/a4nDk4r4eGDBTFA0uphUuoNwDkiy1cgCs28wJXNmHquGQ0Q
qDWbKL22cWccXvZfGQ8hshfMRO+kHnQJ6IfqbUxbFw9429nVUYDQ5neeBTQ0cS+s
7WRn2YB0wADa8zJ+p8vH1cNohX/xzHXrDSaGsSts5XN47XsAGzQb8aSkkwBbmPHQ
D0xyFhdbPIe5O0UnX3yzqCYTdSawNfRqiHsdRWb+T3/nZCwv7zdjNHLbpm+fmGKO
fv0ViGPubuqSURPGhIjxc/RWOPj6gslD4LS/a1/pjHav+W0mZfnuQiftDbfvShRp
pncxtz7ACSi5bYDGPMsQPcsORG38/qxjc6BjBlmc8+nS2K9c+QU74qnFgSf+KYto
8NJqkuu0Vxt3DhVh56q2aeekLgLKYuR6nWYx22ovayX8/142zdRcb0y3DVFuL70i
mpWmuwn0xO3HqVPxkmiyO6+0XsDWy7JE6HH/MoowcFw1y+pHOB5QZ0Qvw+pLUWoF
2QsOSCB9wsj9TFszBfJi78vz6puYMpF5z83E+UJY6c18C968l6MJ/G6HrdhE9wjf
i61EutF9d010G9KVOBMFsAJokJrVS2P7Z9ybAwHis9lYmsaL2IKQqZtK+mIxlEM1
Kfm1vKbSOaMZuS1Dhipdw5aAcrCdxAtXlGHn37s9woia9oEZjWUy2mphueHKghVn
plLCDj1Urw2H4uH7oWDqVr7E1Jj2tIM6Jj9OlErzMZ5bz7UxRTxHEbXcwuXcYBE4
/EwVTgg++1gKFf/n9+5eqXF8uXpxuwYWf7TN1jaskM5OOkxKCa6qZku/ljQ0wkDh
OvtRhTfdD+IHq3tRwkT9bOTZjzSC835wuwJktCniYPJSiVXduIKSWSfaTcQ+pQfg
xGsD5W5EcjNXFBVRJnJkF0okyHQ0gpJ/bpxW0lhm5PEudpoYBvNNtvMrz51Ic4NI
uZu+i1qMQtB8Jjn8TOsLK5ftNzFkYSzyzcr/TOLvVe9tzxvl1TAq+Z45cuJTpyOO
Ro+0i/zEHSbS90BWWnKGqsVd5rCtH9YvNkMo6krHPXj4shrWNinn5s62zymEJSMl
jgIEq1M2Qlx5jGAs15zOXNqTh8PRDmtIgZEPxWJNG/2CGW941QJSuKaeJkjmtVca
lo9OAxkXeVTMiqTxCLlUBQto1pbcZtXaMrPt+9zTvsgdAcToi8M8j9+sEzrWYNyJ
0pYe6FUxW27VhPIXJvYc1U3WnkOVdYuay+BbwkylA5/XpDF9NpI6zWn1dOnT4L6a
q5AXz1rl3hGTLoDTTxkEX4up/gVIU1n99yXARK9vkIGsdaqbaol6DzklefGQzYIL
p+kRUYLDN5AgCPn/oAYW2Ayun59DY4IbELl4tbJQCKBZ9dIWdyzgSUxsIcMNbCT4
caUsOVRWTDozYQhel/LAhKJ9EANtEW8QHkjhMb9OXRyILmgVaIiQjbnErPB5emu0
z82C1QVCezLYfWUVJD0Hi+3GOLmlXOZZLZO9mEGEJANPu8FYriRceIfJRKF+W1i0
DYyq9wTwN7dMSjA4JXGZHoZnv/HdHR8bZOiCGR1c2eHGFYwAjhnDHfuqSFGn16DF
nKg9xvw7rTatW/am221oLJZehz2FZxoQ1JqL4DbIUlNPv/EZBzJvr2egGvTwxGaf
93pJkw2QjkK5O1RXrUxX28AWNK0OCbnawAuEfw39WneyshYzrKzqntV/FkGrJwZz
V3mje3bo5FOr5g25STkslarg4z6Ts/5OVrrduiewMtcFfXLKQwtgQ0dvNlgzBBqU
6JgrQvUa/e5cTmEzSdOhP2Bq1EPZ01qSY/NM6+n8OQF7tHZ4mqUf1oAwUMYkevPV
1KTGKgCgtsKfh1CGfkDP7LO3HMPJXkn2KZ0cvaL+eNEI+oDQ1ScAQ6adHql3YCUC
fVw4xrDUv6SaTq3PoGuKJQr5tUPsdSo6xmmq5TxNv9VFjPl2AkA40CVLFGYlQuVR
MBYekVfA+vadDUvZ26lwQ9gbNzLvKsP4zqCdnsTX43qFfmKkLw1OtIODwVBKFG8N
2ee25IubR96nkXgVhbU4jGkKJoop8GLushne2Iz6uIiMJptgBrVBtcDK/ndlSLQn
X6trzBEoNolyDedNuQ4RVakOaVG5hVuKWJ6Lk4vrw+E8jTsJFMt1WULB/TNQaQOU
vubVY11jSD0/rktFpbggHhJ8B0f1t9CXSmUKiFE/b5qeLG2ELYG8dPEChitXmaN9
ep0VzqYaJiqj9PJjSSoHO2bKFcgvMySM0OY3i/z7rY/QgjPPqGUrVlfAC6s5SQ7B
oYWzwK/4Swg+egMtWjDJTJVo+/KxTVQNJl7MDpfqPOpYsSXvK/2egYIb4bz8SbJF
4d1ebu6FdvHSO6OSjpn4oePPzRXUHfo5uHCEr8V3YjwY1H39IhzW4nEfv+E39TLA
Tkh4Au4mBYs6G8EOC8p62EzMQLPCIubPWp7D3uMYbbcezI8YDXPDQhEs3d+JgYpz
JiUdp1ueomi9ISSTOK4vfkq+HMmf2Mxeqe20elRUX6Yel7VCGdUJx3p482h3yPJ0
Xw4Ij3pwR1tAc1Z6oPEe3Us2w60vL72LMZAUmwoiTKAVLc6WhluAjCl87Ytyv4AQ
czMzcRExGIu1jF8B9ot1zJvFfPqHLPI0VyqU/C+94dW8gBjrqNaq6IOVCLZXjRhU
1Hisild+Zz3n9LI/jo+ZcLcddWQS3DFDAl0XfyOoz7zjWa/vlCsfQrQfCwgr4TqM
Vlo+QqJl+1gByMdSxC3Til8u8SNuPT4jsbJqDouSn3UARC6UeSJikzmo3OiUoYUz
L99SGpWxbU9Qjeg3vtbyqzC3xPxqESKoS6vQQYXtsWeoUyiez8sLnlWBK5X4iy+p
lGtxgAiy0k1wf8U/qMB9HCzfdOfmmhPUc0+J3gwGz0+vG1rYo/tJ6zhoUsi5WRLM
GAtrX2xvdjsItmo8H1j4MBqeexvfHu91BRvu2d7n9c7Eb6Btm2viw3evgbeNTCqg
d/OMyeQ9yAEFMdi0of0PskHlJ1gjfW4LN1YdUktjU/hPs1ZvBc1PfO+csnW1AlXk
tZG5LKFGiN1aC88H8mjKuSloXHOVY3GWs48F0PqvrYDi863P2vZblf2ltfWF/T4V
4jyp5En0VbUqDSsVaHSUozmsQKxWPkUCdFlbQikKjCZLFivGbG5YnKdO54OOy/8v
REq2OgXroJAUv8+gCg4UKAnw5NhaujTvUC3Um+ae2N8NvKGJJ7e2WvHwS/d86l/r
wU/ZSWTHpuiYrid4+OWiP2lPfhubILhvr51KIJH1Tv8PYEcft7+ewklMH0ecmy8v
k125JfE35Qth7Nx0bawi9NB+yHMe/Z+NHYJPdCSAKKC2etTNTzQEKr5Cy7uLZjjz
KIX9LwC5cY4JAidk0GciljJPpHgMQ2wlQZaUnTmofYWH4tWb4+baaNNVmo0C464e
qh/Y8sxtYdVu2S7O72jbtucHDcM1u0sXU3T+BR4vMFe6vcZrhJ6VrQhJ4BIB0+hk
oXTpdJ7cq3ET8eHc0t+wJj36FPybibHebojM7mXPkyjj70uSd5htnA+/R68jbB8J
M1J6iF4RgeReHpSTe9KQ47hSjukxAk0WSqApfyW0J6BkRjg6djBetPFSIT6InYo5
EBSZ+ZDvv/ky/z7H2guKb1NdKhw2c/h67tBVFmHPTlfi/xUBgRmelFEfcX5JBdvL
xbFswqnq1RXvoWxIoSzY6jv0kWPK4NNyODjyfx/C8IUCYKrJWd9wIL7MJrDSlkVg
hgLRVp9jKrh5ulUeNnRWdMNj+oMVjHtPzOCTUyFC0KYIEp379hhnC+VYEVOduhyk
JRxFaLWFN8ejcJiwXANLmASrDPsPQoDxBK/vwgPdD+GSUa03Wwvhs6Ijk9eJsVQE
Et/sEpDYeerZ+eGR2VU5VR/+0ZYgnNsJaDhfrnq/NFzwOHw4z+IrZxvDimrG/86R
vruqpZcewyJKUUyMvYklboWF/kv6nhRN0Cz7PEc7FHe4ki4kSor+2/7vidDuZXgY
CBzHQO1CyKLclFQyxK439zgZAozdlinzp/vxQ5cqtRdBk+xzvDgH+ctsU+Wo6GI/
TEqupAVhez0JDU9oLJ71q80h1GQlg8wyFM0LWYH7V8xcH9UYxJv++XOaz2nxS1tB
E8eFsfR+J9W7e1AQ7SFK1Iz6YCgknVxKd68qjLAf4Uxa6JMAZzINjwwYt1CRB9yL
2pRX67CqeZsMNEd0NYIlaEY4TLuPYYvNv8I/okwh/x2WCLh/cRybyp0CHeqMJ7nW
stMvZuVn5sA8U/QnRraoPX6mXm7RukCZqwUfgx24u2oV1J16QsblB0yrk4sw3wpQ
p5NDJuVOSOix4cdr/MJ3g7YKs/8i+9cxqFYMsCeP2f0xBwwgN0KuZXbXW6xDzy42
Rl+4Hppu4mc6rmcNkjCI3OsddXR3RfcF7rQnWh8TcSWEoqY1m5zf0yxTM1tS7lfk
ZbF4CQKQvnUdR3vp2nzbVwYoj0VB4Y3y/UIP6c5JC5ok1kjQAPIcF96hkhyBWWf6
nNj0RKd5XaFRGOAe4FrDtDU0TCfIyOsl6lDnl2BIsDLE4ARsEbZdi4Bm8DIxUOCE
0KwGb/u2Sn1trs/bUwuLz/6IJic4GlOHBhvfiTKs3s5QdBcR0xmm4l4komFemQUE
vob1GZO/THkf8qiRzsdMTRNKzIR095rNG0Ie0fGKtolvmdPpr8YzYCIye2cf9Y83
+Xzxi+3oiUNxySIhZXjuxAZmcHqP2y1dHA5doAY1cl/sxa36V/9KxB7Q41OiJ7+B
Hov5r4ZnGA7m0fme4xyk4MDesJC3zIBNgykX2NeLpiMkxrMlmtIy0h4r+7DgcGYW
XnIkPTv6wvyB61iuyZyaAH072C8ZA/cudA5xsrHh6tbSdXExKW7PBqdE3md+QyH5
Dw5ZHfCkvAt8Rj/SCv3UvnHBV7T+GLKcktYsQEYEITQWwW8NoHDANRmVd2s5Z5t5
Hrrq4tXVo9WFbUydySaXs70xwFqbaPj075uczgDDKS9sr4kUTkGWSmHs6EOKTGUl
k92V1hEw3QPJF+WqUXmttUuMpjXygbFE2a6GYbGxxg7KTTqxDzcl9PhJ9iSnRcWh
SdptmPGUCphs4dCLEIRml/ekZVq1XzakgnqeslbGr59O0e3d9PuDLt4QYz5nDQG/
8dqtS3Xw4OOiL3OJPXcwo2hiWnkzo8tY2413TgkteSfHjSRacY2X18c8ZPphYiqB
l1rOVgj7TslpXmtTw3syys5WBPF8Nc4b+EXefg6vQnVlSd/f4N47vaa2AJ1KKD3N
h/Y6XJRXOkYxxJvI9VBFl0h7+T6IEG0AebsJu64ySu02WgDZ5UvNipHXcJs0URKm
v7hUASZ3FaaSpAdiiA9XWBADbnqgay5oFAexV0UagpQ5ZdlbPSwmVxCHOntPH/KJ
uOuGBa29dg9kqnDD8LNRBCBimOCjGxDPf19/GqLbW5EUbEyi2AzK8U/Y7wayPLA1
931oi1TDLsRk8mY75nvvheTvHsAR3f6Y+HgTHMOBe0Ywa5H1kcBE+QZCQwWGjcJ7
e2cLAj2LWQCIX/BkxE4SMSWrFyVys+eti+Wu+qvg3GSK3F+nFCLEzYVnH1CvRTA7
7ckgka8U2nqMTsL4mZHFH9Npw6ep9WQc0U/XzNxBzahZHDjSkK5WnTyK7C9aHcgz
xaPvE9uQV4viH6g7gT+iQJfGd99E7tvr5wp/GgmeS5e59eHWMHJ1ADzI1uqyMzna
uVLtexRpY5FqqyUpTItxvSVXSPKnXz7LtwLJGzBvw1tzTxU1Ny8XQOCCPufSANZB
IhW4a+68GRLgVj/Y/YsIMP+nMNqW0qiojB+K5VPtuPBDCajgYsiZGbCaEmLHBpVP
P+kwSwIy9fi4j1qxC5pBZPKd3H5iw7MBHOePl1J/4/AWHy2UjLMmdJS46g5C1Fr7
etwIw+GQ1tSsk0xQdlOLS+OugdaOnekFltJpG6RN8RpO1GKlqPHPVX29+orvM9QO
V+HJUnRnXDdpmRRNzb8uWvQY1/sz8rxLMEyUXecIOG1HCQI6thy/7XVlgq1rwqnl
aj8NQIadMN+yiD9yUgyQfN0lOdqOgqRPzpRg+DY6jWUcHJf35OonHfdNEItwnXNM
JmrYyexl+d0m1IRevjGb0Q++R4v0S0bxwPzWkvZalE+O4h9UkPfpoLcBUOfJ4kop
4XuNYMfm3gtCZBCHCzXghTdociF+c2e/VXO760b4JEmWGRiH2ffxXvC48ixaoxwX
083IA5HkDLzx6+pccQka0R0WxoBOnOD56nqfoqGBwdBCVjcgG+gluKOIV/0TPHg3
bEygszEPwFsi6bNXSmdghv0xi/gfNFMH+Lee+cA9H6dG/4//T+pnejFHPjCM1CqP
rHi039/Geh3PejEOLxXDfj4BpkpoNI3OUlW2tgxeglmv+uhg7qLFlb9ytMGKZx9z
MpXuwa/RvjZveqnjLOlsyda8wI5kwTdBWCz8/EPjcLlo2/MAULgTlGsmhrLoxBPN
x5uwW82aztgZ/qmXH+OzQW8V4CSnfS+J5u1bUH7B/RRkA40h3xRd3eqXOC992tKo
WaM+mn1uk1dmt0Fb5h2hlRpZt7Tasj6pTb6Zdi0uX4ltZ994fvKROxotiyL9o82N
92ulpViW4FKIfA8srBPpmmY40Xw6+jSaJiEjW39LGP41A+jx2FVolOMrjVd6fXbc
lgLgS6T69XWHbuOhyYVLdNjr3QaGWpBq5iWVCqpOvgRzedWFNO2U+0Zq3yCc52GP
2VPm3asNWLG+zlVfB2AVu6iPjDDeiqJJvfE7Yp3C4dQr5cAwamG2n56sJupleFXg
6oxwUNTtCHJwEZRsyWFbTbe7BudpyT43KSWDPNTSEnsOT35eab7G/dsvMIUrOKDb
4bjvUvG+NgGSCSZWqOd4AiHAkeG2CkDIgvynchYN6iPC6wBy0uwCeUgxD/beVuAf
qBZ7LAnYw16eqgu6Jf9BH51azvtfS/EakoHafLnGacNXjqZHQ+SuLdoqCBsLhlxW
vY1TYyC39B2+YGw+2H5NHoggdSItY4FFSh4AXTxlDp6T2q7Zp0MBStVHwoztz3Bc
47o4jAp3TDe6f8cadcSaVYdCo6Gh5VZZOKEs4qOJwb9cUJN8u3836ur6keDP/BSd
JxDPQ8/+i3rlgzP0lPgpYOB0uqowFa4Yb7Yv4CimEp2oRP7JUIWE8Q9WfAfJRmfv
wEwqndlLecENlkAAA2Xg61p9FB4B/0r9MMCC0+OrSHHwzwjTEu2ML1Ujdj36pANO
qpVrqV9gxILAeH/K/hRjf85NsjWL5t9B+MzSF2IaYqzv/NAU07KQjzeVBfPzGAFy
WtzZEMhIySGkgkqEFv7/aVdm4rTLltRcImX42e4QrKxI4okYJrCgKI9LyLBTPjUu
hPIBez0Gqoha8rdlT8WHfmPUxxtr6vJ0HI88yq4iQmlCWHmKg44ECw9VDTFeu7eo
ex4KSQ3X/7uK5Ede/YTmgwQPWyIbW7foi7cYKi5ezXvziR+fIqqRKSy9xwl1MhQ6
NGw4JNkYriBoY1Fdmg8o96Sn5114xkFTLixGG40ORtAyp4hIweEk0+amda/7jKaq
hzmrRXz9XEOCzmfR4kqC9LyEi7hNv7yxVnSHcg5YV6NvRhh4y/QTU+thgGiltqPo
jTa+tVyip1Mr06WZibvoTL+lFcDZUaf7QEfr4aKOqpWM21BCql9Vg2nvbzEUJHr1
i7WTaXmFbHnQf72pYsCmIP9agZ82GCm5g4ncVn8u6uibIJ3xlZdD0T4oRYvfmA4w
ntDkaliT1C7BcB2QAiCO45L2o2Mmx5tFoBLuqGASy028IbWWqX7oeyaeXYnmG+Mi
os+uLAPNvB+R8Bll42SPcI38LsO3HBcpPA7+gnlP6vN3DNgcWqbE+Aqjo48JVUFv
d2ZvHpSEO/VSNqVLYl6dxB1CdbBTOKjxBJIEN+xID1FyrmojJcuvgNc+7b5mwSN3
QzuBkvKhK5yR0tCGx8YRnOn8B574wNfTNToqlVjzB3/DiUN2pyQuq5HaOHwJuwgN
TqzskOkb0VNsI6ZguNqlwclFErK0xYrgMtPzjYjFLs0aueMQdT50EE2draElszwz
VlRi5nGI+jpmpDZXpB4FMcTKEe0It6yyFgFemAxe8teWkfQ8xhHe398UQSa4BYQO
KmMlYo5WQt4CBh61efTI0xiyZ0ol9PORHGhijE6fX1mZJimwcasYBsS/Cv4KrJol
ctZEZLu75/1QoCY53lA5j7xgZep+VMRVkOaxuf0gau32fVCQMNpFg4NWyJElCMVJ
ZdhMEE4L69O+IY1MsaEm6ufC48OUQrB9xcIFDwRtvwtPfq0RVTD23rJhGdA7uZbS
KWAzMDNnMtuDJQFxSZiPoUJwgvg98rEDeGP12hOrz/W0bBNWYXfaHehdAUhhWyv9
mEXnfGZSeslSxLOShdDlYvd4t1FkTpmOB2K4tN96dSg1j4f4LEzmrd2dzKw2cq2C
ftM9Nlt88zAxIGev1MO+LwQXYTSnkL/1rR40cjU0NZ98NamwZMDh8Ur+VjeyYs6J
+hfDrRmLgPiqB52QF/xZXboHh+XXt5t49piZYJI6wIX4Ttsgw0SLcQwKM/HItmD5
F7ewh5w3wv9bxdLGEzozxRLDCt4sJfZjCPsUpYFsDOD0FDVUUfqjFWFRF4LlATmk
OcPFm1scosDrqJH+z66XaGfTPXEm2O8VKJ8Z7kukUbLoSiNJsUr5c+gS3CnnXthU
/enMsE5kBUGl6MVNPooiIrOGMEYcGFiS+Ek7VxTOObK38kpX/8P2H9x6msw5Htg0
x1Dwk/yhWTPjXke10YOcO6M8yGrtqPjJcElKQXy5oaAgQJPHrjHD9lTwRXJOLRZv
b0uvnM2FN8MZD+OBJJHVyJpgjbpvU5yapdktpHTGk1fGMMqIiJPSkfTk3lwoGS7O
5KKYjuRRzeotWtO3iAM3Tbo+jt7HK6x2CTPxGt9hAmxoqQKjGsbNygmimbqDUiIC
UT6AGsruzWIkx4eblHw75BuSbjGG3LyKnJKhwGidzvg9lCiqq8DRxWxhcJyG3VCx
rBXAuuhZJFaGiD/1G64zp1BsJaSu2wjF3Jw+FiPmMWu4rNwS8boCC2Q8Yc2kGZ4y
sTVItuBgKP7azvqD//7n2deJZWe3qtMpATuER2J1aq/dyRlsNNGwZ7Rzk90AbTez
eVMUuYOZFY03Qgqvc5gWQspRcNf5Lw8dZ0mRDQSi2+H14ekhKZQhjBQt3LJKjvF1
HuxOJbFNKXphtSx24Q77hnBcDJPCRSiA9A9ib9ANcJZNlkRvH7yIUG/jXQptXMZK
Q8NP0OqSc5UOZYUyoWgC9PdnKwmgVOr4pC3JnfcfhDbWmHj/q4I0av8z4FeY5Ull
qT7RshmxTobJcV2+bOXpsqsozhPh8fe9cwlEpeLd6egH5gSQ0NZW3uICT54WHooD
FIuIttys4A3xWViYOKKgIBvKZsqvCqtSZrTdLp4jI+2qjfd4PDKcI/5sJ3ERgs0l
XLv3UA1S0MuGFkl2VWdOxIFmRFegX4tQbYLXnoRoXTQ7mTVOp7DdOy27ihwXbb7f
lFDXc/atEvl0Wcb8Ujlu5PSeZUSYZpfnelOFi5Ozt927OC7gfag6Z3100W94BkcX
uP7PZYJ3CyDqqtno2n6/2su7oqztbAb56uSuvkWoRv6a0uKnNA6EZVLw/q8VN5+f
gVeuQFCryvjwv9JeR1i+oVSg6J4YMag93A3K7ZCZLul0oGlyIeEFAuqnS1CYcdVm
dQ9y3mMj61vrMAw9kBfqMlx6yvxwhxqOlATJNIOcghrnsCtHNE42fT/cVHMdklAd
9Nxzg5g5yM+Vmiss841634X3lP1K/HAESmntTG4FedklJhj+4HuHZ5uNscWu/EBo
WZ9E/fQSStqA1KYLCs5iAUV6624k3FrxA+3MZbCfDU6zZRCoBQh/83Xf6naGpIM1
ncm6+2NU9L8Uh/4GOMFk6rDYOAzIfLD1ea1ISM57fjMRWTP3T9TPWVcIn46MZefe
uV9WszNJ/i2Kp+dUXNEO7j/k6MwM6NC+lXxQDbNrYqrTWs47KUloNCgxxI17vC9N
DbCBTm8Jz3AWVDkiGhKRbfamT22py7bx+5TfXOYLpd+kxvmR1nxGR5DgVR/IDScV
S+N+1MSrkfkNtSyAO5AHSrA7gowkUyUYIpYcW+hNYVdjx+YEq7OIPCdJN4LLMJUH
DCLGoEY9yrGmZk024X1ECBrcfKaGUBsCBJtRaNO+NDeYR/3AaMfYWh2qKvt8DoK1
Rc17T8Kmw4ZZ8D0bGXq8w3P5g1d2CDdh3mMwzC9rc+dNQQjhraLo6dH99lsrDeNB
KuI9g118C90vTfoBLTbU7mshwsmFBR6hZfifoL4FdiLLhfbOt8FAvUihcgAhsRR/
14ZBx1ApXePBIUq3oEA8YSyuqdf24zo6JZK348ZisNefiAEIgs3THcSJo3VMOSTt
qHnS2+HpY1UIHiCeL5mv3wkDcNk55QD5UPrhpYREF/HtkB6m8tmSgn8Hk449TNGk
8GbfrFpkg53aChNxqy16s/256lOVaF4ejAUoT2aP07+ccKTaRUFbxbH87RSctJYx
db7+y5kj+ujad9gx8bMgaBXBQL6NMsrAOIyp4x7Atv1PCV1CtEz0mHBsyqgPM8C7
tzSV4oDB+P2gRGRuEcFVg59pt9PzuV67+1SzscZrHZ7v21YTB5CNBG9h3U/L1cLm
CGLwCqaK/1Ub08xaPx1wVj+2zXyyxbgMDEiLtd441WV1SfP+Bhtbv/RMtdm+S+xT
mqzMiTIZqPfw7cPA9tsvTBCbtx2+ZlCI+VaECerpNNrn6HqH7SOfnCMVGN0I5mqQ
VRXIOi1Ko0SdI1CSZft7HaRF4ZJJpgRESxCxUgj2vLdWakpMSridPvVQVF084ZnC
ZmPJLhr8ZxsjIdAzEe4Efzq11OaVlK+6BdI80cOiavOE2zKNk6Yn9FzbnO89xUz9
KH2Utd8XrNzwQ2/G0K5pckkMQ2I3MltxsB3oaZ/XdObOrh6qSgEPXsAD+d0tvwnS
4mLNNLnHR7gaULBNzs1cEU9ZZLOdr833TbSoBf5oOzq+TVurtDsonMUGc0IfHscV
bfNLs2haGGhEteK81hRM/chwNNp/rkFtexEGdvkUiOp4WTJ6KgM8nQJACIb7CV29
Y0NiJ7yxqjiUoyiYbNIXCm7RjqaQ3lULy8B3y37KJfpzSJS4sowO0Omijb9EJ07Z
TQPrHCAacORgrOhCBpn3O1tqf2r4GTQftLbv5ORfA2LMR64R3btHYMRqEWERob7q
KiRovYgJjygWkEzffpCnZ6R2CgcV31t2L30VGVYwqg+1CbOIvWYZTPrCbdHsWpkp
lf3BmT5jsnld8olcLgmQ9Ews8zS7sQciABvt+jS5trbwOZAokAW0t1f4cgsoimCX
ZCRFs42kRCKlT3iPtDshoSkVpVga4+Ak5rGg3z+68ytloi06y7s6SOaB1ka2fgtf
rloQOI/KtqlYfHsHTrFpeojch0ulglQ8qUl+34PAWJtXm4D8aMVJXevLEF63BAPi
B9Ek9Yvzy2OfLAGTIsezX1aF58WKsxELzD3ZXSl+rEkT15AJPfmBl0B7wDWj/Pmn
0JqmxUq7lCe7N9112GDma7AXrNxXgOcEq05RtUcKBPOALWyBCTpqlbjyzOybcGuK
0SlgaCI/D7aCYtdvvoQZwKbbvGcZ5wuhM6UUgnXGPn6NFjRmPS3tsgPN2jfCbsTs
9Ch/GBQi/rwqz8rRMKW/p7Jl1gEMBnmgHnP/TOnVg5KL1/Zltf+jKhdtm8UVn4mV
1eJ9yyJs4RLmrKjru/Edi+tTIUdHaJQL+wFkxeVz3Q6J93JYjA43kZRIYc/K9U4F
P2P2X8agA68vfU+8NwZHUeAX8TbDqwH9xf1e6JxxA3o97BjWTaW4jFRIHQ25rh1P
5aBj/LgJLwBZmgxfr5eiO1jM8WQLe5V7Df9Z8C0FwHDx6jcCu5hIaEIgufwov7jh
/UlgTa5NWWMoeCrrzbC6nKPRqIb3Gtu3XQYzgipUMJpXvHqaW/cUZakVClYvqael
xNBSBvA5V8Hs8FjwqfqVOdsHuA5IrN0D0E94lhbQ6jywav5iCVOAAtrrEied5ATD
GGk4Uxq2b5yFTvNtKaygQqf+VyPZDSOeueW2buIMA1mTMKVnys925eV5V3iDX8kS
+UUsnK6x7oiSOxbw4y+ovey8VJo9+kQm8DpkIWBxp3nh5uaph5IdgvGFZdu9PhFg
hC+3LwxjFgtDTcUp8SSmqK/X0DSx9kQKI734sPrPoz0YBmNjwWKtaJ3uHArp/gNi
Cg84MzHCpz+oiGJ+IAcKrXlJ68qCV8/TTtkgWI9YzUFguH/xyzYKk7sEBJweTqjG
Gtq8FhygYXzqlrGuD2I4sq3hknxzDofrZ0ukljQZ2eUcO2dm3RkGgzK8bmij/Iqq
Qn2BlzST5GRljMsxEMGVxZ+4aMNfpNzaEu3kHtZ9yXGCoPgSMJH0y2qSm5kBrte3
2iSnBC2EkD8qAtXN5dDs6Z8lLdHDJPiNczx1GAVeVcPzlkWbV91SQipAYrU2W1vo
nAei1RMlqjEbG4VrVgdghAAZmIg+sIui09zIQcTberv62V5D3u6ZNlQQBfI/1Unb
WT34sB5KhAY+8kcYmMXUG/VEIbMQ/m6g75wH+qqmqFajYH+ZRodEL0LHzxZGZAUD
ooi89/SEBLcJT46irLlzS4TJfmdK2lLkZdJv82+BB/HKlrU01Gq57v+vmxGtXqGt
8EePL+UxzpMm4nGBClHstLCtb2V0vKW6ndwQHq24A972BHUpl2gSYoLrHutsjFZ/
UN5K2XkP0jeMmUr+v1+Fzxhs9zmGfvk930uTnXhX4btZYTgq8Sp8lRnVhHN+SK+h
Cq8qHqYVP7y+qq2AVYo91rlOHtqyOtuPGuzLLDuqWEhPCje+0qG9zg90ZZnN1fmC
BWDaXMDyr3S1B2bpuIJnK6G86r0QcOjyR1OvgbdDdUW8yEmHIC1Zp828cyYuxeyd
brEdpFUq8i5YWqWB+u19TIMA/PM0CbLrjvIuQRAj7yyW9BFUVmeBuczmZnDIcajX
+gplwN8fLq6Ypj+gz/FAHV3/mGwam0lV7YY3u3UTAJaz1p7xsA+2rgh2nQMWO2tl
w+9tf7pjNxlyd7pniEX0cofqOaQsZz4IP8EoAkwek2peeEQvY7jAQyCz72+xVK6t
xVdjZIW10Rc3G5Zi/q9GFfNBelqjR5gier/dl7K9pOwEsHHvKTSnz6HDkB3xeW/i
qlJFHPYGqTQepDiu2W9UwkM+wF4XCBEwHMEPKFbeLW95LrRdSxOCQ8viWb/Btibd
uDC2b8HNxB/zMiC2x9CfFqzBye53i0ZIl/GU9Mpgapx+Wks87T6XObOCqKBiz+p0
AsRWMzzb64xyEJpaPwQ0lX1P/FLbwECJmkbg0vgCkJVTBY+KMgS169gXFMPgIMtF
wZO0lgMoVhCKbF9HcOrHulVZsN+qPXL5ie6yEfEt15u0RlUudkQQaRdGaiqcy17c
MAM1HMBbEiqnN7KDWXsUiKTQfnipMMfr5nIHaN5kAIWnmeLaKNfcMJzNslrvdfRF
sEQfezbGnv+l2RjrCeg2Kp+QxVa5EzClaOOvDXNDOaMbdIIj7gomFCYTIUSk5Nd0
Evq03CH99jTNILg4vxGeNAyh7pT8mReM0gBSPhRYm3IZKLUoNcMxqEhmyKDwOxdu
3Qqq2w2vUlv3zG14k/IVfidhTfiMDcYoCeXzDTIdRp6qQEDN308QfRI3wCS8uQ1I
Rkr/BONFYjszW8zcWO8LFQ2/+lo2CnPxRTvWmLWDj2z3/Wd1ciKoWm0Un4I3rkxY
3zvwf4/AadiMLhxxcwOO5OwBGATUwKHajAoLMLrXns1l+dhUM6Tp6RC4uqByaE2X
CrkbjeD3OFCm3yv+yvVOQHNM4wEzXb5FMQLRGxR+4ZD8Lc1qT8fmMq/XJ0+cd1jl
sJLyU/aT1BSGtxGYJPBo7jRoUwWweCa0ti19VlVLPvZXbaJ2+F7/xIDEQ8w99U4Q
/I6Ze8HQv1w0Hel4Z1qtH7SQi2O483eTpUZftE2uMP4g5nqaZdIh2lkDwRsLkp8i
Myef+VLHcPGfSZWXGncmEwtBGPxmT8a/jhfpfr3gvs15Z7kcR2LNySdhY2N1ZFI9
3hh+S4ZkdGROa2YmC6bErBCHXlyeIDxGP9+jPr8cpfaBp41wAEDFi5qKtGBVpIhJ
eDxnkkmp3hKPU3eO4O+Hx754WIKOeJ0dZN1BVmGb3GS0HOJl+O0NcSqiiAC9DqpP
GWO7F5RGNorAuibq+ynHWyIxas92dUaW2GqPV8tg1a4zqPe7lpFEnLTCcd1U4C+0
4K0KlPkjOqEd2PUJygfFLTO5sPcml0XEAhjd+AqTFZ0hPlu3aSDHJjvuLj1a9XFw
VV8X4/ybVe/KmdqyPsUM8pBV/G4oyNTBtkhiNCaJu69CkyKLDSJg7Zt0gvHTdVRu
BIB4yIFhmPW36hYMRToPTh0HirMlkB20+VzDbbcTe6T5RXPmbP7SS92lymrG++g3
kp9/Zemu7KzxsLTVKL1zOf/ThCMFIQAVq7FR51NnrFMHz2x5+D5fnvuXI0rEy6TK
XF0neoRirf8UNy2sUyN+IG3dAHusdOMsI1y8ebLF75Au6Oe3GZtDOtg5xkIK1PkN
JR5QFeCckmi2HanoIo1VDrmCYqCXN1jwYX5F4dte5cFH9ea5Ll1H/A8oN8r11AKr
glmSqInRL6bWR0xA/RZjgJdron36JKnsao720aoXFVa8hge8Z0CIK16ORB5YVr3G
WS2OcDUnxO5wk5lAnKuY9lsB0SzEAcqgyNSGFBaytaC6oGM10MSQ9hglpaNFpbNQ
qJ9Ex70bAu4RoCPe8jJpFncUiBg6mlSenvMNdhjIvJNUTC7YQ/MBgxaX12Wu8mpc
FL16faaQYM2VfwcZln9C7QWfn5UhDB/NBSlAqG75i5Q1DJWfbDJoNQRy1UkXO800
dfQxt7tz1blocQ1vKJydcKRPDvy5gNKG704e0Z4T1u3BDIKYatUuCdUAkwHGxRhu
ha29pgFbeiNQ0okNdyi6DENahiJ6OpON/txmyu9k/2To47C7q9Ht/B0ekuPzn+fm
Du6o/ckN6vQVMx36tQf2t39rYrFzdS+UzmFOc+mG7XDqg8QNGSUTmfRl5kyTxCju
i3rvzSQkvT3Rmk5Y4XKYzZKC4vkzLLL+lYw/rKmgj9IDTu8OSVwdKxaPdZZOipVF
FcBpXq0+B0aXckRlqo0rMb2WxL3L+FwX6vqKkty7G7mFdmZ4kO2izSTObvujWY6I
sHbjqKgo6TCkMdC/P/gGsCccceYsUzd7MWOH8McZB+ot3nTNsqG8jdnwWAgLhDwT
5phDCQ9JDoClPehG22JW/h9Y/caa0DC0L9cBgmKCHqZ+maPc5mfYl2rdy11Ts9AP
ppMUsQpzsPDqt7/6aKAYU/4UES6iDjPTTdk8KQQsM7GYrriQaAKnU+6yBAN4AZ+F
yUMPzjiDxvwoJV/yZC8/8FX7byMVvrYGN8CmRQFxOipDjGxu7j12vyPHJe/5dW7z
v0LtGHumw97hblXzn5oT3dKfki/2BSSMu1jYPEKuNKbidiQaEZhehWr0aNL0fkYh
XDU9olccgQHeJqAkadXt4KoXhthNjLY6GUUCuTU4uQPJyCjlkTVfjmlC27jPzGz6
OR9VfaG0duAv2gTbvlKr28rScPECz47d87Y9VXoLTwb8a5/UTgKbcoqAb/Tw/4kF
hczPusbYYAKxbWJXYuif1IUuFfZKo0haY2hxohrd/0joDh/jkIisl0ntOr2dwuuS
Hb0buUNUElZb0PqQsH3KcbSZoUid7ZCWLaRhJGVFtuIL2Wxxu3yOUCtnlmrA5An1
Ou9xtZkAEYOUETeCniaeDl4R5M0Y6NIZfxBbgtq0uQi6WqKkY08JsJ3gxcdy4WmX
Md3/f0bTmY9JJn/AuH16s33Qb0boR/RN0tXgoqx2hMsvQxkcYNsmPP0Znm21zvF9
z/JBJFkzQqCRbmnPm+t2zAUf6OKVbGgLs8waS8udh9jAcdTS6evbHm6yJVM4ILRa
0eBWsQx+0lJ7Fp3s2FoTDlZ8WJfX/P8GkEhqtGBXFiKB1jFWmsgbncEg7Yto5XqZ
/8GreYnQFOYLHXTW7fjDsc13h+Dh1rnhAdJqIUYmGG77C8E5Sb9r7Ikmfo2g1XEr
geTeJ+f8HhmnJxOlxiko2x1IdlqLrpC8rvCNLqEc+EdcvwvR6C3zlDjz6lweDMTG
tADQ6CxODZxHWnFHxxswaXd3PvHF1oMEvWru2akit34REDuObg3VptSyUkvRh6Zh
qvYX/hD3TtatK9JPfgVPJQF7wBgHCqOUV4HwfKPo6gAq8ruPAvBUetCSoE7+8xwZ
eXgCrofOI61dbU0WNfyzuzwgB5WBpVOb4urQb7LF+Ou8HsSlKVzLc6wYODiwGVb2
rmagclSSRDCYHbq/jx0zOICGPjy2Z0g05aPFSDDSFP/TTJ5Fk1C7CXOM8NlE657r
1lltbctusXPdhDoYD+kE55SnsDWYuZ/nWYTqm0eM9tp0bc9klUKAatHC74PnB7Gv
TIBJUEQWp6A1RwYuAcVEYI6sQ1tiJOXkjho+4dsON+Rm77ucH4cUWmtzQ3cOuxO/
HaMRSVfOwJWkOtCsMDYbEiGqKSZ8WJhyIAe8rCWs6AHxP9Y8K0efCWg4WBfjVJU+
SSKzB4mW+y+taNmL3F3DTfCRCP/KPReqoj4lH8yKa2BIRAsgkRyF0p2zH18rySL5
z5D5tFVBz3QMZ9VhglPgGPregrixFxPBG+ZKic6ED0pBYyfYWZvD8thziFGiwNNs
lQNrZj9w4D5DIuXxX2mBrJWlnMUOv4e2LRacbWBRQdGE1cz8Vf69pYG/m1975vlJ
7fV/Vn34aatjJbonpKldmFcXcrDvOLrfMVJzjFlif5JNzod6QhbrHAbVvecwio2Q
fb0JAzWmwJmKDYKmxAFrJnxxBLlS83s/OBX4zRMt08oo+RDmpf0Hbzhi9XDyrsB1
UooT4JgYfksxabw2c+hs0x1P2EcC9lOx5YfFRBwRx7ykPpvbL9T9JGo6/H1z5thJ
nLFRfhL0Ab+1TL3uerho6f0tk808LwDzn86MhfiqjM0YqbbKsqnHf+O1fU82KNbu
OUbY3XePR8mUzdWwL0JUGG/LZwB3ad1ts1peY08YGD6eUSHa9LmzFXfiAgJqV4hC
1ZD+0s+vTpfA+TsnyIB8Hdl6NTtKuDEhIiSUgi5dVjgsg1jjqussBmUkfZMjVfGH
nBq/4lMYWGU2wKb7k+AruhfSrukbNeyTKNIeVOJmQtz9HsbEwJO8IZbTmlLypoJb
yYeXsl+V9H+pm3NgIATWRxtHZwH5B0ZU7QTopUCgliwJbBIrZ5zqSPDbE/ZGN/mg
1Bxvk3ch2eAo0Vq7tPySbqMnxqnfZiK+qdVmAahNQv9Zo9DffBnEpwuJajtU7diY
Sgpb2H1RntMJeeQh3elL1V9MOGwWVtVLLANfo4+hnKkxWV4d95UU6y7fHw1+vQ8T
gfMUwe3upvkemqxfAhrhaFsqvqJitVWHfPMUs3fDGJTyVOBXl5CVo4LdPoZPIDIK
EOszrGkRNRF1sEXWGb5bFEBppPl9a7HtkA1uyqSGJ7+HY4XodhSO0Q+i3zpOzMvo
CKrhBxDjW5oxQznKhUCwKtVbeigjGI0pJC8+SJU28OrDn1QjRLGVLJPjeW7Ejr4i
a/mw0TrtRZC6pu7IN/fCF9c9tI9rILgdrCqYhcjGsGA14ry6SUAD+R+pQxAAsLht
Zk+Fj+lnoiP3Hh/harXETbew0SjQErkQYOPtv0cZumg3g5/uOeQ4sCj4rBH6sxgV
h470ulRZ9Uf13nu1hAbNfkCzMIdvM+zIw7j9z33mN2Wji4myLNlpZBLQXVwFTmuh
TGBXL1VFDKHbFgM5CS0J+MQDXHKuwUA5tNaZE2wZoQkGPIb2DGVtpH7Gus1UhQbF
42rXIkOyzIq5n/9QFmHihAdLN41pbp6V/xR+MfyGwI+XM+RIoC+I73A8vQ7Hy1Rd
Ztr9BKvWIcbZZnx9VmRW7Pd4euX7YoEVEYHl94b09kZXoYWWqvmgEFa9ecOtKS5Y
8sVbFaRC41XCQdGSPJwsA/fLYPMtYaePXKEczJI0wxgRW/C1P3G2g1yr03y+pahm
9/RWbbzKMcqRYorqGdxLatbqXABlb6jyxQxkt6Zq1O6U6xqFMsKNN2FU+wcYakeC
rM63Ckik7/tSQ1Rc1KkW0vxN0nrbF05lk5rPzWW/JEBTPmAV5jd7XdvdyxgEhVeS
6kcAibulzOiBeYdOe9qG+ACb8wlE7+gpucWP0QUwHylpwQ4ON9APq5pi3Qb69S4x
6R+0NxqKLaouWyGzxtNYHwiL7klWmSYXL5LDJPRX/vPhUQ/eloumMv92jpeHLQVK
7lAubbqvvQ5O2meTnoaf+Nd4uX3hMMxYKcK5KdsnS2V9cDAgtFMziGv512lCPyT6
4SCjkeoU9qINf4buaFseRp3nEAGgBPKrhokeliMutax8NRW9mMiR4x9Zm5B8iEAM
qiKiXXwdriCUUt8RzQKB6Ca7l9GisvmxyKdvIu6jgd5Z94+PFjIq7w+dz12Lwzk7
Rvr9iPxbyKr5qpoJApnJOo0NPlkW94gYlr/K8UtQ/6JGRZ8gDCVA+FJHnFSdupkN
HCe/7hkkAi6FnmBVJOc4UYliuisrRKFegn7TBG8GU68WbHsFFn3aPjBM+4owl23n
ZxI3JI7XrQ8ItjVz7Ea+A97RCUN+F3t9cm/nvAjyMGGHqkiz9oNjQ+knu22ENit4
LBECnTf/8DXIFD9VOZxJItbKrQGd6wzN3PG0QfmXq0wQlDhSrEltFWhaykNg2ioK
65yHSk6HgrgVdIn9M3F6/VKzyUJoV5XUed5VIbHzmkhleR9kYKQWRvkCMbQ3QfgI
dSsrfK9tbCz+Pujya3OqSpznUF8cXJabQd4W4oDaQ//ahthalboQoV7Vb4RE0/Sx
iC4DUErYxhgfAGk8Nqef9c8KHKB/4KYehW/llOMfXSbArpuJj295BpsDMcjfBxdo
i5fbL5+Ibi26G5UZBTw1C9LxRE/JNqYuc9UgRuZWijmC8i2KzJri3nfohQpvSnot
HACATM43g4W8KOxGcPEcfFb9i8N1W8XvHRuDAbJWupWjjwQ4tirZtV68PFY71cuQ
Kqn7MjXv2BvWzBC+D3tX7CIKP1UnNjkYhV3/3kITyvaDnu9iBTn4CVrSgkVbn9US
HxstTmhKHT6s8URxlBiSa2alXRJtTuVpNw4aT45YwlzGb3eulgpbmJfMH8LZAXXI
u6VNWrgNLoSUzxjNS8LL8nu8icWRiOk4Vw3xgIx33Q7bq01iM9PXWbi6ntDXozZk
RnMUaYPfwNecMNESRsXHh/bzUwSV3MTjoxpN9vKB6283c0jOvTz6Zvg0R0Hp8c1I
FWhgoG+bKShPo1YGvpVMPoRs1M9C4tMizih1KblP4CERckz/Ja8oBdUATqOvtSyW
KN3jaWTVselYLFtUDSDOmYPbsgWNjTNKXo5KpNvOAdzhfPoteofoyQxrBQ8UByBL
uvsU+5GeALWtp4xxvBe/yJfQMuMAe93fsBClsPeI+RQly762g8I5sBE56/d9Zu/X
Cl7XDgLBAnS75EGEvmKemFP/31talqVcxRC8JEH/UxvwOyQLJkS3NhKH2eZnlgGQ
fCXJ/ze96ExkfIFFyW5Rl+gOGZy0IBJKbAHaYo2wsbYL3FUlSWEvtQSKZqFY7lpL
T6vSh5A5nHxuHIZ6ZKqeqyC4VCjKIrBYEpPcjUFZlwZwVZU3lHUd75RZ4DFiqKpQ
o1s1AIb8lhzb/MGJyaKZxdk27VQznDW3QnfWKiYeK7zT0gLvNy6CFWe8WqoYTdbN
z1paWJxDxD+DwxvsnFCsbZS4B4T20aAr3T49bDJwmyVZSGoE4alt6Yr0mEWGU8vo
4JmB4EnaPS78O/29cq+zmuldxKk5y6dFXR+YN0dHZ2TgP5F+yDGqHL4ftzEWAAsc
TzrGKUZd1O7dbS4yWZOgogeXMBsLLGreTrDFNC0pGpzxJxP+AoSwXDHkIWfcPVi1
uFmbJBNj0dJKOJs7IafWrOHy8CTDco4nRERCimMIZzPnfdV+shxZr+KGLu8yfIdy
mQLtGxeJRh/l+dYhntCY/M1fwr4jTXAI182Y/L+Xv23s6PPsx0IlRXoAoD/PwXeG
C6+jQAG7Nxc1Xhz7oPeI5+9V1rYLIxam2lPTMc/AujF1sovtlmmBbhw9cQ6cDZOS
BnEGMSfWdCHgRe90Z+bfdOZ8LTD7e1MvSuPCiIGgYA4dptq7yzcbDZQUmSIXSA0V
ebw1xSlhomBU+1dLxF3s6MFiBtXPUCCiZGCMhZ7ufgTlj2OgdJlsmnF5+Aj6asQy
h2cPRhhGAZ31EoUmGuN/K45PR/31OE0mXqgSBTHdfB6PF8dycKgNTG0r5iz0C5YL
if3G/MZhdJBnHnlDV3klFudKWVBe8jWednUdTbl+S+HZ2DU7lzktg9tpz9gx5HOE
+ZM0VsgydKua+1tlrC7r+AIJQoEQ1Bvlkn6mTLDoRGYSBmxiuLOYePq/kKU74ODi
MpZY/jQz9XGzUkEn+mkbq9lsp6cOhixhVGoBDbhUwwahf+AMJ7p12kQbGQco8TdH
9vsGzb9ZFKtgmrvS5OoPAu89zOb+5qOWrqlyxvNLTT/g3J/U9cM7+FsMjrCtdBQj
y7kpo3rG4pIfHL9Ggfdh/xVqLsaMZ+uN+moPow1SYGahRx++ghb9lLnOjpvSbzr8
uggiQi7jIfIA9snWbChJeg1Y9ZEUOQVeNWCXEFjnYTrKT7UqwB+Xrb1uwrbn0SqQ
URjbSq5Fw4TU2FiDSpcX1njaNDxGY8qU5dGr1EaPBt/Np4d7kVODaHSBHWNd0rY6
jLon2Jv1anWc9VylhU0X1iluugA13mHGn0DU69VGtgrC3KLkbR15cY5T5J3/z598
fMQxg+SoPW2WgT1wUlfQkp6CJG1ghhN6mC3rEWI52Z8rzwNVf4HX3xdnlTLce4UJ
SRm/IS7Wm7Lx4c52vX+J3DqquZnFpehLhlOexh+h5fwhExIuKSyZg7CwtR/GjJ4S
zqcOsKWZc2BLeBs1bTB6kZtBFQlGjLbNxsp93B0lVNUbhVx85jLmrzlnXcksBh/7
rKO4xlCSFXobZTUYCveq/F4d7RRjfzJR5Mv1iymY8IdfblCCZWbJsbxFrf/NO0fP
fPMXWbpCyPnAKp9vu1cF+6eCuTpjzR85ZRTb5RbD6YF1eCABlCkEGcHov5EHNWXE
kwONP/NjBMkPZD4xSdlTlxhc6t/1qzrsdmuw74o+xnokAbTxuoQqSdLhV2Y5LoMq
1VdOftyXDzfOX6IOURa8BV+oAtlmgugGT/6gIBhjowBJptzfpG4CpetUesmVYCyR
2ZXgDvwgtlpSKty+OUM0XNHAKadkBAGUOJC6TRxyE+AiRvvIG1OnWNfl0fgNnd0O
F5351xHaMfI25brLx/twj7g7IofHbaCrTocwJczdwx60WqccnIkTI0sFz8mITCrd
u+4WBE5hBMjIgFrqNNxZQALqeYC9A3/nCIT4PGMgoYWVqWKRcqsaUVQmE0FPLpv7
hWXrKdPfE3a1rPDjpp6GTw+Z8vAoh6hnmCOylhLBOmE69Jn9mavP22icHqnA31BG
OmGs4rCriF+37KRBTXQCgnbZTTRCcHj7J9MhxeJHcZEFVpsZEGEa/KKfz9zx1Srb
qqt3cSVyOStb0em5cDeJxRBrpdaA0NMZ1pHyeGV+G8MyAJXNxsBMxFeEqCPaxSi9
zKR5ka07gOoLasDQY2mpaLbmJoiMpmii/OBq8LVKZtYkxltfiM0wO7odnddEQh8C
I3/ITn3z+7v17lORml0a7jIyqRSicfXNBg/qjDIqhUWOJBQIZmrmrqlC5EgAlGow
qiYu+gXMXSzn1itUhVtxB7ESI/pVuhSGa6qKKhNb2pjRCY4Vp9sdPScKDV3epdf4
p6x9EE3ErSng9pHP7ftLEJ8JJOgjvP2xywbrZyxGrqf6hKiTBRoc9IIbh3FJOs3j
UHmnVkMfMhX6TXJt3IjGYn+sbtWqalFB1MD9l+NUWX4c5UJeuKjozRYwX592TqMy
mtUmaKxrHqn+GHeGN3bUGgD6FR3fwIMed2XOe9QtrjDPWkZo/Jm7NFandQxTYvRX
EsyhgavA4nXxxcgyezyo/EgV5rh70VPzkbiQ4FIbYTdMil+sKi3H4v2IAS7OHFxM
pI8fNunPwO1Bp2SzVeBIQWhti0LkgGncmveoP1yis9+iO1GngyYimyOBoa8vRXhU
eJaBVSpZvddDVOh2NmaCbouPzq1lsg+bXaIagp0uOhh/gxNxHQP9HqW3ov9N1/sP
q7TDxIUWBVMaRImBBzfnTH+6g9iekrmcftaC6IxZyyb4coM4U2LO9CXgQgXJnr4v
6CuCA6Yqo0esjNH4YlWL9E70U/OAPAE4fld0LrWEH3xaAvlJ3OCohRyvcdxEb3/w
Llg0A6uJtDhQ6EfITMNnrhVoOM2Q/8wiWxcAxdhy9/al6e64QqXRZJlpD0NoAdH2
KvD5LHI0fuNZN3WAuychl+VwNNQ3JPGONoVkXXemnoSLXkkdgjKAno4T+321H/4v
EdSDOkLFZ01X8h8nxv1LCkAmvGviCh7KZKjieZkNeUIli0lh56lycQqPy7TXaWQZ
TpJ9nFdXV10zA6tSBBX6bW6WbkdKeodEkXbCReB36pTJ1ovrJccHqZj+Q/h7t+NJ
Fx4kArkn61t8rjvTXoOR/KeqH+m/Mx6UY6xt99ljzNzxWBalCNJ+8CfwjrVXVuwB
thHwHpQn27E+08bQB0yVzYhqAz8DmAEGVo2Aa1VVOdiuYtREZriGYE2HLfF0X+Qv
ZeUrfqWZ0FnMkaiyImZPSSb6V6pmSQYDRPceXDodwrcC+T1sLZ96z2niUKSi3lUW
x3hXLMFMKoV5gZNn8Kx4YHpKVBMGILuj7lZEKfTtG7tek233hP8rnZkEcx25oBtR
PIJSl/SbvRhbDsH4aSG43XM/m99ic5cfXu56hRKu6wla3lXN/ygsoDLOg86sqfxY
MnEbGKZRhK1cLVpHCjP2O1NPwh2aCegj2tWnflDBsWbs4ar/pRKzdSQyVqFmbCRl
BfUelNzghI206v4Ykw2Y6iSOrusfQTCSHF8KsUa+Irxq58OT+FrtmjsXeWlY40lu
BblWnH4J6CAeQSrrHsxyJTQ75YGb41cIuBytGzTbAHhAk9XjVyyB1GEzEtM0yale
rgIreTGv/knQRMagsiTGVwe5XF7oHWK3jL/1fW7WmoMPmCPoy0+TmL2AkUvh/J2/
Avhk0TbYE/iW21VSwDOPlV60HhTUcBPLO2kfCi2IcdHhV+e1hV09DL43HmcWRsPP
JY3/EAih+pIVGvnGpkWVzqN/+J2DPWMLnXSK80K3dvHpaovfLRsSi9hGzwwvx1Q0
WCSJ4FXJYCEPDUOp2iTHZT6xdo5v5OY1n7DtqER+dA7ywbQAHzSLWgZeWhzYHrpT
bALteidHIIwMBXclm50WKpWqgEbOjxLuxea2hqKYE6Ed4zo9+bLr3bj7ZZDGYmUd
YfqIh5QdKsI3YtsSvFtcM1akIQTCM87rFCBnDsmwQ6rM6HuhpxmiYWpOQvUC1xqp
DwEaAvuW9rrcno8AtF7j8elI+/Y5I7uIH2ih2T7yT+MPnsqLWHLYSgZZnoTd2BNf
2CbrSojckuf1DtyEFFbpad5e1ucn3m0DsKhIBNyXnXF6jJyjY6UV5pYPo/jyBuAU
LqMuZaS+Prvd3pg7O5qLzGQ3igM/QNptgoSfrGeg9jU6qU3hUa2QjFN+PA/sgsaW
pVqa+yL9m7XApZ3wTzTW4mk0FlYvpUXXGfIOkLQNOWmKMYaCBIS9EHg21KFABsWf
8bMY7k9sERTlqoHw3ygzzCLkN8kTzdZfR0IOhOgp5MEtwsYkzsqRMLKUF6HUmuID
KtYKQTCF90lVCUdtYkRgLSRzo1BkZzIXN8lFBg6WvIV+Yf6nNkpAGykSOXi9xhlX
1p/RzyR9PCe7w+LsYgRNJ+Iwe25ACIN/HDG76Fk//QDCtE8knBi7qheJhmweD7R/
rDjyHmYqk1pj+u54K3A6xCblXo2+euZ+uXcoaYMq3nkLkzO2VjlIlt2d2CTz62c1
/t2kby6KEMuP+MKqDI8i1AzB76uWeReLDd476DaJ5NizRWOQHURNhTqpNGR6KxMw
rIXEcLSM7Y5ede5KgeTsYGRwa89DeKdqS/JsAnn4tLohIn5ZD5f7zGLcb9rWpnjz
oKZoQg/sivIZ3G0C4fAvD5ldZ5B9EP07Gd7PhIYr7BH9HPmPfNt+3rjtN2fonB7W
Wd5GV2OBC4IHMFyywL5qYBAf7aWloVXZVeRjA7iKwlT45GIjFdr+eJk0KHHT4td4
brssysnECQCRbBpTmnE/lzgI6Nz9PEx65eTT0GXElpAAcd4xn8TlOy0ZWQ1J5XqB
i4yI2EPT6CEaZaCFeJxUSYYncwC+a8MtsX/NlZ/FMaLNIyVrnwJYtJdtARV9QRk4
aO3gCiiiuIrRUH42jkxekBWT6m5KYgmJ5NxdNMo704S6QtybC93BexbKDx+XeszX
TRdjZ23VSQxR7ltZ/3J2juI17F3jhvkSyJxeD5o1V2tUCoi2E3kBe3EuMsbHMjdt
iF1mOSNiYbT52dSdKFyOkQT3vOSzkjbXzS8SKuHeHM/UdjuMNPuuEnEVgKmCtPhJ
XraVGgV3KP67zHmY5cGqrpTSjVZPVuJnhNgSYsLYTLFzHUtZ56Guf/wLzpMOc3ad
Mr8b8acHsq6rD0yxo6pW0v/4pY4bR2/Aesha23O9eZHpihNlnvbaXKzMjaitF9PG
zUtEQUVXy4/8VA6Oxu3zfxUc7JssAiUmHBJRKP8ql/c+SKu8AW2cugsJXEIpdy76
++TM+sLNxY/V9arTsqpeP6gLlHCD14cLAOBYaggjC7iByH793/1QdCMvb2iutaxI
0JrnByGvP3MW6lyDRtES9acjVfvKJRYEVOW9WwgQNRdg/ve7ojZKqPu4oaBhnrlr
ZK9wyXrJqRVqW8G7DnAZkaDhevtF0rX/n1D2wO4fSC65mJYhN2/DOSxbVqSlcAJb
5ZzsKHjbyabfmFVLjZ0B6UXMt5iUEPkAB8oC5VxPDCO+VWB+gwThS7HZ+ETzJJzg
A/7omFuvxVx0p6oSR24u/hNOCNh84+3mI8cE0EWQMRToq43natjJlcku1Su7tOsb
1+slbd1uI4BW6o6bZKMthskmS4Qi3OJXl8C6MhC1K055EKfWKk/7FWkvURoezZ0l
4Pz4vNYstO5vfKIgz2LaZQ5CCUyCy2Nv9X53mV8ozRj9xm5VIKihxY8JDN+DcZrK
hq6xcGfHsPzfPyWqKqsy9m+RTC0X8vqVrWeOYyHIsKxVMbc0qtYYOJlin2yZ0fIB
jnAU1C1PczCHoy4ITDiy2jPVO0RCIh/uk8vBwcVKbKNYf+dxmk0jOutuKr72e96o
BP43T1fAKVeiZ/eYdHlCqt8g3y6YDaxmtCTcDHUJc0G2fDX+LN5K1WKhjybxor25
BdNwNoc7jLzoHoPN9daNmND3BVR6cIwdY3MGxPCIXefk+7/+nX95hQ4wjtepl25g
eEBhOJVujJY02mSV2PnaIBHEfYGn0GH1TsAO4Z4yB89V5FB2flmYrDg+j61NnB4D
MivkITrCcJm7thA8cO1BDHmPuTB7Uh1dnB+R1X6iJFWn+ATwYIYWRdjlfTKBRMWp
XWEYMXpno4axOanu1N+iI+X/jG06xV0CntTAAJxhUW7Ca9nZj/lkSUu+NGLe7ClK
F6UTo6y6LowXchbf77nkNvN2rA4Quyf/gHBRd8traMaen3awFdRuxAnUC04Lt48k
oLOCmb6CDIddng8d3fF9nfX6P5yUIB2QeIaBQxlMI16MI81LMNJgfSvZ9v2eGbwG
B/cauDyTwJ1RT2qs9JoMG9xyztoBX8ie7y30tcKSYtX9NiyPqWVS+1mPY2gBdnjq
5GZqiIA/YIkw0WOIHz2oFmtxCCqxTYPc8ybHEGRGNEeZ0Gy6ws0qSy7SCuH6KWK+
IWR4jp3cGxuxWMGiiwyVySFcC+yufmJhRr59aynYNxPJYT9rkzfzStN3apCkNFGQ
+vEm+0LJT4OTUbH2ENx1Grskhd0hvxnrPwKpNK1jbTrtl3miLXuQgAK1D2tl+146
aEu2sGY7z0/LUVDzrRqa8K14v7KxiYUzwtF+PK39/BE66xF8Esp8Tl3dGqXdB3Rf
z73pziCZPSf8cLoOWhuVcUph1ZsfFKImRwwAbmwJ3y0XdnR2kJhhg4CN/nciix/P
rFExiNnclwhisJJC02aI9rvbpU4VSolrfwr7rkQWe893HfmjuFKOBd0UV3V9Wgsr
Sv1qOHAKSgSYvF2Mzhgdyz3n2QehxnvmiNF8r5OqR7LNPjZb1s1qN4JikOV2e+kf
dHaup7WgN323yfs/LrPtvSny++aiC9iJMdgJyDysd0F06OXX9nm9GXtfKtmpMdI6
EKTJcVOA4MKUbqZQjlpRK+TJcX6Yu9MKWeDYAsqkvdvWcFv8gWJWqd18zp8y+XVy
iFC/JRXF1gS7g20bmjfRXHg/ipD41joArqRkYkPUZliZP8v2AFSc+2GCdpVTmlrD
+jMLvFD0JLjHl2I9fpb8d0SMDfsBD/tM1M/OZUKVKcusrBhw70lfRSaUPurQYxMJ
4ZmBN08M+KW3aRHk5nyCuoZksIjubRXhtdpw9WDmz2yvvqpGO4nx/hP7WQtrqTK9
FpSmTSzg06UAcYgh1GNNSeIaciUGEuXCmW3dWEEocV9REIISGm6V+8fkUmiN7EmH
nZQs63GQFwkwauYVS/10T5d/1thEUu8Ei+QttP8T8FZJ4qcTggjnRGVX9ilwn1KR
bg/zBSAMnIP/QpVINBIQ8/ld5kEpEXMynTWKA2gJBumH/5xUaFQaDnplgWteqUHq
7zYRFkN478eAHJD/ittNpmkqnc3awdCbGHAcEJuOJ1WgxVznljRk84BGzv/2yD83
XArsWeB4LDX+G0NsM9rGYxLGxBx6eL44nIA1cG1JqewiR5Cc0gzqFh1xbEsSGb/s
ThBB2+zd0MURcEZamOH2kKWyGfGNsOko4atgTcPXk2/3LnnMdPjfdLsSP1opBl8E
2kNhTUz5psh8KzjWwrMXs+ulaq48L0S+cADa/oKfVE3lUbiuzkRUBkx+Wk9JxvLh
ylfAUp6ZVQp6MZmMNhBUFxgMlWCwNO0ND8I9iyh4/YqTrrx344DiNpWiKvfFJY+i
KFjbFomTthnzgxQeRLn7XdVeh1Pery3wJut/A+VpdAlzJI2bTo7O9tTB2iqQxHFQ
93NVHVTdj4FXJ0TA+SR8PaCqfT4/jKPTiZSQIvBQpJY6dRtugYBAhZ3GUlPkVbVW
B2NyRJFtoRbZo0ESgHSV1/u0GRVEQb8FyIKbxrun1zkK4RTONDWo2l8qsv7uvCgM
88IeSvD3tjVmK3oVR++A2PKBcJEOWYKqgwmWm3lgRHbfrNHDR0ahJRUhxBzInfYU
v7ZAIMXD4uyCRc3b/3orxiLtsbEne4WxXW9uhftIDmNPPSrWfLVrsxIH0F4LgPAL
GzxTwjQi/yAdjsrKEu58ZqZ0/oOF52PICgPbkHOzYZ24qAsmHdY4uNXiV7VcxeHG
hWRN9pAZO62Ba7695QEj7f3LeDAePh8SGDbm5xYA3dLDG2OOuX3ozrL0Bu773dhj
hRrx60GTR/WwjrERTktFeLfH3Zqp4m+OpkwBf2PIENbjVUdR4Z3gBDXWegblnhnS
6/GJ6mJEP/MWG/wxhyM7QE1F0u/mhI2h3glMjIRZGK913yE5NAplvrYqB99keFkG
7mtukXw26k61BAHq/f8iKPR203J8ozClJjk1MQTYIXbfU3GKjypUNVCYjgQYJEos
VJgnSkI0wG3OaVphu/R4y81zEHULEQhcE/apLcVlvQ4o9qpqT7yHUJOr6wYPj9Co
IUX9hpJ+d1zj96Ez5tmPyOzJMD6rlPSSz24ZfUfb2L0oudjOuCAj3sDEVUO8ac1W
Mc0Vu54OJ2mFuAB0FrXtXs5nqiEpOj/J4rUEwfF93y8WlCC9TzwIO3OcxRJ0+RhV
Jg4PSj4qW9WaxHXzB6d27OdVv9Bblvycd8eLohsYeO445bA0cNsOzkmitDs07dUe
bWStbuojDd2ZfNzJ5oeMbeTDmMZQxsRkC5kMN9E0+cKW5/qdezl1vjF7xT/bexxU
1QVNpmYfTCvxsRCNRWfKjfmspmEqxztfoShHIziK2jM+x66OgKkR0i8qFu2AxGEQ
nIJ34CZevynPhzwQ9RPv897naIw4oAyRZpyL2rx5hyGcLbEfFOV1lSS1me8Mg5ke
wp+BfXcB+KToO8AHmHTsd5qRS43XYK0hs9AW8FaiqH+OBU3pf+NIUZ1Apjq+8Lh0
PM4E2sUbaDKLGQAQ/bbOyBXA7uTOmFEnDbP61EKgN2D03qQ+pld0TYL3ZieMUXB5
AeZiFT1Hwjoroaxq3YqlJ+NY/CIkTkocYOuErejpXP8cZTzeSasy/iAc8A/NP5zn
Y3zBqvepWxun0XNeAZd6A347r9+pAhCT04K9dJ45G2RCDXBYvRX3N3U/K6lgJAPs
vedUuzaQK2Nk7ijQLzQJLXuVgFSuJfeO7kVoMgTv3NzOLccyalGWRWY+EbjfAv8o
UaWnfRaEc/WcIbfFMY1DZsM9ZbnC+IxIlIF4jUT/GMjyyuqQEmszD8PR8NNl0r5q
Jw+IxAJp827E39biFQnHr2pOSuAofm3uG0STACEnplt20rGYBMwiOcSriGfTXGZ5
ddVpKeQLP1ZIOyPO3ZeMKsvMsF6DLY1IbSlPOWS9Vc8smcTGky6jhBekNNuTb3Y4
PeDV0QFgZiF5ApRKoqf5aJ9EE3KikOxMaJeEOTrNtdYCEB7PtxXT2Os5X9fwNB2z
G7bBcPQK8PkajRrajwn18FYg5BsE84VRPi/5ggQGvwlKlzpb8dQiVvIUZHAUM43X
ldO7+wGXJjvQuwWmI3YhkwB9Rv/L51wqWeTCjVCxZcyI19x4ijNLPUTEaaMXuxHr
+y/warn6GDwgQnINiBQ6XC5bzvYj51rA4zufnhFHMcbkDLHNLWWrXGEZUwFZG3Zm
qNlLj3M+ju3J7LAqY40YIFx5vlj0GO6gAM8tl0JaCNtOGapsjfZ70Kfjc4iYK9UQ
pPrCgurD8xt9ac2UxeW+uj18EnzFX25PFCF1yhnjpZ/P1TMqdjzq1FcaO8kiSqJg
WWQ/OQQZOCuEb9ShsPIgG1p/jHeFdxWdU2Y0V8MDieactBmdgllTV6DzFUo4HrVu
NuhOGWwVqPNmZAr+tM9vxCTo3g8fWBIbixnyQ0ycPX5xlp7AMgOnZOks0X1O6sk7
9zH70j53IWqQFJz+PN/RYAAUKVAPGXXOJQAw0quOBLADsGDg03by5Dnc5B+Xw95A
ceH9P/QyCqToDybLpOteOg3r0OCzgW8Q9uiCJ8ycb3/ffOkosO9vhm2nNWjghqki
i0vyfvKWFQpF4Z/qAWHhkUb0Qn1OjAnrE4hUPIkdtluJA47GWf+/SygZWVipMhpl
m0tZ3w9cYxTniw5aoSsM6RJLZ7r5fpy8hejfm6U/MvbJiPOtpUbbHASpHvca/MHW
WTGqhnpxGGY5xmPID0N3gNpZKk9Jmd2P1jZ1lwf44KwzIYmHufgjygyvNohGRUfb
BFhrDGqTvVUQcBCQBchzBElsOGZ7rkDvFrKiyo7QvuPdRiHfZbwyMuz5xujVD0kr
bFwWAG4kXf1HKzTQjcK9FEogrsigoENgCyj6n3Lj/tT4rcyEXxfQs1DMMWuK4aLv
rkZOjT54OJMg0/mZ1uBYb90x99jfZ/eSP/XWZ+j8/g6fccyxioRLXf26Q6eA7U7s
pkr6ju3wrEZ7YhJtCfjYED1pm7h5O31k92yoebCICAysT1Pz3be2q8AQG2DmEbBi
RDWVk41Jf1LTin+iKEwHiziAVtSal0dkFkJgQ0KR2I2mNJuJ9Z4idgIiycM4lcyx
/+Q6VbB26phNe24m50CvcFDrXOrsx3YJuDPhEpLMtLhEN4eVrL4F5RVtk5WKIDZ+
XeEboZgKv5POnRnMDkKtEntCrK7Sfg4rPk0clBam2Jy4uPA50xvoz0ddmUK7+g8k
3cx5axzTAOdXzybvzWQGWJJ1USkF2WxlNVooKSdZSNDqFVLVKcoS83bd+JVrCNZC
Qd5wpB0cEAPzCFTfTQvVhAEtWG9JPIP3uGIKV/Wr7uFwT5LIMBskt/2RoZ1O+d3w
arvRBW6Pi0MZdw6Ug976XN1qGR97o0LxfX+EfnrEPyWNg1dHJpbWMzWP0nTIYI/y
u82E0aZFuhJJY24sQmmZ8XVrYBGmQW5JtBnzGhpUlAxQKeDmzx/sttopMh/agS/5
dtoo9n7UHNXGYOoV49sNOCWSsxkroKqrTUaRR2Af0E7TnKNRh+cK0/G7GpHJStoo
Ox12UUwtdDy7xjEIEfukZKk0dkamc9IWnhAauKcykag0+HLmYJDxa7geO3cX1rQw
2IVIpHfAX75ZqZrOy99sCKazSc8OoCiTPzZomHJtQeCEEhK4qO4vLwRvA+WJyMvh
BhQ0vFio388Z8v2bdQErag5y6dX3D0l/jOuXKMywdLs1c32k/iuoy80q7iNgHzTr
lSpXYduTkc3XkP+EQbOgRDRTNFfEZXtxbN+ncSzbhSneMIIughwNUpy2cyr9uIXY
zhFJOdhg2v3kzSsPn1KkZBaWBCY4/ZaV49ruDZDmf8jif3IbCnlbjVlPZcrHuyM3
y7VZ7jCz80WJLELBQSd2w3jiZWCl0+zMpQz0sm3kXpH/NjCQQ3VQbm/57/qGRcKS
yJpOft1udubzcS4VC24GDSHZkFuQARK8hRp6WhQOudsT2xsVG3lKaMjm5OTHmk6P
G1G30w8YRU6qq16syWE1eCVNqI2/5wQFoavuVVVvc/FrGb1C+LZ9CDquXnWBPUFc
V1yb2Ffn5mmNX/Vpq9PkdBsLDFyHerHJirnMELTwZzBQkt9+0gTByY7Enx1P8hY3
DETrARoovnLqcLA9U8EFxkk5+bIPjAm7XChXYUUxJ9TMZBv1zuUp6D8mLpul/WpT
e4QNKLq2bfNJVVufCq6saznnyHsW9E4bm44Sqf4qfc/WmfRbZjf0svl6TMX0bn/q
R9tDkgmvw2INwsJRtFxpXNAjhMHzL1UnKKRJU360ymXQDAwG/NY/aDN1Phr0vCdU
3xvutiouUEwiTEAiRybTQ9ZhsNY6yNeavuRKRVonijVGNutVVlesZLu/WlGGqV3G
S7m6I5gY/E2Ff4gEBxQxu9pa4cyzIbC/vndF3y76wHYI8YCqNrcFsANXw3igQRhc
Y342UJ83GNFsiGQzmlbnT1Og7a5h17gl1Tb1//FK2qbwUKtcJTR3K2yKQ90+zBK9
dTuSLt9TioHvj6/oySZi/ZNJARSRf0khdN533JIdZrl+4jBEzRfvKnZYJBwaSy9W
OrdC9Hm8rduel/cB3sFmle7L1LXN56O6mD0Etopmn/teWzYWQOI2U2edNJWAlToW
WC71cZzY79n/nu3l68tYNtOVu1xg8WxYNIA+jRg9zPcN5vdHHyyFVJVbhAwN/Q+p
+J7XG/HH9VTMQKWdv619RVWjSazm73w+6/adpXBaQmhuxynMX5YfsQg4RtJUryN8
cBTNuDTvSiDgZf9cz94Yi/eD4tcEZ8u1qs6T97Y8JvgP8GmLb+G35DZtQTF+fL5D
Va6jCs/P+gDYFKLI2NBMFRO2s7Uffk3LuvaRAUIVGQliBHtF4oRyuZhuzV4EEO7y
qsV0SK74xVgarGdgRK7BjumK5qmB7ii6jPlx9OloSMOCQQMEOgpZkHwfWaxIUUHp
wObYNWaPSLCqlFquv0MS6uIu3vTD/+78QDZ+53QQrokc4LWYwzCuh385NkqeIxuT
Po9SAqtaqqE7mHHOorxFUj3vedUkqC2OlDvQXcODREUMI+6urFNdDXegsH1LTGQ8
iDJWNagXKOWru5RyvgV50ArT246batpxzkge2zxvownMUP12jiqXMn4FrKnGqQLa
tl8g8O4ut4A3ig61foKLhE8/0vCAf+miuUqQolhyXtIe/xnzw9ZevAIxoK6jbsxz
k10J3aCln1mF1D8wBqmx0xdaS0OXADTLRaoB3zNCITgQtwtbL7HDdDKP2CGAPD1l
y1k41c9mEEVUgDfBBJh3DRPt4juiHLyhuEbhOJix8bhMeWSX71F0HMGsuy8gu3+G
df1arnb6LSXMmVIqhOM8Z2PhcaTU/exUXaWSRrs5bRGkXgn/1CJaUT8DUrZ55RKW
DWjqKUOWjQXs9MD4iNmWThPSpbSPpYAm8UdcxzxgGcQnbI2dOu5Z0RtgxUtavz7U
Sb5yR+ZQ6VjPBE/OEPyOBoh6uR8DhrD/q7ei/yax595gIpmViMEgbRaOb07yy+FQ
EGMuWRUVpxI/oxCTMtKbnW0A3+CNiV43qlR5Upme90KTOnqGlANE8y3T0AFJgNof
AbqRsz51dB0VioydZbA8i9JAV/N8W5RL+i4x77+f7LRsYAAWDQLsqVZ0W4kGPCpt
gVPFXPgaTonXmD3Ix9rLsLYSsSproTqkK3XO6odEkbbGjhi5z0gVM6IzPpb/kjbp
AhaD9YJYx2nqL7oQSiisTUyLn6mpgwPvXKUE8WEbvyDKyaF/3fndztLOIoIpGFiG
NzETeG7qZ/WhQqXVe5FqiwSvbI4zzJzUdY5b45WsM+RSbPsau/ARPn2dOCBwQC8R
z+0Ftxp859sSqdrZ3vF97pQAdx86YefVY5lKoTsMeZ/iUn387YVL32muVeahQy89
CkzSPsJjNEz6D3qvx1JODcKFxqVoSYFWqbMaw8Z8GnawOlNiC15vO7RjMN0IfI/C
zjLJfTCffveq/bDWlutXCcBIW+bWDh5LOPBZxnqrx9N2yPcp8IRQswMjHRLbyD3Z
QZOX4sHDBr0yEEVWhh8jQRGSE7dx87Wb4EFPtgsaXEuPvG2rhN2Dn28Aa1zDdrqw
TuCYH7+E83jugRDhGfl5PlM7odUzqMu3xmTc/gxBzqafuv75u/2tMXt6KDhfD7SG
xf2lM6tAmFmxJO6F3hhJiRUHyZr3qFkB3VNkUk6GkqcO78/EWsFiXf71XaXmDp45
B8a0p1velDhzMSkckEgNvNIwr6Ro33Wdi8YG/xCQdrXYKfttvi+wUTThWbp7n6b1
KpzyIX1bQDAdYCRdKVfR/aM5cGeaxJgLVME/8i1Nq5rP6WqRin4TLRItFO6Cdbcq
azBz53mesGNW15YzcxjfpbS+MlgC5VED62ohN7g8IiFzRcFUocxLN/irKCzPAB5h
GVEkqYK5eO691AKELMI0Bc7CHQK6XviANtKmBgNJEGDqeN9Cd895Uhmw4rsBORW1
LGSoz6Ci2zD7ld3jGG0/8PnDfI3yFquJ/MA3V5KMU48b8mJe+nH3lTu0tQqIg6Fa
JgV3KrY+td6Kp7j29Yr5aYFuBeMevh7YptONmmKRqdpwLWzHbXGpzIJPL1hLxHa0
qD/ZciOP0scfeYc4JMM00L2pYOA2bw2F6MQX9T2XX5KwgwB5y1BNQcHtIykXo/pq
autoXErKmCNP/a7XQfioTUbTEgqtaA6Tz4r+brDbIXWz1CA3qCioX6kTusQgknyi
LFb87s7hDqv+DQjp6t0KDgbzAlXyuVSoi/z8Ik0J0ywI36WRD5SwrKt8MX/6eNfx
qdtr4o+d9Tg+cjhcVLYN58bk8HFy4jBaaQUeS372eH3MNIv0vaR3OpAxA5lU+2wD
lO7wkyvTDw5GZtUx3Uhh4O7PSWLyZfebWa0TT1xWln4tHE+fNLKWiseQk6cvEXdv
UTYAL/GWwwf1QyGesWuPwC/1EFRPs123lHYqsUVrUdn94ulRopK2jBvB/lclKbyZ
W4fwjOxrU1g4JrTsvzJqrGkwOjbtYVF5CG1EdUS4ve62G5HQ/cOjEbwAZNTJ6Llk
ra93y4KbEGcYyOJ+5Rb3FqzMLlRxbhcGUy+ypSYL8zahq3yugSCQVxLFX4+xT7AX
6ltmQzWgJ94T213qtN61Rl9bAQ4WX/hskILCKnBiycGP9haHbmQITMpyNHx/tjyN
nwcZg0VdwGFpgJU5fdzRK1ulA5cLXQjqsLempfKRav9/e97q9H80CHQV8GS6MUoF
hbuBi2OOMhihnuqdh7KAnh7SNR68XgjqWo1v0oroQ/vZPJywYgBkwhgsUOuePm99
4mPethM/TSsaA5Jxg83Li5ZI4J3MDsnG/ajHMrLN0DNMNQBUyForAnlhpEuxblCa
li5ZD6Toc3D/PsIhn3H/zMBzitGA8bBSFu0X0Luo4xVZBA9Swx9MbL5FhvdOkQSU
Q5hON9tjnSqIxPYIqOWtky9rml0qbkxKw0JB5gNRcaNMznAFgn5VIKiRAN8CyyrP
QKiPKFCcESlQdYOH5M4HcPzMeJaoJT1BE2CLzR1V/7hgfhA+VyhWquIRi8Ro+f1j
qTfcs4WsEeB2bFQejyKTvWjpzsRY80PLS5loxg4Pm7AwjZYWjGvNVML5JNwex9Aa
vBllJBbLlN7+vF2jDkUI1gKX4FzaVDk3pUOPc9ilQjaeKdVqXuy4uG/FIQZoBJTX
wFUcCdv7G5+YIG1mrrW+z60eoM6nIhdUIOpEJvUrANbGhw2RKKt/cy+H/yywoWO6
rKcDpmLppygFUlAaetE/7VZuJBq8WmSRLlshT7Dx234MDMxfngWe/p/vIwfsWZZD
3kVs2Bt61gxNifBHUmSY276RZt2R1Mvcyyy4dm1yjoAJyOc4AnyfaZgIaVH/Fs9u
N3iuuLfLkBJMi50bihHWpfFkvX4HClKPHPJAywinzD8pO/EaQgXHGCBtx03Vwoez
kNrCr+2Xn6LUAYJRh9z1cRL1kxxS1Jd3oap4aqMnsTIAVV63dA9FtFxcx2Ij9Ufi
/ZCrF1VZecp9tWc9sKDRLq+qbGIH6M3q5FqnGlylJ/UmHVhDKcAZ7UjrncAUkPTA
WPcyUpPxFJ9+4U7wc15WZ+VIW9ZY7UJEFPfORwCl79ixnQaleBfYB9TD/tkCOw5V
kbSYGx+E5m3mgMo6i9K7g3LsF8TUWj+ONHrc4AuICMmai6xEYqV69aNNtMCpwH3j
X+PaE5MAm9PyTl2YgJlUTPBa1bsHUC0lmfIo+bGlN9oKBexdOSdggYwKTOcltubH
nJ3bORuvL7QN/VG1lD5zeJMTthWpWcd6sXsX4wmd14t4IDAXMqctUfx62I0OIftE
6Z8jogLwFzEsqv9sH8R9zNVFjMyXhnF50Rpx/+QfQOri26rEfiugPwOhTsLxZOd/
jYcFli8O5WZdJx7dmOs42VqNEIMeycs59k+nEA5kc/UwErF53Aus6eNq2irE6gEa
/PfsVaZA8rjZtwktNEvRa69WWlRMBIYgsC4gKNzhZ+7n/cZQMBXkQ7e5+v8KcEuw
QuG2XBJYfSZzJ9C0NfOdm2NNaGho4ldaPIK3myfwNGi4VMZpreZ05YHJT/TJM6uW
VamBGfjFIV1moqgkFBfM2AcC7lgmnhcKHM9GAyOZWfOvBHHytM5N/yW2Zh3SSNGy
gzRDVPvmIVAsg+6igRyltT3uLJ4EJ6SOCcd27i9xPkVtFimioLjKAVniMGHYjAqi
aZTXMHD9eJeSjmrF9dFtAYQkh2WX0jdjkXVcrWhHmRR4/4sliq4/CyB/Lq8e1xpm
Dbolr/CHsz9WDrDGb/0/MVIMFMGmOckpy/Hblqklxhu6ZXzRPVa29nCOl3sMyoo9
HuKXTxDy7TL9USbcp+V9Ly/x1S42IOrdWJFQD+yDaXfd/oFnqukXM/cqySgdzNeJ
Kzvll2qbaamTutpIx2DtEO1lRH7ht3jyvmG+JtWCBwNB5zd7TOeeTJv/mPkXy/Pd
uJjwNXiW0oKBgShqaUMkXuK3Dc8DO7MRi1bA5fIQ02464UeZNuEsI0VXw9SFWNZ5
XHzJRuzVbsL5/rm88aoCsWP0MeMMBr+ey8PdRMWWoHsWcOvt4yvg36rsnTYpD4FO
8ApNj27wWol9oto6Qy30HUpuVmfhsNdqL6dOhUj4EVDej/l++F7hBOl91F2oA+ZM
JM1wapwS2FW6AuhZwJjdL9gwAxc1H7eI/BwpiIFq6zf4Qh0MKmGpmN2PyGeNtfmq
oDqi8u3964ZFZxwF/s2I5wwRhBbPyAt3Wpa/slWnTFXzOVTKbQ4Gu74+wttA4bgZ
gMNZCTnRpbeypf0XmwZ82bR9caCSOnJBL0MqE8OK8dE+uSuR5ycWpSySc+g0tRqV
v6kYWsBuQNpyZhRzDEeXFNvyZMVwcb+Pq0RGuVw0mMozPHv/Z+A8lHg1qXEJvyrH
qc9z/Zzugrl3lgOYdx3g83N/m4wrZVhKQqLzEf8wohAGoDHCE9Y9dKC9PWXuriE/
WbLLuJ6XzEQO4hz1C24YZnjnLuOYzx2L1aC5VexB/3FTUiBXwTc3PpWQyYZpUXRi
uQYJfSQ11Vq2w7ogcB1kGUlqYQECVk5Yx/rDkGMieKWWOhtPW/td1gyBqReNBpbL
GNZMc0hlty/Qo7wYfrQb1zMoQ3wjMaKAjr2kONxCNivE/enchGgv1BxEWDYJOVci
Jk02IwPvYrbpCVjoK0L3i2cu6nz1typN/BB7JXSleoUS523zvLiGeswL/Adx4WUo
qBCXpB3rlqoxyqgs5y30Bsn4MpFYW32zdrssRiacWchsHX3vN1ln15urH1d8AdZr
HSNZXVA6H+OrHYKcZDsek/6bu2lX50ehMatybPpGmgxIaxrd7/x+YxlWcu3FwvtB
/YXFxn01R3a8rcP6OnjID2HplQTevivjVIJ3cPNbFku3IZ77A34t1m3dWsSX/nXL
miGTdsDngzQMnWI2Qcvs5WtWlKFo+m7eedCiQ8eMVcTO7vLKYT5Fa5tqv8SUeJsF
xH5lBA7GOD23UbrxHxkfbHMGE0hYtQPEf07oAAgrmdno83JBuYIqBp9ffVLGibrr
PJ52ZbsWfvCy5aIJ8Fi0njdu8i4Y+G/HpYwn2pLyXDMXveMBhOjcnTwiWQAmofvv
1HbNNvr39InKIE5Rn0g8yeE5AyNkKZI9XU0QXGz/jKJue5uyLO9ZnmB59vm6FVqu
9JuNmPRj8F4vSWh/hns0Vql7ANqt1Or9ckH3xv9yRkHev72Iew5LLdmRq5IKCkkq
jG6UUjOLuUOCltmeIs8d76gRoYvjzfqdRGOMnU5lMmjgURsC8nGAplwTpsGuaEU3
qNk0y56plzE0YNdyZyHCLEh8vomonWIETnYs9H7ymc4sIVrQDIdZXDEfSlLI5dCp
C7rH2HENrGN644vUD81wIwByctKaQJXOK4yIIOvkBN2TNaSBoIaD9Ogo272eLqqS
CXM7OddajQdxqZ6IiUosJs26h8J9GbzmpdiaDILSRUh7Nmv+0a7lHFntKfPJ9Brn
rS+mrb6Pa+cu/NnemFnpIV4QtZpOEovCM8f3qwNQOuSI5oZWvVKM60QhjH/ZHoxU
Rwy1oW3afDc8Oelfl+ytjubiV0JOOzucMm1AbZMyHIBIKFFYiS/21ULLIImvnAwd
m22mMqTkvKOp4OfmHPN58D6U+07TCWx/DixBwEEEK5/LlOF+r0kP+Zqw61B6AN6B
wU8q2CMOH2DcO9jv1JNSSwyAcY6/qPJc0afOZ4uFl7noFT7A4SOYCXjqBfRyy8gP
NYVa2Zd024qYeUQi7cf2avLa5DYksP3tAle2MFouMDMITe2lG39T/ZFt7rjc8U13
A47QsXUFigU9w06uwTUyOLF3OtTD4fgEKNs7g3aUm/KYBvpkGddLD3NHaReLdUhN
tQMOjTMdbrniSSqebuOXK8vGAuEzLChxRxc7DpNiuV6ntNJmsfgNG2guJ4v2Due9
QMGVEWYQNLIsSEed9kHaXUesnjRGBVo3GRJNS7KGTZjnd7Ayk9uVx1Kj0Ncb1AAP
YZtF1zkR+bixYIGmoTNydtJEfl1xlneVQKfWlsBTEvxJtw+zB7gwUzkDOjUAIrUR
Egacv7328bNfQnS9Ev+KQAFjcRDavaERTqiX7bbHwTySKwGMZqWflIYXLheiji5E
mOJHMyblNILwOCvFrOS0akAtoLhExmCD+XdVRiPCGa5vVdh8kmGpTGtL76QdMBLe
r5C9qVF1mXutmXmZZ4ReSXlwJ7GqECXvVGNVg4+mVsBY1PKJcwTKo9c2wvnyOjGH
2lHUI88DQgW31M6udS1muRwQKBebFPaM6T8LGnJ+i1hZ2/HpqJeGkSkYmZOYwn/D
AyH6SPi9XG4HOqoZdBeIjrBz9fP69yGBRhQL3gqulCFGPj5W6V4IIv6L9e9P5sBz
EeK8BKWOPPSeDWiSw9odEfyM3rxOXCbj7HUXi7qo4YOsfpJlLMCyREZ7Jee7S+zW
B1c85wInBztdRNjvntsOhhEAQFwLt3FCLMkrTf/n+mErRypUas/iXyczM8/HjUvH
bvzBxLv4RGf/aQMJAOOPxUG/gBHXLA1V4379eucy0DSBjdNpAqd7u1bpe/IAmKPU
0kODg8+wj0QkUzMILhc5dO9mUjs0+QWtlInPz/dw/lwQGUnS/h1j45OtpsKIYODl
yFFDaJilhbsRd0a+yL58Q75wQn0ojvuDPJs5zhGITBcK24zlyrBs54d+QcSv4PlY
mxZhtsKhrRtfqD3BBW7IzksRdZspff5OJ8AcWkj1aMot/JfXPtfT1YNu1hiHDZM7
wy5DKIaYZu9U4cFtCr7QgADrDgDzO2BNz8OtiFQYEaCyL8g7Xv6m51I4z/kpOgaP
Tgmxg9EUYzr5SI7tLFcWwRuYfv5Ub0oGLVBEy64oRVDF2zdPW7D9+RT0gx9H7olH
nvElGDlXjuKLS8gEgNFnZOFoDVIMW9oYQbPgLZ4ulfAmPcNStEZOHn3NSNAQ2Mr6
x3DtwVBi9F4ETyuX2C1l8NElCAFHDIG+4LeF2qHfx6XiHAeXXqwKSj+oJ2UpuUoy
Hqg3OIP8jOdb/ebZwgSkWlvSAxvc+FCq2JM5QRbrIXDvSBvR0kbn6vnjqD5xEs+V
unqxqwRpShBR1eSFTvimqVCG7CPK9SdS4ycwAfD2OGja4C08LXtkZzUAFPq0qITO
8TnS8KKc55v8I2cr4wQKxprtKeOm8agTxWFJeFa+VW4ZGVjHLCmq7WCXV2enj/RN
7TVem+YzbHiCgvrEPtKgQJ7n3X2unzmYSPY3wo34eZrwllvUu2VJP0L0cgz48HwO
YrFi8rx1G0lgYzLQR2HPJtp/XAh/pj/1FzIdWTZwBKEmyxrFiNcwdiNpezveue4h
h/7eAo2THEMa8amrwlSXLOXWogNsRDTQGiTvYTRiyWyGSxMS+esDuYK0QLjUrvTL
4Q58SSVfeRPVtfSmmvtr9W8n7ONKmW+z2NlENnSK7lIfaGYEK+ZWJIg3cwryhnHQ
aSxYt7i2Wi7HXy2k9KM/a+DiF3tY/AmrZ/3eqgoD7CzI9xHqBsmknXyeqt9DTQK9
sHhbKXh9ZvLzirgutUbr/cIbKotwOu8riLFdvq26CHd+6saJ9/2ve0kVq7CQg2yF
iGFDH3RYm+dwn55mJiph9STP0qXRXSGzElJxhwETvQvsAdU3GzhNl86pboks/h2M
/NRUKFBdElSNrBZUkOVk0k6pWHPkruRoXaDEU0mMcJud3HlBFCOhISTCXG46AChQ
pQi9MIgTDP6yOk++i+oWCy847pytIo+o7U/XdKPvM9jkqorduLbgmMxOJ5iCIUUd
x6Tepa+k8aVCtlfOBRdiu6/GvRcxeUYXsmYDkVbt4GUxGUq5f1V2vUUvELK24Exo
6BYHFQGtYlp1lfaw+4ryGpPsRlslU9iky2FTADw68DmXi+g63FECMVqNOD9zEgQ2
++QcKYhQ2+VCL5uzU0Mc8Dg5aQm74TmwOkz9M2u8W5u73lxKLm4/KYa3YkjsfSuV
c/WJy4GNaCB/zi4JUPr9xOIBIRjnRU1WQjeLPw1+xd+wmx+Xm6u8d4HCWsUwTq+Q
6Cki5N1Hgwfs2H3gCoa00yudnJmBfFTebcN2nVMbcsRcLaNqeKYrCu9nr4TnC7Fk
dXD2t3DQlRyjXz2gC2c2QlIbyLESoAM1dXIvwC9ZBcDb5wghhWJFNgGc3EmFSHta
MHpYTLaO69d8HEzyVXStHTxWZKSYM9Z8JGa7Oq4W9rYDhCEhWgYyX/myF93oy/2A
sYkfwBK7rdSkNDrGHM8J6Zfyozpjw06LOwRdCcQpmuZ9g02xUfZ9QOiji3/O1too
Kh/43wLoSgvpZwCCNyE1eJaVehcFPR94eZQPbqk6ktfJZpDnT6tBU/+ljgWOXUqA
Wksne89y3HzViy3Vmh2E4fY69nZ1fjRviXAeSaUASfrOQFrMI8ImI6D6RgtC4CtS
UhgVegiajfQC7FM++ToGPReG/jJT4Q+Ux3iNNIQk76kHml5vWR7cWXiH51Q5itHG
EeHyOgGMogNXc3pWfEjkXnTf+tWFaSyQq15jAUg2NCWP3yzMDNrDm+QObqyiGaCg
9tLxQhL159qtOCBObOT5eOaA3gEppzj2iWhE49lC1C6ETBkovVuVowomDzd4eiRH
X6tbMdBl3JiQB4bQGGiV0Et1AsmqGcgv1QyZiUFUorhD+xTIJvbwoBcxXmxd+7uh
L9NissEGuMYvqgg/UB/nxha7m84Zf0VnXg1By137cm0GEaTnu2l9IOppkp53Wbzv
gPz7X50NBzd2gCFrhY24WuseaRu8hbIyIeBpuj38skYSN8bRLLABM2gogxrDpQiY
pzXT3siRfpv/a9cPYNrkJ7Gf1tQV5GuwMYRei90wI858omsoMggYer9bQuo/gInj
0DowDUqxRLmanqZnkCqeZb0QrwTL1pUJQLXlsZzKN1YJq84wgGLTLQhtiuhB3HUQ
msiUv0AxCaDw8+XOs0aVNcx5OVS5s1qY0vwzPWAsa7bzfiEJXDT/Ews+Qvxc/ivt
wdX9PGssHDlaFrM9tUHqNgN2yZ8UbM3KsZKMjoshO60bUPp7D0wQSeA/dw2dNN6a
pQIkVajEqb+AAsnOLqpqxoBM+H6V793bW3O/XuOW0eVFwB/S3+8lb+IStz9kfeSK
0H0E+JtK7gIdfv7/Cm2tuGDYJUxDOSiGBBYaDsTm4cWKVEn7zq6tE7WT0UsfEk8t
/WmODicsfRl/RvgfDkTYTje9mrpPe9MdeKC01plgkrssocC3wgCj6QRfMTsfiLtV
JUkGLl7Hmj2l5uz0weAOAmkxGT8Kc/lwePjC34WeRhWD+vgKGRI44gHocMJ+auOI
BB40Z20vhBRpn5VEy5M6eaxFaOR4u+ie6BcH7gh3JaHVLVRjI2RPVmINtfq5egOW
wuYEz4qaYoJPNQegmMn1tL9fWOd8O8TGY3g9qpJq9qCft7YuFIt4UgSKJ9i7QyCV
ofiAdG4DHsTAN/Fo65BmEF6d4kQtcpugsH6ugqg3Mrh1gTkATb7RD0TP7cerDfZr
ll8h0JU8LaQr4yiK8UoIqRi6uC7zscVPpx5n2VaY5opcNjR6fDEDHzHVZyqQStUx
IHgryotwARoK6d0iSfJyg3BQUYzWJuEp/ZHtDc2NLAsk8Zo5TQ+gXyF5IXRb8Rcd
brG4JLIH0IpC/ZblJQtKOACtFnXWot5QzU1b3PMFeV2dL8x/9CWINj5+EvBgGIdK
wR9mbBgBoXb5EgLhhc8tSgbt2CUyNkpN5nkq0mGKeVWNDQ5OumvKklCBdpu7xW1Q
NHV+Ijr2Kbkg3D74ZQ7/a81l/cjUTPIlTfa+yEMXcNEnGeMeXZ7adFy9RreYlC5S
X7Avkv3ShQnqnONwun17GXcSbpHlrlkviLSmvfcW3DywZOjDiUiTmcqmgRi72uzM
WZefPsMtzsDXqYFLS2Cos3ORSu9T5JHnHuKCX2apO6CTD1YHj5AJUs2CEozoP8BZ
6wIdw2PFUeRWvXmdjo7I7p63jyeaez2Cx76qg9uZvHNi/6TZfR5kdNYrb7xH+IP8
QeG69ew8CHLWqBQH9WWFn2hyL2kXSU9zSAuGk0UGEdznlsEwn2QRo02p3Yyb/2Tb
7OAqhma8+EifKJxjThg+BxsYQPScQ4lbxnpNJNccRPwS/Jzr13+IpHWeI8lbgK+t
W22+QewogVqqX2mYGlXJ5+qr8838YdgjsdTqhxKG1DvqYO6y0ztoJoFgkoZtTt8L
34Ylg8TaQQw7DhHVZbnVEXGrhGUSsYH968peWK3fkz/BJsbO+bDifwuibXnyvTH3
XX+cXU52TY70hRDjZ0LWNu3aEyvQkVvHDSs0/jygz2RON2dccAYehFy0U9WLmRcV
80qx0Ktu8SuIvzoXP34veyeRnb1X9q2jgEV6zUr+FNV7adxGRfxZIbAIcnAFyjRs
nmhA3uFaAitzmbwHrx/80l12testceA1w4g4LA/JDURQu7m4G5DncH+YfJAYEsCf
NvEajpKbAJZVFG+a/kU5WtElVu40Z9m7DTuu9uESZuFso6yhW9CNKI6W5k3I20Z2
CkwPqLrCSLV4ILK8KKqmt3nuRkVSJDatK9BwEikqOpd6niyLjlm8wNa8MqINx5Oz
c8ooPBeK7kwJA0zlQk4alkwgooDKMxcIpIc7J4Xh8f19Wbc7nx+iMqWZzWYTnqmb
d1xmIfrHdz+59f/wzq+Y67C6k7KvHt1sX1fY3vY54ip8yx6t0WuxjSPfJNraCzbK
ectGqMYQSkLBrkyfZ8Fj2fiig5E40u3vXBelbi2TNMxgs7zGDZYlhLugHqdiDc5I
FkBTf/Ny5YPKSj8nNdBGO5a22BJWaWsyshk3fmFyPstkv8Cz/59uDMc6s25mcMgt
OWt5Q7wms9evS7jb2rR2+t6Y1fyRJ62qkR6XzSrgzgbOaN7zMEHmS6cAVo9e9Wby
jkxU0efJtVwzA6wJ8ZreiI+hgRr7NTdqCknjD/+DBs9woGs4cMVH9vI1uhKqKAY7
KH9XXqAOglfFAGt0eo++sCfbEZALBuZo7G4fsjFmSpmMfEHax6BRSzlkfcomnIQn
EHDUS4O7j2kz0Qys+2cNRJqxmVTPIFTc7ZsiPmpzcyrTm5c3FqEAUYBqM4vR7+Xo
H0BV+NGfrdMYvcB5+3/mpl0XDKeDFqMdvoy6WOfIgoJvkdPr2PzfP7VByc65otyT
BxJpXZnH2cpYojVfbml6vygsyY/LLgoj/wEb8qyczFkuMRi02pc2Uv+reV0LHJi7
hxHwgFXdYnfs4PcmbOvVQTSsEvS09L7sVAMSZXk0wno9S5L4A1S2FIpO2Jqyg6yk
+x6z2GjwgCwDaR2X+SW7ZfCYzwpAg2XIRm+F4oLnVp/3xpsWQTB5MPhKyYs52P9t
SaapwKOviXM/+T08QlgRfFO6Yb7cWy6jkfZ08ePSHSH9IkiC35DFocv1XRLiUkX4
a3K7X15e7TTxbA9cMqgDgNkFvmpoRW0BbxXJ3/zu0pKuyrTQpdNdYyQ3Ruum+EH2
9oFLYTU+fw8oWDJu6p1MTRRhRljB5WCjhXRG4hsOPscPfrAjQ0KQLSCUJmz0qoxd
1WTPA32937bWNVrvk3GBtrhMfbsKrtLpM3z3KLex6rMzmUmwkrGSQN9AkyAZIoB9
hia1477ytDa83BXnE2po7xNaWXxg4odNCj8ZVXzzLT12+s3bM1+B7KbW4m5Qs1CY
OREG1cj5AlsKUp72MvVP4/ofB8xx9XlsM+Lhdnhu8fuo5OQIq7wZmJlCW8Iai6Dq
FQHMbl9Keoflm8Uicyb47hCwOy79AsDWHcHMbkDl9xp1HkTC2qo21KUhF6v+Ptj2
miTwvulMZAek9J4PZTnLVRTG1ADmxs1gKjftLFDxyU0Ity9wto8Faa4MrKu7oqNk
ZREtoadpgwvKWGym8KHknD+qnrgbZrU8c7QgPnBuaNQ2oLjipsZe56fe5XT8+jOA
TScLEv7+Jh12sidtkVVZZ3J6+IaZS8wAty8qRpaZUwhobkdTNPRSz3wuZ5hHFOOK
RfxRg363vyNukV6T5o9WlfFHt3U0sMjeV3x3nMbV7Diq2wncP5pR+H5NOA9UGCXY
64n3q85mp2UhIPiYz6XXU+RwlNd3VBWYAeTtgtTvtfVqERpBY+Zxp0/f1Ctg+lNt
FZBomKnjlm+a3o6eWNf0iUm731GcO+kIP6UfZdw49XdwkX4Ry/4iz8dOw/FAQQQv
cDYnpdQxJTPkTLa/FgWuvur4WjMppEBfs+hNE7LFOsZezxFcfuWb0mrw6Xfyuhbm
hBXMz5KigiYGq4lbcbEojrujNe6QsPvvW9cRaQGMnxcJIdWZ3N+KEtVTG8VZ9pVV
rMNeN0piGVIFzt8vKJvsaaWR8sNCzNqC2Z+1TnZLt2woyeMmnHd4muqKiOv8EMkU
3n+WSAhDGVx0mRcs/JqFh5iCfJfiBsvATxlaD8qnFVE69uiqUNUcZnoJhA1DDOHa
6qxvha49ZYWD+jjP5Rda68EqqW+r2gihyKTR1ybW5fCJnelL+JVFCiFL6Z7RFCb0
nOxNsGXRo1PGhDh4ZS2gNlDfHKMkSpo0641AmUGrHqyELaRWCanzyViWkmGW/Ye1
eTomeIguvqMBj0dklnqj0fmcuzAJS04cbGEAl45q8mxpb8BADDY8O9OajtyIu7QK
2x38HyJ0YzZW0q7kBKmSm1LpEIHiPJUSf7lK9G7nmJ8akLc3B6oDARSv2OVAw5iH
KeBgTMKIQsBY/AqxDN6OYSIlTAfIaLFaJn2BWJXEBG9kBYyLc2YLgTBzU+d6kHQ/
fEMMRNlMfTw1kDdJytwPUXqJlHM9oVkEaMYSm2/QHuOXlXSAahZO402cOdmXUcn/
hCRC2UbRcKO9uF3qnsIqDMN9cHDAxLaqXf4wC9NEA4Y4we4ZuW+doUc8cmEtOgE9
9Vh3jkr9Mh6Esu5S1P2FMd0+TTTLveLHIahwUSZIJngG/1KVcCc7/1MmoowGJkkb
2frLw0mragHqdR+MOI8BCuaE3wKmbaDJF+WT8AtMhVCKLuyaxICf1Bqm9k+XkUFU
Duru0YGYVUXTS65pVJcGWcI4jgYUDkqoJrr92qDQjVjyLNaHLEcKdz96AQdnds1W
RgqJuKthZ9elTinAv+WG0v4JCR+gP/U1LbB5+UpDy6d5pRUcqiPZfYbIKRZCBBwN
u9EKb+gDcC5AOtxzksof3nPPYp4RNzq+wPcFHbB8InM6/lG1QaABv1YlsVJ5iCSt
V8YWRDJl6sU8ykmG64R73NizPS26FbLrjI0Sy6Q2tVESLT3jLu+xIclvF4nC8FEx
EOFtNS+mDd+fwdN1wChSUdyXtGY99QWozXvppNkg0ABBL74n/dKuEYBiHfhlmCt3
f2lr9p8YtFNqx45KGZ0K0+zeu/3FX994dnpjrVHBjH/Pbo9/ZFXaBnX26nhwiPI/
faWFW78sH0++JGTm4ARppBR73M9XoWFvkTSTTaL+13NHC8la/1BIkJBahEO1esoG
ucGW6SHVRGaQcmKhwx3VOrz6TeU79ZiywWJ7lwsHMwoKQVQnGMhhgowpyWmeybTk
mdIl5FqA478PyJemfcr09qVMT2eYFdXrokpxdZum05DXiAZiGla5sl0uVZV8BYiB
HgqeTzYc3R9iCOhDR3vZFWGeOfR75G8caxSwy7TULvHLnKSvI2KXGsLfxZX1vFeY
LMmAayIBO1B7Jajl7Jt/RbPZ8sDweg1EjG230/ZbtT+XSOD2IlE6hUlvLZurjz7H
Xiz/p3TNIVg6glge2/Rzd5eKrKsaKZ12TbvoV3+yr71+FbbbUnXMomip8dxAutCJ
U+6TgIqsrMLYCNMjAvMfcPbKDKx+Ek0Ax7Bu6Hw5Hy9Jr+AU+R8WO5m044NkHj4B
jEFFSiOLVNdmIQ0/HKLmKeEF0IzMvLeAme4+L3uqo9y4TAUbDRzLj/CWIYKP58LG
tScbdaQ/Etkm4tAVCg4FZiMtl5/BcndbVE5L+G8Hvq5fYCnOz+XXvdX3BPfBo4V6
dqZ+Q+xnU7/fao3Gv2zmGqG9Basma02dRfNdKJhTo46kmynw4n7vHzvzSNqmn3gc
k2FbMz0L/+ufOO31oIzOR5l1acj6U9NSsMd0i6KYGPBj/HReugeaGXTo6exRMq15
SPi2rP7xVpbqXoY/ZtAQsZ2n1Khg0G56+f52ZDMKT0GQzBcaRq6tfxdbiBuh0lxD
ZKU1jfo9yYaGb1407l1iZTn8sV3tjy0XB6kN5XOX/BJsDn2IbXuxxmJgMxKh8WWk
OgM7VpYqf3SUzoxn0MjuILpL+/kDR7rh7ZJlFUPNErKoRbVHCR0Qy0EicnDg990v
KTIojetDA7ZbIjyx+1ubv2ejfQO7eyzxJ6nED+ji8JZrtZejXhiOLGXSHeotDtLY
OKtRJMnXAGMDl1WgGHEemhvu7MPEnUyKkJxGiXHfArs0cfp9PmU3S4tgZTZXaxel
A6H5XM48uirYOeWQGgM45sYMoMJIbGVbyPbgaHaiFa9Ms8loAq9+E7X49D5qMMNz
7ikL4FQtwVNE6IK+Pj2uUE/jqE+8Tm1H983i/iVtO9le3qWOIlgU7xRoeDU3/WUu
K1jAlq0hslRq7BMlJo4FkvY8ASj81KKuarlCM2NlLCjvfTOlfbzIBMJvoFS4v6//
3zln4kF4PIZW26PYR4tSFIHCGPXEJeQernkYSWg38xBKxI55H28lxIEUhkbl0XlO
Ac2FE69tL/LQ+sbkxX6msKj6ivBnKw8JdymrVWWYbq5PMIRbi1kRDvnRUKAdT7vl
UeW0RD21LvNUwNvVi4srzHw8ujJwjCq+VaPc2fFk7b2ByDr9SlmBuyjXn2qvMvD8
BAjHpcCcKpd1EL2eVF/rnHHrZAZjsKphoqMmgEsulJFAR2bQC7p7A9+7pqRF7tsS
Pc3J2uNZcpTTk7LInE8+VifHhh0sGrNsxeeLabTWD/njiIj8YbvWrtccBIJt6Nkg
d5DaJDP/Kv+iR6zuQh7HMoUmW7hplZ1+mRQPk1m+MJw9fWnQVHcTYCcEmOFqa2mH
B711+NbH8Npwq5Dp9Wx75tB34wREeU0EARoj5mGrtupCahsHOAHGKv9S8r/F1kSs
/OpeEYVC/dU4H4J66BHc5DaWHgILuSZ6oxvKjO9o9i0YFrVTIKnLWpZhiaSgcpdr
jqn2svdMkTsqM0TsfpxAMNo+9+VbEOnzXbdB+FlMKYo8hg5vMITXwQC59xCQYpnZ
rPmMZiKnSmaXjsuNFKTxz4PJRO7xKiVjkeH5m5GOmFq819qzYGdTc3EcNpNKY29a
QamDFPWaRK4Ku/tZ4iDXiO08Eept9aV+LaxjXLuY8zXcagh4aKAQ4cGBb9SoNuQG
dWuAUWrcKqzaCGXIh7A3AVBBxkKgIXPzVrKk+8GQavX76NCtDtG8ALS3U30S39ZE
x78woDOjwOZJ7ruAxWwfYULgp1S+4geIdNXal8iPaIbZTbRfw3OqxD7i3KaOMC18
CoCw8Oc61e8NtPWTdHeM+c+7ksYadJ0OLx1LJNFXRmko7sKOv3Z8plbsjRkLPEeK
zhFyBK14FlzK8QebCAQSi6Rs/dudyrZ0MVfGwPbcfJpqylsQFtLilQoqCOcU/S3M
K1bVIvc3dH2kh73lJ8Z8EMfeJ7zGn36diJ5b/S9EarSBkU4n2cfLpxq3pjpSMp10
hg9wTgvN2x3c2VL6VCKwD5uKhixpXYNtv7dDSP8tAgZCNvCCwdbnUGhhV4+x1ZaU
5K4eXky2cv4zrGE2nREOeTwsjsw0/eQbjJtYrv471DAmbEpX0LUjDyvuBezCsczh
e59r/9LV6E8ltrhpPQQb2L/RnEBcP/2kSf6u2++zZGZ6QV30TNyzrK72dUgkh20p
wSGglXe1L9U2S1ITLB1nbMk9kDbOOcBpbw9+ciO6zmPiWUUwr9QQJ8e1JHeVWuz/
pUsV9jcidFHXDplRYiAc1vaYXXF1xve1cbSQHhvwlNqRX1LBfa684DhD9/17EGYY
uji4h2gKYUQHttRLzC1UcamkNDMPa1tPTBJCz8V1ngLKedHQ6f6pIc5JD3wgbTop
4nIe8lAe1gGkkJue80OXbuQ5G+97hOs82LZm5Z26KTA2w/n56qWV1YAvHCMoUHgz
81jh4BKYtrNApEUwwNCEZI9QIjhajvB3nGCGt/+WLag91hiVt2ZswZN4vrtPpvex
Snh4TVLT9wkarrxmmiCXxUCJpCoFK5okQZpbXDDsgFk58ac+P0lzFhsmZcxQZgpR
vqtpRVSMuaMzcQqZftIGMd5qT5t1nzgo7oSNKDskWNkqKE4LgPg+uy3mMPLVru/x
oqmTbVetGFSqUpJ0rBXxlCPsEUYDdzs1TV0nD5U+YjiC8ljqAZDm2ML5SVZKhaku
kTEZBWHWdjkzBUSxNNKERmNT7OuHS1lP83Z4VPQZfejR/PkFZtw7Xi4Ze7uC8ukc
43+V87UTvVvSGTfeZR0Bm5HXCdEHhPDYnJTGsVy3RkB3PZflRMQ0oiavPWgOIAtd
o7SPk2cj4j1iBPqMaMSn+Kp2ysRnVB2vKt+7GJcxxLPnqunrOdL+X887A1VRbla6
3tsjjw4cy2S1EnlTT4u6Vib2etyMAYQ28X+MHo11AyrI67PqtP8bu2IdupneuEy7
gndPuxUen9A2Sz38lIXpa2qfGWlNJdWk324YWA3wOscHu69H/ZF1N80M6bxfs+nT
clmC+eY4SKsHABdQEUeEJc9+3IYuaby9hGYoQxjQmKQasoLPSoIGDy6pWgwI/2wX
2RcD9ZM7uKP6X6R0Fn2+ClTnK2tf5PpAtqnDoXjXzVwhIoJwYSMgch2jZZx2v+3f
MhkUSjQhKjUU2WkzomnaRp6nDOWjnA2hR+LeZfqYLmDq9klNacDK8TCErjGGF7Jw
T2LSxAIQv7Oh2wdPHigqxfq0sIcEw5py3hTGTWaEDP5nSNUvoIgOVtoYSuMf6Vdb
AftKiQ8tx4lekkt5MqUfzpiZLkbFEgXcSQoMMLdhSYoebymlASE4G6qLXEK8aG/p
qJ6JVECdOE2m7I92dhroQryggF1sk89OUGcTNQ3Wd8sd/ihqXoXfoXKYl/EJNjYk
WM1etIzMZinykX9o65A8FQAgkVRGVUoFTerv+FWF6Ui2cRpUnNMAr31xqTRewj00
rFQaZY8lbd5fqBxFOKife9CgCytzxPHiydSVhDUJ+onv8SPa5eXE2cXx+Za/cd05
m5/QJEVFtK4m29nWPjD5AfP+myntuoQBRpt8Ts33SEQD7iWDdGpCwCdOzqtFW8nW
qCQLjrytBYY4kTM0ozJUPuoyhNJRdPSOKWdNUla+rnmR4/mw0MbZmdFg64A7E2sk
/SHBH8PxAtei+jVeYq70gR0E6KHISxWSMuju7oXdR3hBkkw+hGY87yBgTn2X05lu
rqhUyplezUUgT4EQZEwLWt3csW/iLhfU9YV0db/ntXknJxzuVJtVQ1vLHdZ5V/+5
X4yjI31tf2XLtzxf+Pi4z0fc7WuuhHR3XI4XeF6TwfkhXSjjWcDnBIGks9uDUw6F
Yrj5gwPF2f1OzUtKjC+uiGnRgs62Ce+J14O+zSzFWymZLi54f1shI4nUjiaAaK45
9ejCp221da5WctU+28bOZRECnWG/DT/03lHWnFS/UGPxzg78/0AGsVZP5bxODvYu
6nUO00jaVwqUJFpMS01HPNTA7yA/+7WvYtaOA/W2xVQU266GTIIrfcSSw3ZmQ5RY
afr6Yaus030o+0ArdViK8CE/4vE5PKd9T8XglYhPlGuFBMZleLWJiTiO9YGFlDT3
7VobXuoEJEKCyV2VSSZDX9YEEZYZnuGKjUqiZO84XaIVfxpWI0KgeUwK1gHTu+qg
MLsgXN6kiwqGQHaEG6VLjndSOJkeMKe2oZbo1O6RBF0xs9y6UwOw1Ux3Q9MTWGLm
xo9ElsiYfNZ33MX0FtvTXIGHhAoYChMrcubBPAfm7p7pG2V15v9zi94dT5y4kTeU
bjJdtq+EVKBFwzTOtaiKOBbComluBh5PBXTfnquNqiZBLOgcp36kgMYjGKR9vCnb
lYbR7ChFXXPIDnNV/pVIxArsTUvugv2TQbteyh5djUwG2+0Ccw/1IzzdfWTOmn/N
os1TpXVg3/Kp8tREbPKk7eoHvNnSs4fRcpBSWTi2OT8DKdcdzAhoOT2sbeqoFZwt
tz6rY/Y5IUBca9Kdunbt79XBT3rEt69u8pq/AchZHrhOmVGtK+Ptv3ZLI7UAlUfd
h0vt0y7ioF3i12qtk8bi8GR6EyWtDhVm9AOGpCnEQUwDUXiIupe/tTCrId4+jqgC
IeCE6KAXQDjlEyCpv6QkBfnR33M1y5gPqYyzg8dtsKO2aWyUAOwpgCfYqFGsZXj+
sZ/XwtQVgxTmAOmjoBFRYtD8Fdv9DCTv0B48Yo/lVxJ0N/smZLb3MYeMNj6XgysD
5Uiv/tfAIzimNjF5BsHGgJx36JvKPoPB7OIbWMtgc1pv5tWFlx0cluHSPvVN0Lw7
qKvQbRpMIx+OG9pk8HNXmR4JH9w8OJ6v+5yQi6GLd4/2jYmcUKyjNygSSMfj6C0j
v5xYypEzw3/BwifTMUhi0SZF/+IAt+gE9h56d93UAKBueh1B/FNePS5MbfjRSFMb
hbB3wD7UPqXciJMPBQHTNR2GB9ZE4aJ7DF6EQk5cY/Zfh1atkboVtGuuQfSIQRgE
jJA2YJTKYv7SmtWtaEr6UYYyW917whDQd3cJPVr+f6ie9ApEF+7Vr/6e3ZAddVz3
kmt3G7i0Ixgv2qEnulyXw5xydK3ntQGCZWhngapuv4HulCfgnxWvaCGaSIiMVCm3
eOvuCU6yOEZ7DICd8AG/Sc8fnlvE+4mziQIPxaeZV0t+RCgfozuENDYTb5htUgeh
W/PtN3of3I2JNnMuH+4+T/AmdmghuuT9yZ4cyLaOu4nHpgFFK5EpaZZp/i9/APUs
5sZfW71Divtl30OOPNtgcOMG0oUwxoBdQeRMhW3bpyje51Gr0YWQJl11Rz0OqQeB
NpO17niaTfUIF/jU0S9cO+6COOfJYYAWgUkSZ8uGkiNPBIOooOm7nLNdfrobD8DW
E+6aA/WzIju/0e52ke778yjHcsZGQUlScSSCukZGGo8jjKGmGfOMN4d5/1HqRo32
3k4T/I+5pQuaOkjU/KUbYn/dAYMEYZolR9Ty5IAGlGIYlaONTxQye667sLswatJl
GtRFBprBimOwWGMG1RqWU5NIbabDNcxhGsMyHASrH7WjrwT1ih+nOPk/yNocsBvE
fXRGUPlm78In9ptHxx3zZt5PeZpG/bg/L1zNoYmH4K7FKThmXNy3tLt9m2AdbZEd
FN7nY9ssgWR4iCuyZnvQPplGVDLABj5EmX0enAhs64WeQhT79EW+YhPbVLMlC9IP
GJrzgl8uHqrGKBrNvriescBKnD7MAa4KAsklCI/Yul9HikHDAn/bPsi5xyIOJCV5
o/zi6VxOpvgs3pk7utSToN3U0IiVbXC0ZEu0vufp3/J4mpgxAXWQFKOT+RtXDeqM
KwEGzVmpDcT//ZNi3iUcp5AgMBdEBg9EZ+PvOMsXwIFWsqY8VWktIEEbBwktJ9nU
nDQI/XbPON3Oj4jehXnfY0tizI/m98PhHZUl3iPhJyWd3cAVpEPRnlD6b/Mw2L+f
awGwKYLKyojj+yKMg2Iav2rQ0bLCgWlxoT0EbZIs/979mZwfRBLbiMvs/KIbX6oD
r9cIQv97bda24Hsdl8q+/bFFHrN9IsSEEA1vIhsBC5RPzTvLqzCt+vOj7EJwm4lG
IXF59JXIOjEc/wVHK6GBi2WO0VqiZDVVIn/jT3k7SahYoEqLffL+Q16fl8Om/ogR
Zm/EG/UJz9P6pDMZ1SVGi9+4pg468g+9hnnHx2rmGYPMt3DAIOTRdOmrnbqK8yp1
39uNy1J9YsvNobUuMoqXrfL4Xm+pl7QRNR9ihxzQwjnPUsgQlFnRbsJbVqDgBCvo
q/K0xltPXKLPcKIKlEG/yTHGuKRynQGld6SD3kmLXVLQszpaWHzKRQTUXM3I2Grx
Tm05dx+P6uLSNABjb3gQAft9zfJ9rasO6S/gWtqfkQ9st6U/9In0ZCQxjYWRhVcH
qcfTEf/RO19mq4ZXfbUVRNXJXB1kvzRVDh8Lxgcy7ijh7lfa/wwA+sKiP1ZXtriW
p4el00VkGIM3sQXySZFnGJoJFxrhV8JtuKcKAFnQNyPMBfDOhZH2tBIzsP1nq9bi
BYMQu7SBwHHWgFMIpVeh1PcW9jqHvGmoi8WuotAbyz8vC2+/I3DKultAbN4Sf5Z4
aRkPiX65Uy1fvxT+zlMIJr7l6sOI1s+C3hUBtJi/bvk7G7HLGZlFkWIi+2n6EL0d
/4otdVfZ7M7eAxZocd+8OVwfG6b/gNHGTQJhdXZJbECb0J5fwCHnk3ziJ5lNbXyM
G3NtazB2qptaNqpsvCuhPOtoRg1ngzet8U9cBVjxxBowUrN82TcQFhabyH+yIaDh
UvAtvS10ojl3ao6DaTqy22H4qIagd+A53hQpc0Cvi/3u61bpjms8cbCpGtQfOOYX
50pnGkshcowKZ942RgvgmHBBePdG725ni5NvOC9VIWFO4ztHyqQ9vsQYk0m9IBrk
fbD1cyI2/87/AN3brXglIWISCcL4VH7CDZ4svJsyGJxdkZqNkOFYVPZ0MY9O/J7Q
O7KddiLzqGqNwbL13ed+l3b3AdV5O4zAuOFpkIkOAas2V6MHdJJnQq3zsxqmsYLF
t85xCW721otI8u6ix48hhHllIPHI92n5zA07CCbzg375q850GVuY5wRyerUd55l3
/LlH+6sh/Guf2rESfFjwaQp9wK3Gbz+5Ceg7W6n44idibQTFELGGavPl2Ve33dJf
ictXW9l+H6sCQIBuhKcoo4NmAIRWGyJ9+5iHO1LYf78BNSDRmCoUbdxC9lZWGFTN
sLBuDXZFjpqlb5W1mcx3YmLtv5UGlExmV4/tHwYKTQNA3Hms0oGwPeNhNFDX/umW
6jGLexOETsKDKE5zR8JtEJzN4G67uLwR1cwcIz9HDb3Hb1EF5Uxjx/D2z+npfC5o
GNgQb3CbvJ2aTUon+l1zADegKbT42T3Wt6IAAMkiu5DW09VSsKxLIG+Gj+/rGymh
35twnwvNu49c6VLPQfV0jkz9Sxx4VzZx7lRkZpXaV1tKMJ4pRUzGx8yobPjaPZ3S
MzcFORCB/y5AcJU2855PBLU3bTfg3rmbUMpd+ZjAD7IG8UDVL8y6I6ooTHQbTFlV
VhAUHZjriiXTd40gkHHf7vH+sjkSA0MMeVmDrb6ypRo0ylkLlfdg5HB7dlaQfGXg
EpIn3cV45MOgrQL5b2KesNpEYQyaq7sfOnfsoVekzEE0ERUWyKWevSuLpJ/MZjg1
eiShYdv7R9EVoonrCrMTO/TWMzF2Be3q6SDLuE7jYb9hJ8y4V79ET5af24FClr53
0xpCTDpTw62mxMC0XtJDna3+zxS7dM0SbvE2iBf8fiYAgGNNTMOgNvEsTuHB5opC
+kZfprPeS4/p+0rjpG2vA+xhiBFbp+slls3qD/t/mT+nRBK/dwXIY2Z0VfAue4zt
I89B20HOeQPGzl3+e5CgZPhMG3ZlRyUg3r+932HBg4Mcp0THBtB0EuhE/OtITVaz
xU+3DhXDb9sO0XYoYdhSlZX+9dzAgeUp6JyInNNfr/i/E9UxVnH/WCwiBhjXECyd
1CQl3CY9xKIkI70Wb7g+4bEBJpWP2eLwqhyC9qDTUp/2TAqvhdgPgr89gYutoRiD
kCLwj2iRkOomo1uG/uGo91Ir9jXaN8MfXl2JWp/SAksCFABAU0Dss2jwHD3P91MZ
eeztfRJ84rYsgt6JD7dKMBfKbx6OPtwhsOxTYBqtRmKbslnw+yiMkXA7DylBqXAd
qb47Hrd+F2rib8COpPUxDJRBjkC98m1kS4C67dSLhX2chBIC5WWFq1WmTy7C7BcV
m/hNZcMymfPnyyiq0dJDPdEILwhANxQ9f1o0whxY39+TttKfZvAHxzu8Pjxa/h5C
Gerkwutf8FvD4X4zSgOX4RelH2QNdAg7MTwdHbgzoZBoB4X0jdZkcK0uuYaNtVrH
o2NyM2c3RWjxdbVsuiULS/y5pyUfMfpBZ/ydIrUJej9wxV41rbkQfNQJoTeIr9Qu
KSk4koIBkiPWG8mq4DCfIb2h65858CmOmYrg5952qlO++khn6MIceWmI/w05qufw
jG/DbDHniLivhuR2IsY+C9qROPVHxQ33jthHGUsUZ1gZNP52WyTPvgOL4/QVqHcO
dqJEFay9VCJChnuFjI23MB5753XO9wHy2UTrhAgWMJwFEUGXKcQolAJ5vLw/18y3
0VcDPDxnZ8/gRvGMm0rbJwB9LxNvyrScRgKulnmO+rrWmAMTstaM1QEGUkviWwW8
L3A9v6Kz/QugofrABr4gg868YPM1e3hnjdryUqgT1w0Lhdf7AsUmKvN+KI7KnjaK
PGXXOfDBi8U2wNS7w9Kpig/Kypt8qyLIVzUqb0m8Ox1ThXDpLxzpSzswepRPifhP
OLUGbiBtf26a7luwbT3GpboidKv1VDeiyvILZVi0hsuSpXOsGzMYg2mk6/5NgiGE
XgI/UX1tkc1OfE0fAeeojOOsbRSigEy+L4AoXsXIlq1ySmk9t0SA6ruN148dfWsp
u9yYXosNPIYSG8c7cZNQBP+ArNtQCrrvNhx7egxWTnhButqgjR7ogrnrqle2Vmt0
xQT17B/VADOW+sGam+X7L0oUC2bHmbjQbL15s2AcjrttTdM6jLOfXzQM9Gt9gFEa
0DJOcWBMEvFsvBQwAWu7yz3FvH6IlRs0Qzi03afxXmHm1yWFZKUVuz4jGhmbBg+P
n+FS5kSzDn3d2CzqINJGpa1KjutiI8OSbvCfZG9yfwe1B9KK9U8gpHovA/GHFhya
WZKuV93WQ+2mDir6BPPov/yNLmwgjzgjBiyMCfrR0CLvKfRhl3SNZ9uDM1PHOCNX
D9Pi/EoW0/oXhGgCbaZId9RnmI0wST20G9W0yOqPBskRHo81RzboKzqJmPvBldx1
da5juIc6B+9a/IgxFcmzyoe8stZ+Y3/6kLnR8Qn2PpJHtKHtEnEIgto5IvBOYOR9
9mLGoPJRaz6awSQUdNlUg8kNwFqi2ZU+yKUtUoY9wY1G9agrByOdAiAwukw1VZYT
xOQkGXNyc8ArzN7CcuZ6JqyGTrqDMtwW4BMgmAr9rIFsMictNmPnIAF8tMKa3bfK
d1ZUrSAgD8HskzWCV3Fc7+EoNsuhNXmElK/LNxjIy/OyCSRkgF+otZd7s4Qyg1/a
159kVZHxgo5OnC1+jcxagY6vhRBbG1rKXIJWBHczQCgXSzL1pHDiLsR3jgNnjI0d
yv8ORUap8tGezpIuQxkbA3OTgP2dzOayBqn62V9KEgZvO2cwKY+S9g1iI8K1dCGs
2VOMV/y+ZpARcXTzO2tVT7hgURMaMcdSh8ViObdyrA9+hAslbJW2n2fbLVanQDyb
W8EuDHgs4lsiihW3fBP7yyOhU5L8rOLiQPF5jg8oHsuleG3FIfRcGgAFhJn4Ht/c
PtVRLw1CBYwUjqLWd5inH5lqU3N0UwV9YQJ6IWxGWWRT6nlNh5TpUcnxn7m9NN79
9GZCAzaLQAdirU4VvBaSTeDLEFttpxfBXbRDdGbuUYVzQsDLdFrZlQEheGi7oMAD
HXw+t2LieQLgmSNjNmuh46+IDl8/XUGQwcUK8a2i4eiWlvRUum53we72I3rqoGPV
vNHxUcecxrXadvuBo7rMOgvpsgpWI4qR9/tOdlxAomXqToqD8Jc7zjgEJA7tN841
g2DLjlf/FRzXLj1AbtzgCtLtMl2SQNRxwXSi81CXGBee5vM2dpsXEojjjI5rYm7F
beD+Gs9lCcc+PnDa0+G6yJDq3b1RXmkMJqQemtHRDS2oL9xAuZVVnBamN5nq81pU
KLNfjahNNXPJeLJrYvu7ypOu6jt2w2ZtSKk7tzGTWNkVcPzU8LTzo+2RAjNOzbs8
w7WDEdzOdoLvTb3k+YtuiA2gYVAKL3r3D2v04v4kOo/h8dysEHN+fQLihNNeb4lX
buaqWlmPgUyDQ24SLSr6ajvaXseeOlnjTIUu9k17va9XlTEL89hI8BJa9BWGgA04
EGtfwvl3xo+XbBmtrf1fWdiGxRRyoFABUttKY4tYJOjxWYfRydsVpKx3fPpmM5fA
JHss1R/AZKFWjCaFPqpoHZP5O43OA+90yL0f/BXIyti186igIDxERX9Yt7IZY6ot
3F8SV3/ITBYSApzwqCC3kk6kCg7BqS+vceDeoUNkrxwBP/4+ecbZlYEm79bDEon2
EXNQlt0BA2YV2yPVtoi6OCT5xK1k7WZRMYZ7IK8ke8P5G/owdu3o2it/UPW/Ikju
7NpSFVAvUqAU3mG4C336YwQMKPj1Vy+600drX3G5Hg0AzkDerXuJabqK78tUH/4n
IgIRD4ce0NBBKVXRNqjN92KAIDJyIz/2brfkLTIab1TA5RTeZ6I/KNtsz/d25MZt
/LXvPepBMHkgukh/yMDrjw6gcElL9YrzMBarfsafUnQzstv/rYGDA3lvbRg9HvZX
0TQxpCb4Y0+vXKDVYL1bRZNzkVvLKytQXsN8U79QoogtqojeBUzIUtSiQl/nE8Ja
ZgZ0PZXF+DBsCamIwnDcsPbViE+iCIUWDFXCMubprE5v9Vke0YhQ77JHQiTRqs4G
KpJpTVJq2Y//krXFiax87xwZEI0beDiczHQdw480X28et7XEcDPx/WnELq8DCxTO
8q0A8lLBhguGjKH/cQgmFd4AUY4UkrZp4bj5ke7qfoNcy3oWBzg7I2cvtMKLvJN0
HfLqLWnLzVeaTpqPuWXmUlZRvvnXyHhf5WYAcIvSlxQk/SR6Ek+vMlqQueQvDfC6
4LSfWPfY1wweTN/93QoypPehxHG80kr6qipXVJ44Vvf3Eoz4IsshsJPyVkmjHGC9
5Rnpiyt2WO65VvPKSxmOp4hj9g7nnvrDeFBFQ5f2cpQjU4vFiLcHkb3AVrcFAdDj
W6JNGSif/uWHk12ErVgEkM/qiSVPZScvLy+i3qreiM8jxsSVjTqtAxPVuB7Tfviu
0MC2nzbOvdz1S3YIQpgbaAnnBsk5SGmzmbBMAle0p27pVCRQRLfx4UNaZv8KRjvp
ECGp6Iqnk45crgWPdgmEjMJm+ssmEYZRec3p9VaJHrd3F4s9tvudsRv1kfedBXia
/L/QVB/KAYuvcjN6ACdg0wTnDg+KGTLGBTfuvZyOSxPcYK4F4BjI7ZxEVWb9RgQB
dYf2DCId08kRjr9cyFn33JE5OgHUInHetg7OU5oEQlAk5ia2sx9b01KPe+fgwQM5
7MYvlOcP7Hxt4MlbqqJ1TZjmKmNWBNL/sH963Ks5kzM3JcXd+Qk8ysOye8zX0Cm5
E8cf3YvLY3GP4OvIQkc3DzjDNaXmSk5qmTA7bVu+Lhk44QggjuPmMG+UcVPM2hnK
4vy16fAHjY1AORKC8oQraxMkRe9EddcigJQbFiXi2heP3eicE/tbpBxtrqKz/I8V
AHkmoexo0Jl5nKoLzLShf3tdD1u21AcHB1c9fxg2Hn4Ys+jnOPKyZU2BuqqK4WaF
MuKD/UxbPqBXhuFHCL0nT0kKtCZgweLWiRv6flVOo1vpUEDTvzGLc5u6vdSy0Hu2
H4Vukdx9LjsvRFBP+z3r06UJ6wD7hUC9lRRG3HwBHqvOhXJLAaj2sHfeN1/eWiR5
vPIVdOg3I77HTpXAPeGboftxWTgLDMw/SOoS93obKOT8xJ3qvLdxsXlsxLqy4sHT
nFo65DeA1b2+hUrDKPutNA3IzdlqNfgilQT6qTR6fvn7GelG60jydU7nLXFA5lP/
QSKAG0GW/IxxnTAkalFkCE8rlZU8quWiqDGnWAMJVJ0r1thG9J5tM8IMrXi+XVU2
CYgcv91eb5H/yZfVJ5Z1vNpXslttY3s9BkyHeonhjKbEUY9KVnBXpj2fLvmzzud1
a1L3+sBA/4VqoBD7oi/1/v9pxbvPyZyiO7ctLyRNl0pEpx5i8aOYIlzXiDEqq9hk
XdOvGgqO9fK+x98p2X+tRSbXtSLEDTyns+99EcZIdQF1pxYCvwi/bW7aWJZDhkki
UUZrIuRzDeqHYeDOmabKvu88WJbk2rS4WWEcdtnMplQP71wgV+7SaZJUShJTPc21
a7t6rCVo2vyTRs0bkLTRJDSH/nGc+UNWRRsopKpMv9E1wKVC3Ze76DFbA2UgVOxJ
gWcRm00IugtY5yRZ6G8RIUQ5jgPcFuzaa0YYrTTWgFaaF6jZhOYjXrrnFufIeD1U
MXk2QPKGdsfUXhF/BdqgF00Y1gmwSFHaN5cBI9gny9UJUb0Pmg3awD/xVUxd7H1w
3h5Q+gz7J1hkvkx1sqSAZ/Xp0r6qiCSmerXA7lG5UoCprXoNUE83TbGCnQdmeX9b
gTxnB3Zz66MU7GAeuKxARWFa2szP+EY2xryGvrWSX0eqxjlJZfEYl2SJzFj+/yB8
1PnPKxsGzUvw3JdteZCIvrqThgmNnqMBRt7PXyYpYDxuJCYFYO4P+JKZ/+FY9dBQ
4nC2GLE91TwObQQMSZPnDTfuByyKtKR0X70PjcMHzbxnDo8Sm+/PAxllk9Yxp5ai
yS8Tbi3j4dXWu6YwZJ+jWQ+ZXaywz3iaDpoftYWK5SbT8ta6zaC9qwA4fs4qsyf1
pgS30nuR028ZoF28EDZFSIJSR8/ohv16aJFhnkaYfKby39fEn73ehadpouBOtLmm
+GrLRYzF3p+mxoS8aTz3J64jMJrJZ4qV/LSKmZGwzfFlN6GIriw6hFxrMwmTg1sv
yRv5T1mLMALj/ma91voDmZHaePlAvCR+dRrEGBhgTqyWgRxObyvEm3SCoofvGeZz
U32n1+vbRl8JH7w+SSywYqoFyQz+bBx/Zymx/OXjZcRo6rODMqxYNlfaouA/Im33
XdeLLdOA9z5KwaoKQWantZ2KcyoUYD5n2+ego9yXjtekY+jDfsm8bWDORuTBHUvQ
WmKOqb5yu4TIad0IGzYTMn2EyfKTmO7jg8uphWOD4t7OzGAufQT7H8pXiMk2sVTb
EZLUNJlUmykobb+UkZubbrGphzZYjS7b+xrWqy2EkKaERaTF5jMfxKyG4r0c2+dd
fs9ghpXrY+AApR5Hb0wTzZ7i+BTQ3ymkIIDaFy9Dh8gcOD1HKlXeJTOwPTNs8Ilr
3aV+Ff2AbMMMo3YXyIAFti15Iq9hFJdEJ9zqrvyaI2Qg/o2QiBi7oq6jKWo2GPtS
8CT0qkCe6Cr7zNvJ3ywql6cnZoKZRDpNsJOiUI5I5sitZl8WVrYuid3RUOP3hKcc
EzolrkkBTY0OM2E9OeMygKyllbY9ru24qsx5oErwbR1DW7pfNDceSmbJ1HpmhQOZ
3cIcTVVNpfXoYJUCEJLltEJ4/qHLUWB+aoodpAYmAL5RSg8uXvUbXEiuhLHCvdif
zA+g/oywSlh8HFP6QvHQY70gZUZ/bT4qcNWVR1RJ0/puOADmLXqxKmRUKaZJfNwx
SMsqaJriHzGKCCZEg0Jwm551aceC1jFwj5LKj6qEgULVZBu05u7vINOV1jk/fIuk
5NDEF1WbSnqHUi/Kq2TSpqwksg1Vy5+eWDbSSTpY0RWHViZ3jC3Dpz2z5LtxbCcB
SnvorDU779cqmlgQO4MM0iPyzrr5qCUuGFvE4SMgbvau3XUHk2P75iL+v7VNwYHJ
T2UdZ5CAdd2b9de24kIN+v3REPoSxeh2S+EU/D6F7ByQ3xNSuYE0VBaYQUhbmvKg
0v6Cuns4aAcgutY9qQHz+jeP1sVhaPwH6VNOvojMp35J/L4dd8qwnpH5oldMDyGR
8rbaCcWoziIY0tiIItgDC7SU9pNAGBqyiiSQl4aZDEmVr8ZIGHOEvDrWA7KqImRG
XJ9mfa51+3wbCjcjkaQxVlZbnzQzF/b4BpPam/EKJBHCx+CVFrBVXHzJsRRUm+Rn
nVhrkFladm0Za2mWOfzTUL9DRnk7UoSuXRiFdv5deGoVyFWde/wlu9+90YQAUbHU
+nrpsdDNOtm1uC8zzWGzgprNBNOfrhSPsTp2bhLjPUzbfGZ+5TUswPtlKQvrc/NO
twHNsJU4dUpyfpRmdg3ePulupWQii/u/kI7Syiiy5mkyuLgmcYiswovriWMi1ofT
I1Kkx1J7B3xCouD0k5s4VxsAn2PNdMywpZ8eb2lt2QDe9S/cP9ctkAT+Dw6bJuT2
kOnRo0dNyh2Fno+ZFRsL5Eo3wpBcpAG1YDySaj0jB43mxwEVG2VnE+wdRjMKHFa/
2eoWOcNuI5Gt2QeryuSP+luRmfzTS2CYM40fqMQ3tpOnDH282EB2oYUxZXdGSNUA
/jKyx9Qayl+P3Al9rMbGPnpHnB7gjEIIiVSngNntNMlucZ1iw+LkDy7zp4qG+0Oa
z9cNmk0BIlk+uGFuou2DQO2tL5DU/eB+6bMX3bms2MllMxdN83KRUXpU1V1y/cIo
/iL1y32MOuq0DX4a6nw2xH7T+3GrW7q68ROxocGwZo1ZBN9tPfqKSQRGnqdO0HzC
U+T0DyeaBIDszTjR8ToYdi6xV8cpKfLS4zu7UIx5iLbjfwZNzB8XvEuBcY1HHN4K
DP8+q49OnDKS240VF0TwucACrnc/NuWzyboMju08/THzvU894ELWqZh6K+MW4ddl
d7RVOZO2er91cTefCxYJrX1yIpxZmz1p4jORzdSD1d3pPG/JB7pFE+uJDL0DW1Mm
T45TDq8zDLvLLXsmRaYLOBjUh5Mpec30Fa1U9IaHdyl9cfzxr7zbcO49Bfpe74Zr
mh6yXFd38mCVWkeFK81mKBkmXCJj/DfAYUQTdQo+fOnAnH3L+Mv7IuSqQZ0m7bKV
g1FazPgo1KpbL8GI+W+yPrD4X4feBb0k61QzrpbpaXs9Ox3ESqWZr2vfc0gX9dnW
bLZL/sOGUDnAFfO5eYDfLJn0zTJwTy+YC4eHkdeb/ZzIo5dSq4Oo9y8HPBAY0jfx
hZweF5rXANBJDAWogClwTkcWBBobCHWk0ToGu72bCwXTCZbx/0orDq0TMl7P+UQp
yfmusTOxbVRtBYj7ufp2BESPUuIwak9Umkvo3s4jz55dc5C7wo5+0w9Oqb45lzvB
5StE+fkSRGYU/xAWgqfiW03cvsuQmbITMPZ7aK5ajgtQRwzEO9aj9SSGIqm7VsCe
lG/ojJdKKgg0HZW7ZuebWHXe6k4RIAYImN+lHYVlsbYI6kdrnOCTZZ4aQ7Jd4rf8
/uNUVIN8wNZBPK3h5089PJ6daXEPOuLitFNv1tOc9zBEKHEQMVFmONXugUfKsBPT
Rf1Se23lKckv+d5921HaURYxLsdS9El4W8dNiahl4YXRBUTKtCmSgSGJPaalxXbZ
dPFN3KS6lY1iHs1AkRReHR59WIK5+K0JqMJBMTIIuh2MGLduatoUQAKMaQma5dKH
yPoRKgjaT+u0/QQv1IWuDNdyUGvpuOoDtUhwYWPA1qz5VrllFFD1YYjZRSd1imOd
xB9PWDxKKpbZWNYfaqhe3ujtKU5igUbNxFswzk1wpH1UIhSrsUOnxO6Ld4AhDY+B
PPWgGbQw7QrhBJKbqoSpze7BFEqAZ+dbYcVCF4i/qVQmTtX7PSc6tDqkQUCRj0kY
Rszp9e9RfsSv7orqq4cgkh1GdaO++f6Ipyo/MXTDb6tMWl3n8uDbfV28wNZSWDd4
Ss/U9BuqUwPobveJjeekHAkXlHadYlaPUS5Tje6+WO9k9xAq0s9aeo5+MGG1C7/8
eAJ+7Qlgy4zIiGOML914vIWxQ95rZ0mQClftBpnXGiKbBJAxyt4dSL6ZNqFK5qar
lJYWGq5jadffPplFatRgy3i+pfZb4yDtECV53iu4sCNllVqSzYrZPEwGsBJ5+TC0
j6PryOpXm0ZccZ1Ge6EU1fTJAnn1UwiKwxvSjdcBijATi8UQCtquBFoPSh6Ih3BF
+eH+Gv7v1Mkw/vSw/51b1qVkPQjpi+kV/iJcRdJiwK67VdnA01KWRqE9XnZpFffA
XtrzQsU8Z6CauRPq6yr4fxS5arMMxHg7u6ukcDNHe8A02CJqBI81uhgaqWzILD0b
mQ6ZTr1EadSDEhWRmErRraT3e1JWkO4qZx/8AOW82c2g7iTbXtuQCtvtguubiSZ8
6HECDwYTaUUDLQuVdmLobtG1EYRkjaJGvP7kA24JeI50hlabN/KKWWpbkszOcmQA
GyA4FBdaFbh1uYpJq2IXbZYFjEUWCeV5oCxPty8ubhwpAQSdIvsNt5OI7jyVoYVx
StNCoQppIec8qHwXrGvOgnVHJWGK1k53W0gesSg4hYMxYEzl+RrOD27zA/IFj0pi
6/sqcaCZCY/X5gawAvAgLQq43Y+CBr0c1NKIZFi4T4tL0rlLSuncoAG4JJNlTb1D
jXDYiIlLQ2Sz6BwiWcB8KPStbCJ7BJYemcg4EtM85wtWLXADHaXdhgMGhAzIkvHp
k+zNXvNl9PDlGy6XcavgURZSORonmGdoe1CYCZnyNy/3BNuMbc0Ep4RbJyBFkbDQ
5KYYRKVW76G29XBqB8q5nBDyL9BpNNdU5DMcF09nBPSsvlyM4EDfDNhWQnrxSqUy
NU0vkseg216wj/Bekc3j9klyocOPmdxG9bPmWszY286lJAJF0k4yjJPcjdsO9XFA
/4j58WEMQO/oKLmLTjFVX0e8oImxdOiDCq5Jy9zQjjV1bgYCfd8Ew2vzfgOxa85G
thD6I6cqS3RF51+tm01a/lgDJtyCj0I50FjfPaG1EJ3lrYyjv5OVPNp8zYPyxLd+
fXmQ6yfnOgP0gjsOZrfGR5d3ZP7DtcpHoFrn4ILZdgXgqDR46Vepnf4k2Vl+aKMz
mdbqSv6bip7NmiSOHTp1GT7yWqRzHSmhJgR+J+4ff0OtjDTM+qemT6DBK1n0RBH5
nWvkUES/WOI+5kwGzAAQbShWBe7+qs95cnI7b1676JodT2y5oEAMRrzWssdbO9O+
HYhAVdJbPgT8kJ6PfZoAdfGN5AnSWaEMc6REG6TniDNaJjYv41r/T/5K8beyvABD
Xhz1zudL5SS2Cjprflao0UPL6DzcCWHGYOc99PiAEAcI7FAdiLpwIrCGq0rghNMk
EwKbWpyN/V5panMgh7YwnAbpHgJsmGWjIati+AXMUT8BWgavYIMBQBKsZ58ZdrBm
2DKVgS+Bplu5R/5UkSBGo8i3QhRwtwTSIRpJZsrYne1UWfCDX7+9/nE2qU/51RSS
ajfGJVNYq01uLDlT9o7iTd7uOzAFwY4GFNf9DYyRFt6sq0qm//KOnprN0Wqq5syp
vP/50RJPYxrbs6C4mwr4GxxwbszBfygh0BC/j4sE8l89WBvZiHK3D5ZO7y0OsP4I
QcMePmgq3goh5QIubAUO5aJMDF7VKjW1EyW06761cx8nPUT1ObHpwRNeHD6HYBXX
RxIUfWDdAzTvoFV9QPaReuWkN8j00GD1DT1Tykghyx9TqTMtFZX8uQpQSZ/e1pFp
smo5WyRENWM4vi8pP8Hen8Urbps1dH0zy0QjwQioD9iDuNNt4Q5H5D8TEdgecN7r
GVlh/+oC8TLEmRCaxrhyf9YRP0UuHiETBt2a/FxJhJUjndxb4p8nNiikM3EpJCXM
RrNhDefYB1sOKpFcBjTLW+sIsGG5ijeAjt6zeOM0pXQtt84kWj2qY+gJrG/9+Kwd
iUOivxuYbIm24PrmjD4d91UXDMptxAMDcTw5xIOvsmjwlrFcN8nW16XkputRmcpH
BoXNK1YvzLHrSitEIlM2Ci8aD6d++/JbHGNvlV8/nl9FCuMOkAvXJ34BtIe1+kNc
De/34rCGM0QbcbaclV69dd6sGw4KetJWOq8+Ur/KclDseftuVo5+dgNSs/bcR2Wn
rVcblVAzavGomp2Il/yPP6B7an82XJwHB9FJnIsF2bnXsDzOPDpdu8X8slKUZkCX
ZeMyEVqf1q5Zg/m7INjh08g5GBNcG7GvFebI0edOfhEF52zRsneMQHWppXl16kWj
W1hHfpoxkljqhK6SJqo1ZwA+AG7kkSsfQAQrTwdbGvemQdvECP1YtheG5zCyxNnu
SvnTgIutDXEDyABV9mUxQUG298oO1ibVb45/742rewWfwUi2srS94UycQN/JPwdf
wG2O4GR7K3hEE3RvJtie0TUBkjw5QToHeACahEKz00MK5E0KJkcPRypos3KnABpB
ka3/OaZtSRiXs2Xb4dph2DHWa8HJyJhe92OGqI6ybaqJY4Swak9pkQ/rZ1y/gQn+
lnNhMpfB71cBua9DuLaXgYG/+xSkH+KXC17nvOjKbx6g6dm7/nLYF3+TnRNWd2qK
biC8419hGqrgil4K7Ua7ecXhohJORSO4SdRAUGF5YwgdgNOgLzLR1B63UiVTOlHP
znmKDWIoSl249lQXnyRjm4QSNzUL+IhHHz3RuC1F2E2P3DRaGdt/PLndlyXQGI5M
t+6zlMpcbBf6CELk5St8fUDYtVHMpI8P98UCx9c0xAg5xGGAxcXIFDZNf0+pGQsy
zFWgCh9BC6+LSomK4G+NHFrWw7OxwACCeVGb37jTpsdma13WMeVhzEU/NgLGQCL9
si5qLEXJD4/7MumZUiQt6v7Jk0F1VBWLQutVYlyrKl1kDsUcManXMMORnulM0A9z
tnfjNaS8B+/SwkJ23Mg0BNX7dcLfF66q9sjYUwAFLaLRY4aZcBXkId2TlKvuXCt6
jwD3hGkhHrDMsffkJIUzU26l6R1K7bXbqfMAO9/E0tHCSgMQEVeaDUIlg86v6gam
nRWkqBjWMp8ZOzpfIWs3wB2nkKpWCx3jB7WfsBAM73KMy5/6XZjHQDFE2unGpRwk
7pYv3LE/utQyl6NTlTprLsVt5RWGonGbrX+GtaE54ZzVm6tzCXcpnFEmelulqXuL
P921C1xH7VqQfAviZiGV9tGty0BeYHjZaNNi6XaaOXhdkcVmm0FCribvsVqpRpWJ
YJEauxkeTkuegsl6HHpFQwNPka835EvZG6b1zV5ahY/S7WfYYt7N6lDwbia+/DH6
XcxvR5m1ovPjUjUT2Hvu8Xk3vdlq00WIwAhp1424WX9rQS0JcqOPqvBsLgGqQMUX
1ZqFuvSIzeT83HfEnRMLcdzOcgixosPwUl/K1X0HWLOC6wkdgsh+59QzdOC/zBHv
TuNEpg1wmrJ0tKoACJ+7RiZBxm7xQ2D43NLEYNsNR217/5pvn5HTNDTKXZm1mApI
DrobteiKnDCbl8ZFTM4/W1RKN55QME55g7VS/B8NDZKtKDllGJVPBnheqvpGjiyQ
5uiUfiWwskjb3U58P5R0Ox4eBllJWWGX5OGu97iSnoEBBh7DPmshRBhz0UEimNLZ
/LtyNoyEbVGomIRN8XoGaMMyira7mubQG9x45RrYd8IdsxgOOm901YAQ3vfcChPK
hAH4ufOaZelSkUPtoi1mwFEylon5o3KorylOoesNmRRpC/VD2MgJ5mnXKS0E3MPq
PXoTvs5bk9YXr1HZzhEkbJoOEwmy6SdSVuOFlaMlcbdPgHGpq4ja6d4MdRW7ndjz
+vr/PE6MOaG8BRJMsgZ03qNJIkWH6I605j2hN737ZPcFeAUKTrgEZjbDuy43Q53U
HJfBagsb2ZuBaoF3JHxZvuvfDRS9DbJHBrd0voWLEcOg+LQO2yQZtUiWYn56yZda
ARoEHTyWY4J88nU6IswYaxhZ6GGSxvANIhTrn2rZNQ4JTvGcyG7hahiCwTczSiTQ
GZTJUb0uw/aEo9EIdTTrlM7dUXJCNeSzTbjFGzdZwvE6ClTaPlH73f19+Z+hF5k5
y8pveSZ8+GKqWrOM1RDdsIY9aHZH2FkPgBgFqX8ZScPLRZ/E7tLhQ1uoKrkMEeqZ
iQxuRvFL9SzBQR+vVk9fvCnyexEqi4jMlCRhx+fstHFaaRzYJSvXrxsIMmTdd4bp
IIXQRFnrQ/S62jLEfEqgduXsnlYEptX3ybSMrlJQhZHp/8J+Y8yi/AxvZXdH5WM1
UoOT2QYMmtOVCXPiy01Q3BMsIsES9PavcAtH3bis0CgzlWmxBIYVBHqhxQhUqN24
UfW/rEErGwq6m6h/Joi6UvKr7rdR8wfImqNZvNKAn06rf/jpXWKfPKKZd79ri+9H
k7prv+k4FjbbuS4XcSaoX2rEx5AEBW1Wc9Kco+k7dInZ32O4iXZVQ8uSAjgEochP
809mnonEg+lKWfzQL2XVISAXa4crqki+KP8CKdV6443lYneMWqU05LpKqySmnqBj
E+/O+S1UHLbRgC03voOje0cXg+NASNHdtSKymlP0QPSk0JDIolSBaDQT4lN1JYO8
CiMkEulFsow2nTT9V/l94XWx9UYFH0F+vrh6gIj2UeqkEnxQXj+OlsG1Y4Uxuy8N
B7HNH8PrMYrkl9NeMyvzYPurznU/sp4sxVX5C0I4nQEvA59eV4sEEozGzjbnXN7V
8hQfHXnJYjB74hiQP+kCr7zfzJsMrmzLYlrfQSTCV4FDAuEwCkRSeo4cEMnIwZM1
MI1LmUUaM41ZoGhnsd6UsAJiWTd7LjIursftHsQ4nnFaEotOgf0os2XzvJy3voDq
me5zewi58rz981Sa8vsCif5dua6QUjwo/zZlhfQoXDgqF0piBhU/9S5rriUh/bTl
bHq35+Q1X5BENP4albfwGbNLQdwwddxvXy0QBxyqXmQCWmkKGYtxrnxxr/klfOld
WbfduCGB4XFQN6BhMGZ9/fFJb3eF77WoDMB/NV6Pvdury5ULilX9rOstPFXbjsez
yaGA2GoLz/IIqDEZOWKogpJzy3PADCk+c8OlIt17QizxBFkYq+fNYLdlzBmofZ7Q
aHuMTyB+3iJqrErMYMdt+DohkMufkPaUiHRr6x2A3hNv+LKP4Qwj7oPekzjdIKGv
GV5oDEB0K9dqYOgxBd/Gn+C/BP+QucfyJFR0LYlHqZr9UOTs2KCENeP1BEeu8IEg
nGITnEmpXtaF/wwF0x3Mq9yoTO901D6zWXJfX4JPHxRMzENEP816WUJsFIpkcQ/q
dI6n2VmV6HBkDhDerwPXrrGNsNnOpGNiM79N2MwRe45eGt+W2wPwyT/+4/9lGbfz
fXVbTGV80SrQTmzntK5HlsG8QaXDPTXjLY0rbQ57bbs1TysnEs+O3+T85V23Napo
GmdWr2cOSAu9hrRIJ7yFTipfC4TR7YGiu9LoGKWG5QeQfkFXpKthHfUt751stxMY
9d1MpK3iNe3+GThb3uEnCeaXKQ8/E+lXx28CWcTYICnXZhXjeBudO7AWJ9D3XMjy
jgLizZPmksQ9kpA/RED+IIFbsWe4HRuCKGWykm2Jeutp2SQ4FosM9Se/ji+L3YxH
O+0VCPIsc4RxQzXNl4GVk5ZBT/uPLSQoqMTpNkHnWawA+L/ciiLtNcMatT0rwWVS
+B/9KGck2UyKG7GPfyJuv+q/DrmU9EZ2GnKmkNo9U2a/IP2qxi4z7zM0tMp2VMYM
087DC/3pihZZldh8gZ5v+iOWGQo0QS3/pAa9/2U2ZBtSPHYk32YvynpsOA7ZsrrY
aHUSaLb69YAc7fVjYL+HPYkwwahBKdUUvOl3uSkkMwUPi3yaDm4MtFvz47iok216
DZKIXUrCyhE+fmy9ttFJUEJ/aZneM5yn5vGx1HRkA6FBtsNT3Tam0KZV85LEpKUu
cLSBNHAdznnUIYpfvq9dtHnNPNljZSQWVO8E/13x90/PGl4hPnEa52fQ4cLqKUcX
X46ns3lFhOLbclXxSGADWvMOWdy7Xb4ep6vGk6TLcmtJTrnP/HJtNhUvI46/5sEH
Yq3piIq9BaQpqM/0UVhUnUddmFCwN6e9VFQhXCeDcXVbX++QgwWUAGYMtniBnPjY
7JKhsDHqkRHmlasZE3xVwsFdfRjWhuQ+QKh9MD94L/VqlFSe3DSqNfuGpYD9jpzl
Wkdra6l52oTPKU4bFuiudCVCNiVOqAhcwpgAf/jA9UtYoR972gm221Q9G2EMnNd0
HZfSycF1nBTY9gp+7OkgO9D6D83A0oiGwW6xUF5gmjapjeXfl1X/s2bv1QuFy2QU
z6qgDPhNIFqMWYo+RuUyExqugtMKf3uD9O8vjUepAuXxF+XVUNzbkqSTWLdrioBS
LLKjZUnF71P11+e+Yq+ieeht45CAX+IxEXdVXUjElrZ41IcpPpHMt3TVI8ag4ecK
s9lOE30e6ytj1TZiyPCAgnQj8DJVlx1674dWBK5hj1bgxxnLJjhyTD2tMEZA2Xbl
93rONSonbXhQqeCnMtSw1fyKO0OR9p4uUB2E/IwkjJLdDYv51RCv/xyC3NB6wzNC
fTqb9CbRvG0RP+cu/I0iJqheSGVoxbWmkY4zBVTPIYQAdVw3NP6l4ETV8iB8y8/P
PRGpGMJW1CQHZVZR4SBeD0enD8c4h858G01eKM3kUKrd4gJ4wgezAaCy2VHM0Fcq
Klo0Gf+/kdG/Y7jn69+wJBRWlEmBvz1sutmjqijueLq/xveMyrH3MtrZgeK5XgBC
a9GnhL76nQHo2JCbyt5zpOkUQRByaZgW2j4Kh5XbGsA/bNJ+57/yAuQEla9A5ug6
68xiBPGB214gotlD92zT3h9NGLHwYiu5zwB93dwY2Gnqnulo1CdtW2rPidC0HO3B
Vi+yDjVByhjhbbrSvSSkXhZCROhFGvMomZ80sxpheZINIQeseuAUswVtRomezkrc
XVG0OU1POoM8livs7mJLJLx3CcLbQZL6CiIuM9ZR6PS2qEDVMMO7t7HiZF0T29Ii
vhphaT30AHrkgCAaoGzKH1i4a0RGnQj4KigkiDQRf8CC7/AedhbwhX47/Aihd7gn
QN+2xzHLvOSTTwYy4qG+KxDrvhvod1W9Ft6wsZsdUNM00BKvKlXnf2RiXrkVE86s
j1YHZvg2TeGDmRfKoEu/qShCmlvyOXxuTtkxEGdd4TviosHebFLZzuLiDS6+NWUn
tfrOeAeX7RXyp0wAFrcIOkrf2mY4ViUYHJ75KLvD/kuhA1DjtEV1rKO8UtjVqMqs
B00KLeJgwKm71Ct/0Iy5y/ldnAf/SZRbdzNLNseBFHbQ2yrvrVCKDgc7oFCbsn2z
GRfjyxwMzAYRkBcoRh9yaeC9RvbaziMaRy0TJab+8K8A0AyNLdaN9+xiOS4OLPve
KOkJsX/6N+9WNa896Sk+RAqvb6wMpwHHkfCOM9H2qxg3ZhiiqfLfVHQTCZBs6xEh
27cpr8+4o3LUfHGksEy3aJ9doRAn/SvEP6IsonDwvGMaaa3Pm3eiOITKvg9JF039
ul3ASp6ax0zodSEH7ExE3zBMDnr3e89oTKL62D7h3IUGNIwWroazuRf4k6AQ+urE
7Iw8nbLrRmI5otyGayIaXjBUfnXzF2mbiRtLFWljxHDYr+FZFRE3w4rUcM0sslOW
Ie2FI9b4wvNWN+auVF47nTo8yEOS65DLBOsKG4bdbkPad0AjnbIkmc2Iis3Gh8IL
9tq2EPltuTVSG54EgxSyoeKzcfT66NlJ3cr7MixKhvtgqXuDU6r6E/0OaVqYBDZd
IUASUgCTL826TcJcMOuwBzyxzjh03GifWaO/U1+xA6q/a99X/OnZSv7k3zUOe7UI
dnkhZZsmpR3bJI8IzJZZhYvaE3vkJMA7qKnOUVAog2ujVverqjPWpUUzV828o3CI
BQ2PB2qyOU1T/AIy2TDBeFFPgRPkXjje6XWRIiCYjgX4NFwpbtEHYZg9YOD2B0RL
5Jv0bRq4iWdcXpwRTX7BJhXD79TVsnVLlbs4+emUHG5RPkcCbTuC8IHlOUGo02cU
xh+o/V1tHKXxutg1X8ytDim7nOc39Hk8kKVILfehuYiclAaUS0Wm/z9rs86aZw21
6205kxdJ8jvK/2h6GSIevECJzME+Sfk8y3KeHGPRmYMCk+YZxHeBRQjBZgz4C4aH
eFDxgRHDY0HvdA+kU7tpp5ZNnCL4LrjWUteSHYkxVXVrPI3pTwFYatFabxgy5Kdg
YvP9nXsVKMfbZb145+JNlI+hp4SlhdgUvWW5UZpiBzTuW0tNtxtGZUKnjaOmdDTm
KvleY8Mw1tbnbjOaRR6Vuu07arPqoxFc0ajkmv9cmG5jo7+yE6lFBkRyUI6r/ILK
k9j2hRnBZ47E2LQT7UmNoDk3AWXCz78vZSiEpkk66rDX1FaCF0qTM+pB+bkGSw+7
AJ2u0TxyciKbmSwUObnLDVIY14zgYSyoNWmS/UJmM2vEPTorkjQMmRqdX2maLjDo
+Ci1bhAea99r0lmb5myl+9CcAKqHDsa9rO1vx55wf8dLOpPWK7ETVj56YVrNGofw
4YJP9HVjKN22nWBDA++jRAkPxVPBgbFSdU2/u89Fg4z3ToW0KWxBJOavNOJ025kM
Db1L7py76VW7r8eNLexnCx6VG5VkqZ7av4HglyviUAltX1so/Qjwt07zDcpy1odQ
H9KAnURHNZhRufPhqKYKItcsF4AfLZbCEua7fvejEarhqa8nRrf2kkv+kUm2Tqo8
FMkS6l7GyEI9kG4nmdNQD67lHCCIoVIfBxOh4nY01GxmcrPMC0aCLpFesBA7wlYw
bRPmb7+ObhvKoNl9oFXnnPpqOJ+ZunkzR+H3mU0uNXbxF0BS021UoXlRETwYK0BN
W+MoaarktkVMro7kQtVPTJJm/nlfsc7kNH/D2Qz0jP6jgsJWaS7AFxdAXHMREAzv
5N58QlQkOlHfqRbdt3C79BXkkmAEnT9hqcZFPbTfSGxuFKGwetVc1jTCdGSkxbkI
KHprevBlTshj0/dyY844ZXtaUCpF9XI2bwSxe4DKjL9rGO+CMG5ZIRCj7UF//vnu
GNJ6JanP2NxLoBY60Q3T8S288v0HKfOghFCuPMJeGH+Szb+CaN3SH7lTTeCguJG5
z8OLFM0Zuip1a0h4W1YGZNlU6A8GWwsuBtz3ywEtrOWkm2WRiDOGaGjsT9mUwrpD
9gjtnMqitD46PFRQgl7yXjvXXf/i4rXqyAFPR8TN4xH4wSXxGf30AYHAAFnXXL2U
dfBSDGQC5HXZu/7BwZILYWs+5J1nkzax0KGZ4FcQrACJbNhWkKahMcwYPdVtjVxs
cMX7FtrBHmHyhwp8mJlwACN+5/4eIlsB9pFjLKSJBLINCERmnzapt92VaIPIeR05
ZH85F3DXP3IO7dkoc34r4L32RUoPYXTpS4IQVlIxgNToGF6Us/lHdkPJEWWwxcOT
fEfr/+LBaEll0DtjA82/7yiskCsrwPkuIIjewGKOO5HESDET0B1O+6FTGQ0Kxg5+
37yTRMlNAAACqXtgINBVG6xrtmvNEBLLEunmPQkff6L6tHIvtQlPmqcKFSAs+iWw
Px5JsUuOUsToTXp5nf8S4d75QQSz+Fcq0wUbHY5JAOIdvoK+YUKqQsVU3eyUJi8M
jBHSU9HKMbf2sUoWqLbi5Yc6glHxhxVfPBKHW6ur07JW9D8QaXDzpVsSkMl/Tl3l
gMjYBk2aokx73mrW8UraOoQL+HXFol9Orcopl5r8/x0dJRQ9FHoNGkaUYJt/vLWW
SlsrQn1p8weFtZZYLcFy70b9hrckS7tNUnIhc3OjFdKJtudiuo4ppkuvU09e/rLA
bEe2mpI9jVqgVhIr/pfINUsLYGxvfa92Fp6txNP5U90GrqjH3f3aJKbWYMaP7cGK
sE4NbNJrn4cYDLsK/649xUu88lepTGHgGqW/1iHzaEv5tKzHwfyg7wwBFQyQ55Ci
dMGhpU9V3vSviDNfqVgNc761RZNndaJJ+5X/RFem8x0Sdv0SczYPL3zjJiaJvSW+
2CCErr2XhE5qW3tAOW+d0xiGam+FzZsO8X7qd1Vu9Rp7+milubZ3XBWdPbcH64GL
LagMLR2agiaIlTLXxcZ7zu3dnN89v4c1s0k9DDxC2SMYrDQRFm73sONN3MmF92bg
DJKIvxJWXAHq4iO52jYUhKLGDUwEuQUk/no7H7qmHy3jjSkuf3mp5DtkoRGZpehT
6949ZJdxo55A7a0gSQdIH/g/J1EQnALJg2V65EHF8gsdxq6pziX8gsqL22vsLXGJ
ZPxpFnIdUAhcplAYY2F7UqWwCpJG36IIs5w9UPZjovK3MVk8ZcTafjw3SK5Qp1Ob
Bankfm+QoYrYNfvaPVlSWJTQOdBn5HVGNiIfEo+gtLa2Lykp/V+M4GiQg+OG3uDm
cIsMIxIjJEF4gOEii7TobGyLShThfXJvMLYUtlgUq4lfx3cS4T71AZHHSYwTgyPW
aTXubDIYLn+HTQpUIfClPT9zv4FN4sGHWVblYcIL1N9JWkOalFU7hyWPXs2+NlX2
W1gMrv4jE5JaDRd8dx9EBF/s9KuWe3lh6VwL2qWMdNr71JJCjc2vF11f6E/5uIS6
e/9+UkBinNaRS/c9IhVfRt/6WPcIfs4B8Sfu0KFGKt7VnUdNIf5yoU0D9KEqx6HJ
49e1fXkIYR+aGDLUN4Kj3w8xbq0xRGW2W5gP1VTEeadWYq+s4Q4jJM6hfvzwaeUG
HzaaBCItYj29OAeBzh2n/AlUSkWVbTGVMggLU/ONcRf48Z1AFoda/iO+Z4QuaGLn
W8AC1Sf3kYDYnFzPwsGZIx1ZqFpmDVxP4EYs+BUDvJakz+FZxQRIDoeoKQT9a3Sr
oHtEhp7asX5PKQSaPLPp+HtuOXYl24sUYFw9VkA9bk1DW8x5oAD7fCLr5SGjzsj9
fzsYLhxSTps5H0wj8WT6RfkYlVRXIaYc71pNNqwTP3pVCAdfu75rNt+mQDANRM3c
MJzmEqzCD7cGcOwK8fCCanRFfqP3g385X1F8mtPxMMujjh9eBoGWXyRLf4m8jeUW
uF/8Gv5VTBztdLSRkf9T8A8ZPCsXaR6s3iCDS+pNodh/kmHWejFHS6eDmm6H2b93
9PPBP2yn9DaNyK2T/0Ov2aoQaODwnPZBgyuc5ZUbm56Mp1YJxBMkHxfIYnSNke0i
NEIOlivmvI41gczl9JMbRNWR3ppqYVaDw4kPVH+V9QVt+xNEA0ILtDHD7BsI6p3h
nrQweHS2iJmCT9NP3bjHAXy0HzS3NAatUL2Zch0HE1CCPDI5Y4P8mQz6j8rzFp+4
KhjIexXlQO45d7xscwigQqJXZNYxs8U1JqejVZZE0DE0VXLd2Ahau2yLotkQNt+D
CL2i1DfYwc2P3fs6f+D+tDNlSXb9S8E7/Vlh2M5MK8ThNlzDgLQVJEcEPRj42p7q
ZRNoB+AUCwdXFldlWLXukBTDErg+SS7pfrG1yoxy4lEeJjt6egS6EVJ/sRqN/ETW
5QDJUDUrhi9c3flPTMasCxq6ZToDub5OsQsF6EWceB5UMXx/f1z263cWNmrqY//L
+2anQaR2w1720jYGDf3Vb4IPH0co/twsu7P4ewCvqPK2v82aaNm1K38+XbvaIQnr
3urTk9xROU6rAE1xFeX28WHz1/wGLmIwbHZFiZgOH+J87tjknR+lS+3LR7jVLb5b
Yzg285C7YBXAw5DL5+cppX6izprcui4/1XVERowo5AkJnYEKMN7xY5aZXFLbHLoA
1ogVGcywGhcIxb56hHEbZlwnySPuXY/GLIcDsgzlT7p/ACGuYZFa+K+SpXGsQCQF
UAkFtVBJzRdHqjmmA6PUxb9PyQ8obQs+YbDcNr5UoaK6eNrIkh09UTUnrbACif9X
7j5MVKBnlyOvh2hmVWs/0by9gcDPxTNrjL4Y/BYY8v6BQEwBENZyjwhbCAujWDXf
AZizTrutmalZJQTYNGAgfafutfHJYYZgxFgcY0I2iJARaTpG0hF+Jk597UM+w5Vm
OTELMVj3vIUjqyymlGxVMbFcQNDNUuNgnoy5MGOqGfi0COzlFOruQLOLeF/Rvk/6
dZsZzsQvxglUa7AZN1hahqaucAsVAQMHotUiX1MfFctp/9nMr+oHpTuaV8mBUJM7
+oCuwjdcvmqxHTP2GcvzeQa45N1Cahwg0yKTGLkJXp6cfHYjj+zjENCE5vu53uie
d9CknAZFlk+KXmRg8MPRlhAVujFNIw4jVXpt4hT8u5Au8+zICoCfbu8qACrOj9ww
phRoBXVCbvCS+hBARtlyWzTqkHtLl4pD97/5me0sMwKSxJGloUne+Flp3iPuOlgI
shaV4Cd00L9BU3xJd+YViM8aYBp+ylqPJoR+txL//OCiEhc24AFhv7ADNinryTZm
mxht4gNU5D4jZVX7ygGAGVxDs3aPZVToaIX+hkLSbe8oORNWdruqmc+BEkrEJvIM
UbNnKWNFTMwzeQ9IC93B5OkjZ79tVcxJurxpvAmgemcKtnP2brIK0kJOXT8vHgEO
ukH7LAG8+zbgdgQ10QaZJy1jwJz5au6Gk2WJRCNsgRihp16Nc2ZOF3C9lmylzlsU
9+puHp2JCY7peYfUGuKORz+YNQbkAJaIfoAgPTZAWqMoO0Q8xU/AwDWk1nnFD9aI
D1uGl6pgUMTBf2JPjaby0rY7yVW/rSGgOlgN03eKBvsiL0qVxyjqRiHTiFVw/mv4
3FyXZXpZOZrUMpU/nbaINxL4GQPb3sxEH0lV0kRJkakjWz2W9yy4iEkgA20X5SMd
35Ca+LyRJ8Wufyq866LSYMXidfX5YsT/08bJjI9cLum4gV54m3HYOFy859qL5kxy
Xa4blrURq5L3+ha0XFITpHOQ7TEl2Fk0cKkBliH8aJEChaUgA8DPWW+knEmq70/S
qJ5at/OKmgsX/jzbfIb5ndyQCl35he6k1/TeRjHfBE2SYUjO8W4o9Xt/VUhEkkUu
fDN0GLvf7tGjkpvS1JJHw70uJVxokzH7BYMNXbWOLsAYMXtGQtsjW4jMxpBc67V6
WDL+1W2eSGuWSOwib9aPW8f+EQXxZYWJT7NnJZXFXuK/8XoICGlZK+Sy1vB2R+wy
NtNZFOUCt2huC0SRO56u2f5fcofwnQT4fs/lTow0FpUsueffkoW8A3C4WWXTHYUR
45RjBsQNV6azlkDUGGD99+eu4T9YNhB7HQcZBSGuCWF6Dm3XxoT2hkxM7xFULCbT
XQJHiSqZj4ewU8UnCZN2MDvG34Ak0sohkiz/eBRFc8B4FiilX77+7Xjfhql1+q0I
RGaBxk+UYyJkjzGPlV7Kqw0GPua99/6FPOJGYwkAcIykhJRhET51eOD461gJqTPB
R65dGQtFOeVqYLgY1xCW8NeJ+R+rijaXQL9Rsz0RWazX7edm5neCLAOBimVrfmBC
ai+EUkQeEIK/th7Rdua5fq0bTt1y7Rdt0aiUvsQoNhPqikc+OJRBhXxWfydvmiQH
ZCGgbfSATgdyKRBx0dl4F0NI+hSTyBNbN3GuYXHf7p3TqjBP5uLcesaJ1mGEiVbL
OPhxiL/ZuZekuZuQqlEGvSxj2zTtR4GhtyTH4B1BbpRWSpRV9qdMtp4SmhPacwcq
hQRkT81pN78uxjkT48BnCwUm0B/yMOmiRJ1izuuDgMAxiXx8sXXQo+Kio66epCkO
SsS+tMmXT5TypZ/OoZb30hXlbEsYc7PeKY4HtNdE364K/wVMrbitjygiS/Y/nPvo
QZBrL1TSvUi6rhU+Ilp4hbR9bMol0csqbRmbHmV7FJ21erMy9qA9IHWaCMgPjEDw
0R9xdOqHM35mDPcYtX31vipnuhNHkIY3cgedfWG2hTxV3Z+XNILp26Bnh+ULV7fv
m6oo5KMlTDbVuDBS3WyRqCn/+blwANPNdGeXp70LW9k8/j+5hQmHqzl8vrjjZzcX
Iz3pxUbh6RrFOKrkJ4/nHZ67jFmH6i6QfOSQAkIgt35Hip5oUN+0Ph+rLj6TGf0Z
X5INp3MfZ90r8jmYrFbwUCY+UoGJBhjItsVBiAcx7SpoEE2KXEELbeP+gAKAu8m1
nCLc4O/5FPVS9j+1+uVT15VgPpmfwIl6W6eiOynwPN93w0ngF3lOxw1e1NIDJ5/r
KFwokawk+azg/kQaCxclbNa5Epu2rKF5eRhTLirHmgE+f2n83zQXRc0wUClgX5rk
UoUEl0nDppVuJNeN8gHwBjNl62eH3HYN1y0NbhLes6Vw37EFm/fQrEAyIrFYva4p
kOA14d3NoA2hm2N98Ons+nNpsMf0RovBK3TRCuMKbDf4X9XhoETlmkvNHz0/NN2M
JecjYr0I8mW/KrvPphsxtbZ2lD+GEPY/og8SuNpe/xipY4dYArmerU4x4/B3hUSF
YPAHnRPoh9ESkWT6FucxrR5C/yd0jTdjLEvHdHr1Bj4CKUevQ8tsalar+mktIVCY
+1Yz1G9YbbKZzSPY6dJUIKortai3j9YqIWN/n/kF66KNs1V7BOhDU28IdhBSJxUe
uLOf+LpEQ0I7UZuBsfIKvsEVRsfPOoj4fPbPk9cGTJgb5N0caKBcAh6+yDgY/vxp
xqMDb2mi2bhdcsWzMasbYTeoULuX/m4YNGaDGItKs3EdIMYgvoJoU3dQ8VSDxAzj
x8pE51gvhQBFn7LFDirQjDnI1o7Zc+n9TAIgKWHnQpVXF+zJIvjxsb6lbR/RpQch
TzUIi0ojxqJqechPglcKyoFLvQB/Kc2tnJo6dY9BxY+pA4JoAG/kV1iQh/SubWms
zPZlv+aT3AqJXdtQBrTKqojqXjMG0peNUGQjFQ0aVQf1ZmeeoY7zwYT8TktIsfH1
NAZUpHQQD4MUXvqkiyw6UIyoLqGyyg1RPGeWl1gqyAE1Iw26N9quDTW2SXKubHf5
NZu/s04LOUL+krbIdZEhclW16B/jnwVACmUJfYqYFmKEHlhrGAITy2W+K+fIS6EI
mPl7ETBtIaH7dDgB7mXgpL1uOcmEbqn8+wLovR8yS1YbU7RavcHqiefylm116e4z
9/eRKNS0IS1WX2s7xxSvT2Ppf7QLIbx+rUK6yZ+zv8bsMRjqHxQZxY0ohxyYLv/r
4H90QHm9JDJ2VP4DRRR442eo1Ia5YA3HAUmARs58ZhIWo68ugG16ohnCWOryPoxO
mPPuiUqxiTTh0sJMiaPF1jpUh3KY63Gpat2tL3ggfdZ6HUe3FgdSKvfQA1QnwKy3
BLCxQ5Tm6RR08vrJ9t+rPJ8GTSFiDqphNRIYQVKr9PCTf2xfz95mbk+PIcFOdKP9
dNcoJ9GuWxbTxb5ZlIOCskvCDKvyxpX4V4xfiiaIkiqlwapEP/13UKsIT0H4nE6c
Pbnj2JHRKBewSRyrNOiWo+mWkzNsJY0AelDj8ifQZasAcbyl7gArp8V7rx3ADdqE
OtI0rVb+foHNvfgg47e4oXmt0YVe9OKGE8bA/Me4d3MDV/GnLa/rN9kaJncVEiA3
U/Lsyb+FTqsoyNPwgIX06glZ944HC8APV9rPZGyqvDbbinTDODBkR6psHe+Hv2xE
jHXWKgGQrD5VjyfxQ3N7Geuh65s1unEajT7g6Rvv0ZddMa/DFTq111BdTVuHq61w
nuP27HwaKJDGcQsnBiUwFpT2Xf9+bcOYH3huWRNNv/6QDWJ4o2irxJdsM9RmndYt
9DsD29J6QLClK4uAB/9EeeBHSoRMXV0ylMxBPAle3agQtctQHZHOm0iau/iWEjj/
zF4B34HranwTnSxsDkFXYn/Pe6Gwi9ZhjDjkFOOVzIZeMNsO0SJ0IJ7scBqLNw6n
xxbCSp8nCSXep/4UBMv8Og7ofYdzMOGP+C0Ob9rq+tgMAICUmeK/Mo051jPWYVk9
0Fg+Tnd2iOJ8UEWT/EekWxnCV8Qo2h82qfHib10Z5VaMQg5ELOgwdPWARQfnjPp2
bvbTszFExKboF+RovsV8cOl7i1mzr/+NGULrH/Siob9KOVTJVuZkIr3TWJX5Xt9k
qOjUtHIpqeXRIOMAqRrq7KMMGYJtox08xrywKiUK9vMP2HTnNL6BYyBk5KFK/Hhk
1THslV9HSkAndtQZfb26VjWjlXiuZM0lTWqKo+ggXTEJ1beULw2XSQDBB0y2hzfn
jtnSeD460m0oloksLOqFbkDeXNXoWzOK/rfjn2oz/mROiz4kRsJhBqDx0F3ljgyg
heXMO+lDLYV7euyjLzoGvdCK2yVm8slgJkSKgjl32TxgIe4le6p4Y4JsUUV5tKfJ
xwc29T1ZmtwNJ08TVHUOCPBOdulU06IwN9HwtBLLQYn+FgaAa3+UlL47+xvHGYx/
Qf4AOHjedj/TDkuecCAP7VdVwvyJD3RUnaD8IcgfJiXbaKFMR9UdDPO5EWlYkULl
m0KK4nNEr+F5dNv+zFHLi5+9r+4vj0ebWDhJfTs03C752Z3KwtN7Jkrro0gKPi/q
zBKu99KEkQIz1/I/lHW0XJBUXdpr7xIuEjfOlds+AMkZCci6QxSEIyZcj4pLNtKE
Dv81pbpTypsx0mx7k9pWB40s62lfc3+xS+OWK5sXm2uCpKbPruQIge79RQLA07zb
Ye3wLKzPC9TqQ2actGz9ea3/zaNgQwsRLrghRtFQ7l4K/urgd4iZf7bpPygY2Xpk
F7rKqKiK0z7G1Is9VFWzfyzW/039E6K1ptnawAxu+naf1RI2+0PDEO5VPaogynLK
aG+15znPgq8d/S8yneIUvw3ZPSQVo1tXdoF9EBtOR/fhW6EdyeAt4EUPOTH73Ac8
1ZTKTK8h7rUervnjL1h9ln5Dr6QidAp5crJnbs9k8QgT+OXy8kLQFA7eePC6t92q
ZFLbJA/TLL9ceyyGoujCyomM/YvaOourHG9y374yUl3iW3KIylAd3gufViE2v+Ix
yLIp+n6utLTsQXKGEOzopQtRxuPZN93toXQ9FltBC90LZZqERQQbOH6ca051J8G3
yT5365XrD0rIRTGdeSq3jnmij4NbX1UOcgqWjB1ZQw8Gs4r2eYvfF5zefmQ3XW3j
n9XLBavTBNphzzyWxcZWOKekeFMF7Ftgnf0ChKaJbSwDcy2zcoP2gCRpNstWTy7H
NzWOyk+svjfBIRtiba+w1Cd1tmmXv22r3B3GbbmH6NkbJZiqcIJIlhClzUcaLMQF
DGsOrsGe7bXOLTPID+frTOypQAERslqKMrMUT1c9eu52n0CUDWojRLBbXfkVfjjl
kc4MB3Wr59kB69foottbfKMxnxl2L3zp4RthWD3GR9ALYaOLJrA8ZnVi9OyFV2JZ
N32LdUraEZVxzI1+ykEvwGjjcbaC1Sd6uH80adP4VwFqu5j2Ft5yGU/ojt0srJAS
CYa5V7HJu24MnyQM+64x0zvFPJZU9MB2Gm/HQvXgZoiulrGv9OHMeL9zfpN+QY/y
wJ9sqL1DmiJKCwAR2cOr11gKwqZk8r/sbAqZGy5ivzlItbs9hr6citbqXDV8ATsl
2A3yO6EgzNpMujnA2JDMUZDPUG5SfZlMi2zZKP5fGzgPiT3z2C5KqtrcYhh6LaUv
fUp4u9CXWsOlxzZTTq+ULeVgZn7W1ePpvs0YW5f0hoJysLSBR9jCiMlYuG8xQFSM
lJytWG/gapfRrBexEuUqg6QdXr0NZOny6ynFnH3A3Nsilp8RovfEBKRNbLunsbWv
Yutk1F+2ON76R75N2PKRc79Od5FCvHos8V46lu4N4GoQWaZoorcUA09irIJkYe5z
KM7mgGAgj4L/UPZdCQT4d+++sqFIx7Qy7EgoGrCMGlTWZpg/y3x3ussv2btKIEqz
eBdr47hWZmua7cTfumPBcQVgVbhEXc5lG7GvInzVvNPRrpPA3hl9l9LRWtxsbPtf
ba6X5OhxgSY0DFwNuoYJfW4A/G1fbwaqZ23eQz45WVQYFtrW9dS4+OAfWdthey9X
7vnCDe9RWXeqavHH6/HcVEjN69uRtGFP1vEb3eVg4ARIfKY27gCb4Dh/7IHVlApk
23V8QYXGG6rUD9yo5F9l3LG2/QmygnhAb5/e+CmnRjFOhLCUNSZI82+LWBDUt/zy
+GaNFS4UDhAUNLtsNqyTdA3guSFvwxKQ7dy0ec5o7VqIJ6ftm7uW/zbWHtPDpdYH
wlOrV8wFSZBuOeAS1PfcPcAmrx+oUUOpg2v4iEfU2tmvwdnL25nsRLeiQHBjVJLV
KJ7ypnCl8HQVQ47JpNyy4KFcWKEBV/N1HLn3/Czrkh82mDZsLIqJR0bAiTnJtbd5
HFTNtt5DoIGCZvuEeHhnmvCQOGOxrtzgOTrr0TiZmdSVt3gJtcsMTU+TZ9rqSQhA
e923z5Ftov3Ff3w42P1Ed2BgNGT40+9DSklKH+DQvWUY8DB3LeWc4MKVl1jz9GeO
7ZxRVSkQaoO14vF4GrZTDjXmsylCfc66YtPPv7MKmXeW5jKHPWsLbb5/4WvmQKQe
oik1o0K0fK+zMnuXw1bPgT/IcM29vemn29PeofLKrD9+emj5MqzKFzJXVslPvVHM
ca6uU1XIQ66tBANVzFq0U5nQMiDr+JW6fQ2uufU0Lf34N8z/W08M5trurA9fV/IG
JWzxXJYeVIK0Kc3t7c/cbxCRctC0oF+6fyN1i7jjYjgK1o+5j3jaevT9oGVcxHp0
qFhlL529d86cLmxrj9ERu/dfpSJeLBLxwg7gk+PZkEdg4U2SPCbwAd3QjbtWvfZf
xNFLP8sVQmbRqC++F/iBwVa9SHyWM1sgvYPDviErQeUo/S5TuHG6UKiwWlaB4BRU
r6T0VHLEThidoudyLct3f729amjiHSzHvrctr2o8vXMgO7dytUBuHhTz4Xe0Yo7L
VVnA2HkdwtotdgmXcON/oTmoyWI/azqD0mDEPF+k656kjcu24x0MrDRMwqlHPaYi
fxze4wd7ZXhJNXTCgNU6eLyZXwdls2dHGUYKWF8Di9ULj8L7aP8/cdGVCQrdA7r6
uXTi4hhgh87cKnBExK6SCX3zxWuyrVddo1MWkoXmKZb2iTWkXSqX7FRMErGUaZjg
SsFE2iDrtCj8TpDzvrkM4/O4YVF89fmbIXX7xfhekvUgUx5b2xZhcSO/TwyT8tDB
qH0lzGytjSNx6q/DpW4mRFSK1vHpaWpjXBokFmPzbciXU7SeJ3TaczpdiYm2SHEH
dpUPZI6aeTuEFTFcw+p32b9YvSWD75lfsiXsWX1ybyP8xKIVRimh/wGJJmDfrKoz
6uE0gCn2h5lybQxvnviz/1xbBBLajy+1lcmT71RUr3ipQYyyrq+97j4Fm4rrfIVy
cA4QizOGRhSNUudTYj8367pYqsqpff9VymHYfPohnTvvAf/5tfApAVRimGj7P7Ra
2cR5Y+dqOTEs4Cdd9lJ3Tj3QvrRc/S0my8S3o7h8YsVHlxA6UGvDfcNhgfEzNtUG
w9P9OjyY3Mo/44xcStrN1VE+gE3I2TpP3nyMzLPOBf3fe44dvWHfUCKAfPtOst1E
pQKSLodjXedwh+vN0MmwQnOZFXzCycVRWVXxTgmxsWOnPqHLJq3FmXN8ztyYiMfR
RPTr2It3S9TYFBZvuKa6BrnFOpkgF2avlF1qtipeub+BcQwe/13GuQvhljcESSrv
leOpjBWkY7GFKe3icBTEVIV8RSI09FfD+xXLKRsf45Mu9m9GWOf5yU09YA5PzFsX
Wc1ykVa0vj/ekcoRiMtVSfyDbNOWxpxEoDIVQ/rbTmBsLCKutdQUeupU1HbJtQkd
ErGQqOa78kLMHPaVEhJ9IiCT8FW+lIV1Fj4WiJ7UiWLBOnW+d34Je3I41WLvPJRJ
xkC1hREBTw2uo/8dt+Rl7LzxEWhIN+kUx3OXuQc+r91X4MrVkjLHV9Gmdx7Ga8Ce
1Y/NIdAfnVYm6yC7CNm7+bWUHu/6m4CTZLCGpFxYwvcLSxmMSegtQgnjMwbhwgZB
gJ4M04cHWAfKcdUCFOGG7mBxgvvh1O9FGWCt+fGjqcXpOYkj16+NZ4y0rYm2VZ2M
NsnvWRJLDupx62XZIvejegof7yXi3LzcKTjBjEMp1Pm6euFdquKIKoOudGqtIuhc
mEqIx4jBON90ZpluCheymtW2mOH88GIbI8VtgmDXuMTGMur2WXjNJfA3fqTaJ2lR
O6ALS+JR2+Xq/BzWMxLz6a3djoo0Zy/hrlP2BKUSxmpB0Vell/3xI9YUzuvE7ZeQ
uyQlxGjVeAUQeTRj2Wp2TvUAyQbV9O5owa0Pro0JHfOSaP9Mh4vp3OZlFSHxPyHv
3nKIT7FD633Rw0/hrGIsdCDdA6+u7BT3+LCjqjah1dfCEBvFd6ppvXFBDQRMfGn1
+tUYX2G42hlfcEYae72wlVSW0acSRdm3VVdlK3vA6XdhCFHUasrhmuP2RLlmkS+t
+moFfRDfhYtyeVYmQgd/JIPHCiRJwm5jYZcTG4+kg2UpdMF/d3nFMuvSZvaR3q6g
nG97EM3pVR5NxQP6xACydcAzHfIt7Iaa+6ugbknKVukkeQyA1YHKzqEREpMUsDCS
irqQBOEYWr/SmqTKsD9I0axLN3/TfYU4FUFxoFzRhj62ZK/Db4WJys+5TS5x+tjl
kwykcF5NtMxQbE3RJEMq23FRaKzedA/MAZq5MLao8HkykqXBCU3Fu/eQlgaXoCXg
Ay4l+Yluj+tfwycnyZEIm69f/pdlk9g03Hv1hL92QZBNFAqck7YWJ0gox4pCbtOR
QxvfxeR55Z03O9xJZVqHuyqV0FiC0/c+XDZK6/rTM/DlmLHjuDi9WDJ5z7idixB4
EdL9fLhp47Qp5XID70S62trTcWgOpewQETyrylv9CC9PTTzm4bMLjJgGuc72zE8E
mnUmrjccOJj4GYUsFmq2VfgsiAQ5VjERbl/fFaSyt/+UYXmO1LtsLcsQcBzejqsU
jjSCPqUAJVUrVlCUOvlWGIfuesQADYMOrWN4FZQWoCUy3p1a+yl20oyokocNiqof
niq8EyuHKD/cPgmu72T4VZ8T4enWdO+dSZyQ9Y8nV0PUaNWsDW9IMdgTL0gMTZVB
tLmbUavKaZEN7ohrO5ZXgsBUsIlllXeRPb3zvemynbpU71SU7+HkvexSQBjzEiuz
6SRd0+pmH17abkx2Polp5bk0GrzWz5fsB2RM3rCI2bQZSEsXVoXPr1WePvNoPy8l
gdApqflDK3zF/02gk/Mz/C/3mdge7P6dckkamrvdUNXsBFzkL+iJDNdpe9Kdb5uk
6Mu87mTejfM9lYgjxQi9szKjs589PvYiOKWJDzb4deVtVgiw/6uQgk3KinNUbldz
t8XKiphQdRYOaE7RIDtjXQgKate9BeoVyCCTB71EBQ/wCJMHXuvLVRYfxjwge2Xg
2bV27atgW+2zD0GtKTue9PXGb3E//2w+5fPg3ie0oRVtwgnujQ/CuvKbJ/KKSweK
TPYZKCmxW0oKiKWhIuNIfGTOsNxlsR5A0Q50K41j7dxVKbmAAnexGlv8Xxsa936e
CPMN3siM0pFfhAxVSrTdSyPB9HNVI/ILbh06zU3VmgIPFN5qZrV0JRES6frMYbau
qLYE7CorCgp3Xe2IPbKtTqIIy0ID8P764VSaaZi85ltbNT7XggyW2pFLAitsIfMd
w9xpIjYAB8S1dZoBFtCTlY1Hyar3HS3JPpPnoof+jGMHWQU+h00Q9ByJy/fqI/xf
qXoMnuiAaUcGJGkPqdegeUdpCRS/Hff4XSg6Tn+PAYQ4yr5FuJcberW/1BV9Zx7H
K3SWCm/w7guEvt77qtfUEN3FVZ3K7SuPkrqp3FRZ94hG3N2A+kHqBbI9QIJnDROe
a3f1aTCim/7mefJR5KEVDcTt+JOzHbY3vxmR55qT7epxKrh4GAR3NGEJn8/6ks70
KXXQdCF8AXQV9YJwdgKpwqJcsA2Lmfndc21aaI9/ZpQsgd+H07Xa3eVar6TBEK0e
DqSBVIi3lWkeV3/nkR0uqqTaTWA3ceo99pZv54Z6+ZcopTcykgJYI3J0zBTzquDW
A77JHRAGYA4DXdH9LXpk98mvcvaO/o1hgP9nU+eXyI3Wzfqcm3O/HK6aJZn7sVz3
Wkgfq6oQYBBLHvAOYBRqcSf8G1r43LePsr3sHENLYCbClkaXHPLvzpSsdzs6cnUM
L3BMU7dbE1NXAWdhU7uPks0KiLNBif4yZOxw6tZ4iWyieob0dvQA2pK53iqmP8by
UcNKh3yMj2/fuKHZgJkTsSUdI0F9xzNzg8qL+bKf98OSgJOzVFEmq6FgNJobrzap
Il7V0wFPWjjwWnGkvyqAmui99GaisVzK8efUWaDwAXbuT8j7Kl17R4sO+PIR3HaG
iwgApXvZkY6eUvb9o/rNb0oXN0yJg+2oVBkV5oHIE8wNS8hU9BYIQuiJYBBXevxt
7vILcxSPfxlJJDI6bBjFqiLg+WGxZKJsb6+BaxulT3AUrqgQA6qd44kG7iFg1U18
Z7NmuhlTZrcT/LtN8IgPyPK7xiNsuSmo8GlxrG4vEG6YsTOGY0fvQ3skiwcXx1cR
0xL9xzHQMFmZsbXnGT7+V3YpN62KElQcuASYAeshp/iQDob++VdU89om8EAmRij5
5D488WKo2gnQucWba8TGhzpccn/HtPDkNDI92uOjcuL5XcGCslJrsc2/zuYQoiJX
sEv6BQvnzsrH9mZLxXXPzfPaf+M1KPGRvfmwk/PMfDNaw7ZwjsSf3snmCl6AVftW
XNcz72lLs0bsz2zDdGV3fwobkYFJIT+hVTY488iKnckMyP7ftKRGz5Mbcg6ZV5DS
JBnL8FjEv/YyA8d1teFIsis9O65/odGZOZFcHOR99Z5qCKO6lhUSYqlL/NIkF2ZP
vHdOGeZXHZxeyr3eyHOqOEsXBAuo11ASifri9PsKE+DzA0Xh9Kh1TCyAX/wyH98+
NgAKhbT/CFdirASKYmU1Y5B1PNEIJbfasa03BphwnOlq0AbZU0I8y95xIOumIaaC
lpc/IyzTpRaAvKHbWpLXvzhLh1/JYA6ENV/5/BAvmns8La2iH9I0O+WmWcf7xk8I
DtdBerx910fm3iBpczkYw6dft2ZYrLnMqflGvkVDsW32QLK3Iif2w6TmapYGJePM
ghwmmbgMufMbkKpRPDjlNe1NwDGgtAKwxvnnzzC/LN4uDch14msSvbwB6+EDgHxc
WPuj8rNj6+45stAUnmieFmKTTCGiUWKe6khjo6bQzRWPkUp8BxDITWNQX2FRonSx
3QT8HabPRw/GGPn/fZnhXEGi8VdDwM96vL4+PgkhFYyb+KFjCzGRhZTz8rZPzhoZ
RTtMFttE/Jog/dkiqRggVD9rG+HfS66TzmIi/BlrnvqgUIuLRfuORU4hwbKY/9N5
tgJ9rZtBDRTtnzDBzI0Fy6rKSLK1MoEe55TsiBReHD9Fn6GEDeKr4NaNjSNNH7rQ
AAcMsX8XZPHIsBb7CrBtZ9yG+Ey3BOeYi/uZP2fQ6FFvXDpPWbDLnOgRQqSSlusV
9XLOgiKArO7ja7zyXbBqXqhWTHNyxqnO+JiL8Aclfsglf3eIkZvxns3ZYPveEaAx
u+7cjgJeJvxJznFjjUE5j/1dN+t8sTHZ0Su9ULUS+wr0LQC5Tnog6BX+8L2vRPPd
ar3eRVgCzGodYfBaj6ZwzmpUMWm8kGKqGH5ZB5PTLcuMHbOL02BY4ndk4ISyaUM8
XWdf2LAdfQPBb9+3MkaD4terIyTE0TslwJAxkyzhffH7f6PHsygu787KCchLYAPa
GllWhbwUdj3SBorIQceDAKFV5Q8L6Dk+AQilt0YRg84TgizvtVH8r2EyoogYXDhO
OuLGPdF0rYyirOT9lL94/LnSeEmneys0m96xOwnzpMETU4yrPFIIPhWBobbdVbk2
1psm49GnLPd77beZpB6DZp4IxiPO76//hXT5mVcs5RQM4saHepr6ELjO3Nolfgjs
Xi2R8DYeXPl2dcoxzDmb2aETRMEe2p9JBA0qONzbOqw58Uh+I/4pNSPuUPCU56L4
0Yg7OVj4FmnirOCjGUmH4RvvKLJIDjDn0/Q237DCh36jgAs0XhZJ74JbHvV8PqXX
KY2GOYdFbPaOTG7epn78hpRflIEEAinXzSDQDdHbmbYlrF8Pq77SehdHbbrmQfm2
lo+KSUGP51zH/2Jb8tVv9SaKSZX7TZNa/+Q0hz689IHruMqbgJknhIrXASTXECrR
NlwKVV12NbKP/SD6HIoruBsiRKGe7e7OHEF5kKe9Fpum0Jy8OwGJwksL8OBwIaer
l96bVD9WOQqjFKuG7++RM/HWTnFub0Uiu2HyXdadRrm8f+byBsbdyJVYvU/8DOpw
123+QxhoFp1KBHeQMy+ZQw++z/I1oOLs+0yb8yv7LjkSwRbTfzJ+kvOIvV23chff
SswXkKzVIujZYTIwF2mYanEGKXH2fgjlqu2ze0MsrN4znp4X8baX8ofovmCCIj75
kF8glwh3MEotJXheQ79FUmvzTcbEbN4H9GMnr0HfS0rmkZFuSn0MvPg4fhQNFvfw
HbS0JYycal8OnlRYkVpIOWHxx/Nlz6AVS+anzIVkfTr/NB33LnpBzi4bkptnYVq4
DJSOyUSApeLihKKCCiCUNbQ13UJVYqgyLVeOR7jS7aaWkWTBjmLARvwQcqTpYcjW
KexSYU9Xh8qYVqMFysBjdG8kX4fgn1QdCBQL8LIxoYOFFe9YbKUDUr/tyyHAZCNs
NGtl8Lq6aU5RgQR5sG/GOiFaZhX53X1cTYCIOUvqL1HllcDXWoIfz/oQF54RnH4Z
LnHPz/gTht06QgSZ83SnqOL0bPVh2lSZCUGoHS6sXDk6npln2WPP6uSj69tJAUp8
IEU1EjkjJsBcGQTP75IU4V924CsFyxs6uGk6a+jZl6QhEjA6JEmrKtzdfd4b9j1E
87pOr/qRUx7ZFleBFrDU4iw+vcurYVB7lJivJ7+YnPDwceDX6yMYfm5kN6EEWjU1
bC1fgAnnYOj/k+aZz92RAM4i1pKDMaIdQ+v8N1lX0g/qbEBnj25EobciQe/HYR48
NzCJtZMQXTH14/7zCTl6akmFmjG8Z67WTke732uFsH7EHqIuZQy3a61BkSp9X9WF
eUqn1ERw9qGtEBEWz37dO5gFLcmSRxTdU6MqwsSFbAjCSeLYukJelK8iWh8v4CcY
8xIksnOioe6hqrga6jca5xUeyL//+PVlAjC9iL0OWMfd6z64FCVwtLGbZj2csxpl
VDu3ooxzCtMz1qUvb+LoBJxOPr5tSgIX2rFgoopyutZ0X27dmfyJLPQQRmnnF+GW
WOvrCppT3B2zsMFC2B8++dI5Dz3A5LR9Pc/4adKzoXzB5ZXGLj8OYhVhgjfMyQtT
eGGC4OeyGGWQdw6sNCpGLRBS7FjOlcclQseMLeh+9NGxF/wOD9bHju88/pasWMPM
ouHYln8rodsi9F5puncYnQeanyPVPVTFdPaIRKjFfcXLOglrK2BoQLwGeD4MjMao
JJkWMtnGQHnlXENPiNXg+2pALuCc142j6bb8Q+bbUq8NU7BlFc92TzBLnCocI468
U3gdylTlcNDi0ozujSSED51JjxghXs9Abgla3Sy6cWpaIf4uB4hDUFN8AVQTh3Uj
Z1MG3MMOUQ+WV2JLHEgcmhAMy8PGPF1hvTdSho5g3tXv57RWvdfACjhMqlMsRCPC
/TdszFxf4uTZqMt5viV+omTauAvZ5OQQ5IW6Eb31RgrHMMj4mICV3l3iR0ZeTtCQ
OmZop21o/qdEiOA0LpwMR7BCFUlRpIZlepRurRdhg4ihUqojnAvaLDteqGmHcliZ
iu7BSDWxOc0xFlceHqecxvHHsg+6uGR3fz5GR4JgBCoWGKeKopoRw0uQRghFLGD2
THrqxOXyBeZUL0awSCpDnuuEXF/4vw0xkPNzoQDNH2sKAubk/EdoHohTb7EtcCp4
O89pvm7+vX5RouMuUuFcaECGaqp5W8oN7UcNAPK8vlFGzWkcCotlZzubxgTFSrNz
U6cE7YtIsvDbKbAd8dh9TGm0dCTJfhl3/YHGqnJdTHxGHgpQ7fCFB2lRMiAHN2UI
HIfh43e8G66TsexvmxUnyGPttnXpGU3gISX/hr+FTLfMWeS3QozEPkMiWIKAtX7t
zklWdeVrEorXOmngBVrFZ0sDJleSv5CirHtiYT1V2qNgtsHWRr9lmOHwJgATSqbQ
uG+V7se2Uki/Nt/BfeAN6yUGRzefqYnWUXC88xnXe9DlpNPgZkmPSY4NTmGBeesd
9HtSK3STmx/M9rcxl3NDPGEwfYwMbARY0UXt7WAD1+ZoOcqEUPWLZLgcOQrk0BFY
p0i671OfKoQN6EoojB7hVEHCQ9Adpp8fjJQiOq8828nEX3Ti6WvpoYrpfrbw6hv5
WKbS0hqO8DMn4inoZGiiqqessYC1IDfzpi8U8EXLUNCbi0XP5E6bmXIxeVmZ240x
Z/HTKOFOwV83Pnikg+p4Tw5NdCG3VYlv5NQ6pjJbAIrZnrb6CiouyGMC4k59MpPz
ZdzIXAUDGS91qoES2ee5ouIp2UDag+PQUv5pmy5sxwvS8RVNgcMOUUAdggrGFDIc
BxLHDdElKqtK08tlk+0MxZ2La5/X6Lx1bHMqSGKzEC4UZOEytLwZKFOUxJ4mq0SC
KplscTqH5SLaDWc9GjeScV6VamDv88yT6JUH9lwDBf1Z53hG9+GIjAvc57aVS0cw
r07p2vSn4foIfLxZaCKeJM7/7OF+Nw71NakjSzWUsOz7hp0iuyVRtityeniQgBny
1qtOlXX/J1500nLeMroWmS8oqwOU315QKZGXlk9MTOfIK50iyI57/GyrnIE9352s
3aLl507mvZLLnuFi0v7t3V2IgIAqg9zb64I8YXYcs8PpoT23CfMBcE9GTjOPjuYC
T/QGbpvTt/XbhLh32MS9S4j6Xv6LbFRi/GIGShzcsZQSs6Du4QrVNd74aLTm6GBg
9I56j5THt9iLPlX6uHmK/4zHP1kkXDHgQaQbc9IzSywsGXI2B56pENtngJrKCMzk
WF/1ZKJMKVS7gCTrKZBXndzpuSnSrHB35xwJXenNkaQsl+WHOEv6EeKDQv+iNerq
cv4CxDRJbWEKRZtwZS6yPAvT6smv6VDIBfbPW1+UwTXfJZ+YRLag1BPMz5cCq6eu
jbBizZkyDzyVvmsGCFwqCMSAfb2U7+oQnw8R77VI7r5iRY5p06FeyWt2+nxy/drf
eWSByTTwVlUz7JUVdIHho60aPGDRTUHNMcpcIuB7/CpvHyFfgRWZqyAku21j3+Wr
/eKX6plHKVtXUWNurCT4H3AoaT+A07QzKeihgIkuyK4dxchPZTxko+X3rxQ3a5MR
l1OHXtbkJtSrfkTLxQuY3iZo5Kgo1it2FM6tf3vjnSo0rijIr+3z4JaAi0FPa40J
mb0+o+uP4SkWjsI/npfz/CY49kqHk/FRVLRqx4d2MN7fBm3yJjwcxNAySMo4xqLJ
1JYJTJFeD482OW4DjsxAsKwO9Bamg+GLKXEYWkLv9J36mIQS/YMsabGp7TA1F9El
iZxkFlQqoYoqGMzOPjQAp0wP3ZLr1vzJZlz67Ba+xyp3i22yaXqcimIjgivco/23
20vaR4FHi9l0Ybq8uE4/JTqA1EaIhxlXlovjmpd/TZX8PoCvbYjW6KgL878BawZL
LZ744CaGSq4ioRrwcmEQjrcEue018LQpUN2C+q7XywHv3OW2tMGz1xws85hgWxXe
LrEXspTXv777rMZGUKORD0Q8VqT12xHhyzLt6KA1R0QKVT6GwCdINffV+7eGBCb+
nHoxRPtI6rd5KrIZrzrFjhG3idCvyEYc0JC/B2CHJ6SzNg8+8Qs6KBKeobj1xXQr
rMY0t1/YXOwIMj2YqZ4VgMY4x/zqybgV1NmRyIDGOatOhOBiI8C+smAleVPn8jqQ
W7NDytWIQNlO1i0Q4OeftWkyWFRYv1QJYg5j219en/B/BbIGqLl9Qh2jQKEQvDbR
fwWeIx3uv3lj/UhOSvVoBjb+PXRFOkGsnoF07FhC4z5B+BXLutTJpzWNtlIjZNsJ
grZLtP2vQmoH0SIuXbHjsHFUrl8FKOZ29KOw4Sxvt0J3As9qfYo44lqH0FMeMSDT
VwwjlXYqaJGnb7XU5sKtC63TP9hWGBGYW2t8XX5WGIPX/RzCzt9SUQoV1IWxqtdL
uYaqWahWDqpWEswRE+WKhn8ppuDjR5wVSoxNqTnAx4zsR6LbfG4VBtil4Oz9Zj1m
s56QR/1dQttG0zETmS7wxTecScLAs+YAO9HWasGFbesnY+Oyb82G3BJhK/EqPNWd
BdidlzDWoob26MhoL9UwpfsnHOFJ6b2GGzqJkImoI1UQkdlaDT4zqBVHAphUbN+f
99iQ7FPfYsydhADmzelBZIYO9CywDabQ1U2d6Wf5RjqggSWpEs6UHjtgYXMFb3Gs
+p1N6X1G4yDHG6g4zkpAcmK44GFI25Wz6PQGFGjMVjOL71a76zwO3V54kX5t5wJX
bx+Y1HawS3K1GGcFw65lCyRpxS3tjpCs8niXia92IyMrVO9Szy7vvAxyHvCN4Pp2
dUFu3oxgOqsOO+IrvOgCLmJ5qr3Bvv9XFXd56zYpF35SnJ19jxQ4FQxvSdoMaAPg
NyIONRDFRtO+8vk3lr7FrUkWgyew2vzUkhc9V1oo2Ouq8IEJzpXw0oeXU7Q4AD40
Qnrl6mMVgMaSmppBvmYN20XQUqYEbJsy1p4RwGht5z8dwwG4Z6u1SSYzni8F/gQ9
vGjOftc7uYqFxmmY0v2GhzyLuSyYsUsm6p8DTRagQXmjc/whUfAiIKqvTDYNgKJR
mL8KJDqzjOFWUrOYxkbotP/eK+DXRxgDeTYh8jHuINu+ZOUwPDu2U+hk0ln5l0+A
fowomTaghNG+4acCl7Ik1O3UXMB68Wg4Ynv35TPy8g8NrDD2xsnrnYtnt8xEsL9A
YRuN1Hl91gM2zp7IYlElQ7f8NMu++RTaRSBQr21efAK4PMn25T3KWI0A5dYhO0Bx
Ctn288mhF4ydRdSb3vcebtMlHNRkb33SdyCN1mRMN3G1HtSTkj23WFBm/kDANrdr
BpPS187celj4yIMjWVGDyKHh+KAa2IBE2nj2A9ZD72cqlVX6EFg1elUg6UTrBFtg
Pau36K9XxSjbGktkV4VpWZw1cpWGDQXvFKFrPCgkhuy5xIGQd6hLhcxw0m5vzDOG
BJkWFms7fewBxo7TYp8lQS/jICqTt24EAROeeY5CqRUVvQoOottOZN5oeKzaIbbL
BHKK8ZTH3yFpwmGQBvghYWUONnHsBGfvH1bU0mXif4KePr2TkexWz2GabZjgK5wR
9A+7UjKppnTa2hLk9ZMGxF+H9zU4yF3EQ5JC0UKPa2tmbhFGWYqAMi7sl7bjJtZt
RhzSysaMFBamhnPZCoq58Kcc7XGUD8K42pTAFfZY094CgS7/54Qb0V86ImOYhUQ6
5l1HjznHEsGwCg+n+WZVAqAKfalM1aCsNQ796ni1dDC/R/WGGwUxnFAq2AZFviag
wg1K2m9RN01pvsmtK0k18fOfgKXEwpzaBIbrm1z5PlIHJwf6TXXtoIpAs33Za5IJ
KqDjwKfqXNaLuja87AN3HJyTA4D34aL7ORXOnR7b28kSZrI2T0uBDA73yE6d1K1r
6XINONEBB1md0AtR2H55oUypMyFJGV8Glad1luhKp+2RE3nDXc8vBnLGZ/faLdgl
ds3tA0d+uX0EbRUjRaMSuNXLuThSkHEqlBidZe2msaxZTthf3QmxpWn5JFg64FQx
Bka2DveioXisWqCaOnpYtgAGbU4xtLNS7BwY+9KGOswTLK1Sg9xuSQ5mZIZ7x6oi
2t3omHd14PWlscrFghePTp5s97zI+pbCWwq5mVukySBNj555zhudYgLqivRQ031E
IEANxGqUujTiVoQyVoInS08Qo1nANYC+ULqk+a0Wb9cT3A/Ndrm2y3nvfFLSd0Jq
fVgXZsr44EaLHwvcq1gM1tqZYvJ/4QgbKlwty2vMLZvYZeCw7UHOZ/8aMyPKMEAZ
3fO1WcMh+ZDk/zuNXoonZvrDPkUMh90xUVNY7Y0plpDFHow1fjI64eGvOij0JXbX
jSkAgAJT2wHu72O+4XqtQP8babjeXjJPfOV8Egy3lZVFfEvCTQh6PbOwlDsygHYy
JJowHiadh/XSrsZgjSpyUuv3sW+dzKkZ1QeA4vf3z9f4zempG+SbBBxUPOZC+Ows
MevXbBtlYJQHpBafCwhIfuJGRawK50+y53JK7pcQW+KmdjWU3zqsxMuGDllFOlNc
fQ90OFLE2R64kq2TAN1ID6/4WGKprOptzypQcH1uusTUoxwJWCMdy+5xl7eaABgN
0nGiw0gh4kKtRvVJtjvCkbbU6k2c05KfBJmTNpn5GVmn/fLABSMGW8jhH+qR8x0s
G8YQR1phgmDgPh2Xm5WEUX7xU3/gwfQWTI76AyLF6lExqTdj67kyXVV+ShKmr/2X
sVmDA2a+UsA+s5cX3kSVwbo0abVEJh8GVP0Cn3OpmVBh4ePEgtuRp0SFeuArNJaI
fj+qK95cJQfeBPEaLrTe0Gz1LYRwinpEcrgB4v1Wm48L7LhizyR6N4O3zl5+GtOb
s8N9Hix3DC1XNyy89d7g2D+GLay4iPlIx/wAGpcTIOsZcP9qOr9W1ujlEfvWfWaO
6CcecCC+z1W50ifmBBu+iah0uVEpHZwyF6wWPCXQVTwZjuYo3tooDda1lzOVOySB
gWm4Cugs+Li4jAz6ChNAh+8NopyB2IJeKiKPe6I014HwWHX/n2CFbEhjNMI1+zGX
tPBxeByHN7ibXJFN5u7FbdbMwmnDL4BOMZ+6AAErAWFzIfxOejE4id9ZOBQqYuFc
kmZKzMPporSpysoUbSdjBCER7Ppl+Do0SGVoFJJtpvO/Ik4jUZR69mFNW4bY02D2
8My2HogbLFDydEMmh7W3qG02IjETSp6gHTy+TW7on4lsQ15xWmuvdx+EZWDGHx4l
XDtcE7/uTurOWnaL7zJ6EIlTzBOyR8fa/XDkWqGYJ0yGZEFLXRDnq/1XBc5w2XWf
tmJXLglM099iH/VwmmVlx0LysDHftd8CBawYx5B99GNK/26rjCIv+LgVlLH9KN2p
TugwB8i9lpcstyCGvLJ6lDwBiDtaPUIH0nGbdCk7QURefKh3pMBqC3QKpMultiTr
KDmVZVnwQNnzEn2KB/w5YkzBSAIIBPXo1naBQ/oXYGOGXwcRgtOS3DzrloR4KTv2
Kh/HxlfCIpYVD/Mrox9ydSE0cOy/uXm9VWefDWZuruFqXBCytotZ0etDlX443fdV
2YMyNTChFq7HUEMQ4/UBbF+rzbZvN08QV1lcfV1auHMHWsTWM1Ix+jRkQCiAW0V+
Te81Ea1aikpvqo9dC/a9WwyIIDQvPZX6xsQhh4k1C6ZGowL3DOzoPhy6jT6VAjn+
ux4CVla1V/CecKCyqu0c731yCCxoWELZnPU7HFsfPDvqcHBV9Ggg+AquYLeva2DP
6MnNaZxHgbxdTcbCrAslxHSfPvGqPk4+GUD0I6cv8Kyy5hemrqxRbJGkrpcfAfIP
7HmnUimh3oNaaZxYUr5tXdu9zaoI7G1T8N48acRinj03cxPoxvN4qa0aeI/2RGrU
LXrzHNp5VnQ/rb5NgTMeo4kDMHocjjV4JibeYanEHYdkqNHQLoc5V3iIl70iphtu
vs3vjch3CBpvs2aNbEBl/NND/dX7HnEnB43TPO1N80yK316Ig/w8hciZY5jrZaV1
ZaH4FZeVKLEgqrrgkuaH9ux9PsfOff04vLoDMoISOGfI13fbvGlBWZyt06GU0+HZ
s/T91SWjBZiHv1Hb0ig1QMauxjOgjt0L1e2VbZkbq8MImar/uVw+L4M7gnh3htwu
wV4KRL9z/i4yGKnfNzDmb6pSukSD3eOdvhtndDzFQTCbWdSaSD/nEsZyihsJXr1B
htgrvAy/Bb7NNcuah0LLJwcgKRFWWBl/C7pEuu5tW9+HdrcQSnsRN3TM2KQVRobs
uK3LZIIo2PY94zDgrnJ8TDW11KFgpll5WBWRjLvU6hLAJ6s1IygzEyUJ+Rcrj+ti
X9ZpnLy+Ftyt3vjWzydGkXnr6RCJRn/ImDis+p/4NaSCEGxxmyT/ujRZXWgQ1nLt
eHx/ag9XQjKvVyZvTsl0bt2YlfIuvSWNluMi3M0i/LKamPN6Xxb2DKa//mOdLKzo
/eTq/x1NciUTijdbnIJwWqHuHTKffGIJlWI78uVHD1C+xyoiyke4dwTEp+iNL2E/
P53mtqYQtHm7jWRkW1AkRGa1hSZaEfktMRAEt52qnjCuWw5ZUod/jjFxAkOQH//L
6hlPNZIKeE37E5nmoOhVi4Fq+MiwhhepujCKRPNaKcMwmb2LoMzXTWMNCdoqwJdI
gYWmdPQmXT0VQJuJw5acNle3IpHUyTa+n2u5r6gjamuYNxuVXNSYC+MvgZuiHn9w
tzOKa5BY12lPO+x3VA1b4VAZjNHM6tElNQajczvK90cl5NSdS1qtavJsiSxcWr17
4PHCidXhae5gjTD59KXE1rXAZDBJ+/wluY3eyblEyeguhISSS5NWw2ifU/KGelbf
O8H+Gr37ab2KVPD+pvdqZQ1jzUCWesk/9DkPMy7f3k5XKbW7aXIEvbiUb0V7nC4V
LSddqnbglF4Ii7USdFq1jdHyY+VugfQbIRUL6IYFTJJLxltRDqhZ2OU/2UvGXF+b
Et2Fa8Qa6UaKABPSvlHhxqtATKhlR4rC3qxh9Iq0ZAb/lLuDuI9H41j1hfyA1Jf/
6OKlR1n3t0vEhC2xz9ELnQ8/fSHBQ8R7MZ5663ZC0I8DA6agfPdX1UVAuNrXxAom
xkLdMVbSeAfCAcNn3P2Q+2rsfCX/hK7RPr0Nn4h1V6y/dkhST6vpYfnRi8LlQLtS
Ax5fZwcD+KtInbkq9B82WRJc3C3IGmq2XLjUwH77l5w2x1UiRkBDNSMfT9+p4sjH
srug1lGUTfs+cNRGJDDpHabskeW76u8XSUODRVY+RK+eIwpe9a/RcMI3QDx+mMJk
+4AevNAr0wTtkU7bldJQFEq2MVUdLFP266dvo7FwNpXMmmYgDa/3U+fJjbAhZytQ
P+td/Fz88jnCgLnJm7KokKgv/GLkJjHf6YMO+bYtZX54dUHvbPOnGTH4lJnxWi0B
hTSaAXxAPbtYLxYvkuS1kRdiUjFLHiLtxrNK0uM6e/BiSi4flXfV1YP1Fsi4WY10
dOIQxevdTuUt/f1VWp6ndhU5VF/SwR/6/bMKBuZLy98Rrqcx0Yu9AKtU6E+dv1qf
rJsioo81DUjYwQEhpO/8NzZwy/P3KqFSf6H3c6OnSjkHp+45ZFU6Aqq1fR3ZF3X/
FceHe1C9NvPJjnH3YYzDSA0QHnUpZWH8yi+0Pt4Q5KIdOOqFRWOpJ6wDx0HUpSeS
LdwAMOuASKRXjHfsRKAtb/ttpLZIX3NqJpM8Hjb/KV/0NTp1GJ2FLeuoIzqMWM3l
i1Nrm6ssjfRU7LiA4m9wxjY4WWVEu56yDMqz347kAKusbg2f2PCeiKMflYeM+rVT
S2gegFaaSmF/htxAE/BknV7nOkxI05RC4T/ljgFHeuWIgWU2S8iqmsl+/4IGi+U0
+CqggLHnsHeM5HcpygjzWPOSE5coDJCLlsXg3kMmAUOudDnEDswz908K165zU/SL
EE+jhxUpnAZGYd98c3e1jfVHC+kvI//Zm9lCS9hYFh+UfOvVTdX+PrS8+Jklou9X
VuvVkkV+88sYUeHJZeovubv/VJ02pfFWXHwwyaVEVKuRftkMjPnpqWcoHzRLY1x6
YiXaZdom4O9aNUb5yPPPkkMHANY/6QFvrhHO5Si7ERu2gU5H+l/8a6IN7PjmzLiC
SibcJPoaZMfzLqHYAmcAHpFLJgWYyD/iB6bdz8VlGjpTUlHEOBwGkKodjrTF4qDI
IP6nLY4TO4sPjQ5zMlDlbvjw/qjnszD1p1ptC+16oR0LWTp3G22nTVMqg33mNIya
vjAsQoQ5JPcw/FsOzCWquN8THYXJfnYoSM1mTm9/uojpW7DYww0X27zVY84mHu/+
b1eqyBbV9te6Y3MNZIjMQWUn1O9rG87MVxU286iFprWpbGzVSuV62PFEWro8Kvnf
Daaa3p9TBgG9DzW35V+U1P1hbVGCw4rjpy6eXc2zKP3qlrO0Hf0444ldgLWdVG6q
0ZfD9bySo5RqzMiyZztAA3DmkOPof81jyyrteKCN2afBAgXrz4YYVt4x+Pt+YQJu
WeI/OdskQstVMZvc9oVCMf7AnuI088POTllrAkUBTkGkxkxUh+eJWgW7VlOf9p+2
SrCb7TJZPoQkytQj4G/pfcYUpGad8CqKpGgi7IUfHYqq+TX0hvuDw92R8mYnbMGH
055IudkL92TWP+aSjFB+NWAvrJtrnWOTiq/cBr4WtgFHX9pUCrLEF8NAKUMMTZXN
LIcMbS5fRbgoI+gOJIcp8PLPbSAw/cg/dyUizDkg+VboQix1AuiG7PO/gH7PwrNG
koRFldzGJDK209hebhvMrbjisevZhGjHWrmwzQ+ySRiAXnynnpAXxO9oFJbp0l8s
AD+oereCKqpR6INVusroJRIH3uDpBtFVUdg5enzGxjEFG7Q9SDk6GfCgovKhPckm
TWqfY3Kd1mOX7QuX0qyJrkV4lvzOveUoGq+OR2u5oX9iXjAkMC8OcgLLfAqU0k9t
f47GXXykOtp15qndubZO4cFhuK8djdpRfF7PONmQFjG3pKzSV9g5HqXYf/EacTn9
BxaMCVEPwFBlij0auUumtS3uT9J8SJMjnjp6jIiBO/zRcnMSvr3hiQ9bBqPcZxna
qK0/t1sbtf0GmugsbuKml55wGlpMBBR7oWlSIZBFEeebCPTgJVaiB/1BjRQVjioI
HTuEyNv+xmna/dSIO+dbk//Q8JBMrUja36rCVmwWM6B3/D7Ojm8zeKf9BNBj6fH8
xRCKeps4nOC3LsbH49W+ULdMJdQ6jzDUe+5/8QYp6GOXXd0dGDVVo2LMo1esP0OL
o60jz9I1Tpn3HS0IX/DzRrp0iIVy0G+Uuw4QLvEC5IQM+J80XrlEAFzjS1gPlwii
8lx/hCbkg0ylEyXfuQG6pZqsTSrHWF0UqHk/Idisa6OuVpQbkWE3H/3oIn6EJ7ub
aY3KBn75ujysqaMAt6AH7aEsg0jHcdoqp05kIBMAtua/BCs8qSMQWGKLz2WWcDd6
wuZuR2X3kT16WiA4ICrozKgJDGnqtY7fDMM6pJP2sU3fhY26NCWbCtkLPha2dbth
GRUZ/zrpJ7qL9Sj0DNwk7AL8MDKSQNR/q/JNt1Me/utYCWg/bqpZ1IpuoE/Un4Yl
PtHoxgrDrB7nRen+bJElEaxvV08M01Hu9YxPyt8ngB/0edDcce2ZRdACVpkoZ2wA
T7OozCMCJ/YQx9G8FzdpDdHjVV946hFcFGrq9dOe/yAN2uqhfrHhLzMjrbQxafaN
Rx1XhfXwSpS5fBcrdqvShqK9OIBWUe8jzDgh+UWCYk/YVqirYmIOjQiL8izdOvfl
dtn3f6A60LqkvwLLMzQwjJrfsTZKhwJMm7/PLJnvov6ZTX35YTe3MC0DpGZekeSL
VF4c/yk13DRj+jrPSc1EQ8Y+gFbJmtTEohUndHQ6AIXnyNfWSbcTT8dShMEtwYok
flpXdCUN0JDWp+NbReXf2d2t9x56H429EQSNca1plelKaNzXsfPG8as2kZByF6vG
U6yJRxQ5GFLh1+DC+g5KcrNDex1OYDgrbPDcwTjwaLpMrgOcYe7sjX7H55nBCRyN
LDLM25Wa3L5nkajKx+XNLZtAupdR1LQhHjSa8v0oIlmrFIakFpD4ANs8Cm0RW30n
3w738xxcFQ2642jOf+5eITDSVf0gpS4OeCxNXT3fmU06NhEPS8rvVxdvVNxmgNhb
Jdr/Yej57AQQRHc2lSX755/y6F6hLt9kMu933oPV7vEF+UARfXoCq+I/Xl0xdAJ0
yL1mCWKkI8jLDaOOZDDuVSDNLkQVx+oAd93MAfUQpHNtuPTiDyt0ELYs6xFLNVkV
GJd4GGAdTxwrz4S+rkJSlZJswL5OPJDAKofb2RU8K3ZNETPZp0FhFk4ZpCGDpH02
6jpoaU3AsBfWsFw0VQX9Omn0H2If1pcb5GpziHL14xcM8lIYzBDeGfiKtxLRwgzS
GsGOh8L9S1BdgPxzJkdoI215beCHErtEDKpLvJkUIM12aiQyEEyg7lTRLLPYtQUg
0VcKfBUryygGORXccKI1QzdzVbrZWvKXsISIM9sie5IRFhMeJNO3f/2RHpgLFa2a
uZakfrSSeVt2jImSGwNV0W46OCDiyf4Rl1rVoYwnwikGAlhsTXWaXk27oVRz5FJZ
60ls5xko1yXJ9T01mRc7KJN0fOzC0NOPsLC3Z7u4/IbdvLNQ49hIiLTTXd+r3p1d
6+q9u86mRqwIf+KfD6Daeac96tTKc3ehaC4uGfTxsqmMn3E5cEL/7LBfgFXJVwBT
lmYprn17VvC6wspUPT3Lleli9gfn55hO96/RFYswTwQZd7Lrw+KL/ulumuQnT+jG
Imh1OYiO8Ddb7odYy0C7RTdKBfUqnYtdkD+ohkpRko0Wf0B9/yEZroqhROVGKcjC
VeLKqOlYe7Zj9X/pW52Rfhp3Tyd/yvEb9d6qg+7r0sI22RGD28r5QXg8gAmdIUhv
Rbt4dgir5z18YfzHFBZbUfGRxLtK57ihQRkJrQzi4UczVfvJXLCM15COhDjb+DZI
nMtqFE09pIpCqEh2kLh0jNKdBMpnuV2XLL+SJxB9X+C7Pkbp1bqaD0eSRREXXDJV
ef5/vI66RdbaR7CLIFiyv8gEV6i3vITgdGPmw722KWUO+rCIR0syADPZUoUOSfEX
3uOShCrZSRvpWOrXDD4waTIvS8sJXTKLf1ogdPrZd7H99p03dBFH2vuFDdZAQg0D
ql10Dg0UxIe2tbdM6Qrof7b3gfvC8zrbMtEToY4gRD+gAYdPa7njZiKn172jELew
+v68VE5w9Nkw/SxHOXMpoSn+IOWYtJj9o6pUMm5bk5vpuxFtPzkCuC+2Y6VTGwl1
ErKRwpkdVIOEE93ZW6pt33EkEb9VesoMpEHq5wOIgHZPa/x0cB3ErpfricWHykK4
nLLxWYSUrK+41x0nBwbJdrDBxc96okgo91zFDzxHpxLp7+nGkGZPj2QP951K+gRp
Gi2eUKZ7xG9K/Rd0sVKxuYcErAicGW5PizvxB+uOr6b6Zh+R0H6TDQPivnzXninQ
bjSQcZJUw4K4QvUp/OJj2IAmekcowLOfO2VLhuZSLyWMDqMci5eUVVJPU+MHyJpV
3viNT2QWUC/saJ7uzXyg3IHrn1DZaFeLh09UYHiDi4QH6Pv05gRxYNQ0bzjyij2Y
N4n5Qlc7Oeb0NfqZLxJ4dIdNETqSqlXF6FF5YA7v4BSlvpGYrECCnwdjDUq9RTju
wldhyQjhHwNBK9lnWGss5KugIUbkyMcqFDMJ6fBsrS5cramNhEIbG42CiNt3tgL5
DosSJYnV8JAepfwcPpZvwk6udn+R6hukod0/b8Z7qoDl32gAfeO3DcX7+YXGgCf+
2nnCG4w7toVOvfQzZCT7SvuuyuVYRX31NMbwDKjPVWQYuAfod8ZByIhlNjKWqomB
5WM5yNNg1NzahxP0keC8EVk5lzza1ogE0hQdrDFezLohShq4/juMZySndDJtJ85J
Il7RtoikVPeaalyt0wYbEMxIIFYIua6EeG45CBf3uyvkqnFdpicP6CRy9FIX6A1h
krCXghU6vJYPUG1ZN6/79UmovZfcQYuEEIMyQlwx1gjyljZTyAR0g7gIhhyiUtUQ
9WRaAeFvOU1FFfePT/E6VfxAPOb3FNw8qmBvuCIwSWcCIVpazBXzHy/rPrrlylM7
92uvKA5pP5omzqU2g2dx9rkbEa4EM6RNDUayXTq45SBaXeKghcJJbwoC5V/ieint
NPCEwvF4idnO0X8l3vou0dVtg6Z0+R8Y0yDlBLeXG+jqevKKk2mdjQcR1aQTLrCR
TRKoZZyQKroA6UnPpIZcBODzVbwHG3hEFl8hFmpeFThPD/ecl2Zwqzwlar4uKq/i
YsNqVaqs7zwj6p5A5g/wIzofiXXHkYTrD6TP8RL+UwYVPr+O4DreG0FoPUlYLslu
zyXluw3ehTLpUwElYJJGCrCrszTa3dHvuh+8BpnbRQgIZu1EQVz34HHJ0ikmyhpJ
lY61TbpqGws//+95rvCEAEP364tiuJl8MEt4OFmlOc+Qpb1GGsvuBx58CFM53Pjk
bPmW52r7B875t+mVLAYg3M3E/wb3V4RWQUI9Nt0fKJ3RBiqAfZeLOMoLzcYanzHd
+DeLZ/IJfBU5DHCKup1j5ca0HQCV64UD8Ct0dKbFcVDhdYbH/q03zktvsWBaq/6V
ns668L07TzsJvdfPi0NDU25vSTLJO7MOF7h9o3gAmZJOgTe3F24v6g8+rh5selkp
medvIBNiPxjlzPx2j9vZj/zQEHGmoPKYDePehXaphoeMOpE6Shze5QMFbrdkkvTj
wHs7gu3Nam4z9x27ffl/1Ag5ZeHKJMdI6yMXRMPnAlb5lKoJnpbqgkFdsLPc61sP
ThCpAOp5UM2lsc/fFQMO/E16GtJ445WXOtdQxd3RzUOb+f83hMO2T4ZI/chS4elO
Zn3w9qcKuX7LbWpEWIO4nVFWzOfOrXGyVxYwTfXhieRG8az4ezNcpqsPT2h5qJ2V
JtvV/PNTjQ2kysTsPyRcsQhMeqQUKXtc3gisyqH5TYFoo/TIcJWA/KFzzbD0x0tG
AuDcvrxcNOXuyeWOj9cU1UCmuGBUIcC1RFCd2L0ysV13YHWZb2gLAMjDGTMg0A82
AoPVHmkXqNCQxfz4K0+j1QJsDflb18dfdEpDNHuD2NLs9+ho6k6lF2OisU0t/fdi
SQ3Q6v89T4G6aRtx7ywhIxRLlpG9NtNkwOsgNtOMpcSOvsW/Y2io9PBT8SGkS1SI
yyM9SD8pVouS9w3C1ua2HqTjzTdaXwsXWt15Zj6oqCQ51zGDZEVv4VtRCSTd+iYx
CMy07hOEzWPdHFuby6iewLdjOn7dk5/+Qj15ETOZh/n6NOMH5XMlkLnKk0IutOgi
74p1nQIZIJZbORosx1B2PN1iXfhJERLYAHXuPJUjdqmLRoSW7p3ixasBezXQHQPa
Ws1m7HXweIPUAT2NWOTu7i0qGMGhi1R8laMnXBNIWN1xgcj9bSXaxK6IuA1Dqk/5
FWEgZ4knB9E5HEbbyq+zRTAiR7UKtacxs1wmUTsylrfEI3cSm9sZnFd7CdYJEBZK
9Ef6wzmevayvJxH8m4tPaWv68tz/47kyYLXbifaZtKVtMAqSEUrmOPHodPRP2dZ3
WuO7g4BsJdszgqEQk6Ty4xuvndto3aMR7k8s4v+4L4k4JXtwzk9cPZRot5XmDv9i
cswc1LcbIeAk5lXX/SnSmrgFKqCOxLKvb/DS3bTt2gRF9fMpreLF8Wl+J5iA5ef1
XBJfiOg/7uKvTTqNJMNPqg6pqqYekZMw/AyaqNSuBO9RE5X1zploc5KVkAczuKLA
mQRvXkQsC6pI/k15m2XOYTjm+s2f8rP45Bm0ZVIFlLdd7iLfz8sgQGHaq2pVKsWt
eJRsetuwTHfJONPlDAkHocJmyp88NCbMwsG3fL43bYCIs1MWjFPC6+sMwAWEfFIr
tWAqap9C4/J6i/Ei2vWgJNmkIYO1jxav8Iwpr1C3I8QEZjeeBAn0k3CZSTxbYLbb
sxT4MBRKY89EQInzvvO5rzzvxOCSYqL2IDhBWw4scg9xqjxcjnffQ5Q4bPnbRsP0
/6i46kFq4bONb4BgBDn4fMhvWM3KZrb8JX0iEJgcvK0D8GwRjhDhIcEW70keBiOy
bYrdXlyi63XwgpnFgQeu7OoLRWHs8rMArpg0CN6GNK2s9zbTolKLJ5ryr23uOJV3
37Aq6WbSfs2e4Xi5Z1TiIMFijxgtXE+S8Q+1U2M0iTmAXgDaYrY7+eEMpuuz6Pxx
vwZFWjB9yXk/ATrtYVZWUrmws4yzAvyOPIT6Pn0RLR2pV4ipT6y7yISPaLLM5oG8
PlYAyRMZtXgeZp8EIuvRr3rqDySmRzoUpfxsToq8p+bA3IjSgF3G4SbTA7DDrrql
gYziNnBhAyHovp25Qox7qvC2sxYrjH7IxLE8VTU/ZCVDGzXpT828HB2WCuGPRCK1
Tvkm0bH9GCj/DxvXBxLkpS67qjmEr9qthWF7VRWkyJyxWFDLnngJv041MZi6hKVW
oSaXJ6WoAgwytbZvEzbQI6/dRUT6LaNWULEd3Mb045YbmY31MEXS55BI8Mz26EQB
06ni81CTJTS0TxO+VhN5z1mutwlDMkDjSKH7xWWbObShqdmK2H6FdmTyzb8rGc9K
OU9Dv6EFxF5whPdJcjJa0793WPAop/Wio33Rktz3T6btkHPY7sGk2+nYHt98iwYB
aUidfpwHKQ9449eAllAOYzfynqT/QO1l0Iq0VwUuBusw/asJlM7zMLcWleAvKtQM
0t0KRqycCLfPlAss2JtRJf71XKoHwJ5RCjJ02zAOTOQIDFvtywggwCOQXw20iVjp
bDk89dEyY1dQwI+HdcSBBh23BQgsYhIck16y8gDseD24iZKbpwVT453GZP3l0P7Y
rwOOkMEfB/8XZ4i1Ppa1PSNFxumsOa5qDNcQ7k3dgiWODr0fqataQdOuejkwyDEI
fPTNTbSkF7AMTnYXCLzXARJZCoaF9fz6qRs+KDw5bZ6H/+3aEnvcut2CLUQBTklf
0sL6ht+vnKeM3XgB2YEm3HLO6rV/Syd55iL+g6fh6JEwQnf6JBpyySh0bNGP3llX
bRtOnoAo0YKud8uero6MoqLuhSkWozPJSA+8XJqrYompmfQH9bIxVtl9PSCzdHzA
94A1DUxXZszAdfwT6ck33l2W8P+6KYGLaG3j8HxYhKbZfCvEhkVhFTosY8nztGYC
Fn9EdChFUFOSis0S+euXc4gS66DtnyY3MVY4QDiMPxufwILOOggBoBsA0wv53Nzs
Boc4dyGLklVv8F9jxliJAgnDdXjHShpxo/rAWDxrJo71vFR9ukr+7cdOPZjl7QqJ
1gcAYiVrg2InnVVIUZetDz1rwcc5EAPiUH6aQc5bpQmoRYwmNnjFA+t/B5Y/Tu0z
k79Yg3XPHu7gWjeArv1wxtwe0Z7SaRZ6iZRmfAk8msR9ECxWMx5o14PwDtIOkv15
XJwsU+QUHKr2ivm4XrwR5IL8y3GijrQjQLl1TuFSIH77wd4f9sjWKAdnSI8ueCcX
ey0AALIocriMQfXrsF1QJwYvJUs8MfubuRxur4gN9UwzGlzcC4+3BocJh58ux3lV
AxMZXcTOHKUhYhMP30lH1cXVCUONaaQnr9Z9MlpDs4uie8eAoNa/AsyGXA8swndM
8xNRdamy8Z66u2HC5SDxnPvMH6EVE6qK79qjMztBYG00e3c+/r3IWkLqHjQ81s7/
XD/XJKsTNUcXY2hGfWDyjyVYF1Lw6SpegRBmvLY6HBmRqF58NMMxBmST+r3xantM
5myVck5u6h7toUAbvFoEkrV/coDbsb/hGKIhPubTPwa6gRm9oct8ErsA09LCWRwq
XATeJjh8M/+HJZ5aNPXGlH2BBPMmK21hdCVMwE9Hshf7jPUwvI5ea/G9gckwNXOH
W5uzNB12XeXyXQc7LQjUFnD94+/SVkAX+AMv5pauiSC13LG3ayxMRTQDWFh2cNbU
TugTKL78DgndKV7i2l+JgyZfFuo6K2ZgM1aZVR/niaXq7a+apAxJ+l0ybiFJGRNN
qDVj09sVnvFlfcxE8a+NozgKJrPLcuX2aGx1S3rz7Oo33Sz+mRd0435mReZM7KSK
7Z390a0wz5sOPiGx3TKJUu6JZeQlOXiKEtES9dhHrLZyq9rvbe0LJbYGkU/SZA4t
bUk+2W4UWuo1dv0S4mm8FN9FYfdGokBGE8DSp8voWTxCaNY1KINqpbC0kvaY6eCI
2HTj690Z/k47/mIHjqgmaI2euheLBi7SewgxjfaJrFZETadK1p+UGwasPKkqeG+D
5VLKgSQguO8Q831lPqdnOZzx0cql+OAFmE5IgRnWiuRxr1xIN2+Fzwk1LVVVQbed
RPWif9nhIOVPHKQVPWoswwbS9xZOoxRiQt0Kh4OUT12GnV8K1ya6SRqRTy/3EOom
5KmX9LjyX1dOY6VEILVlk0jDllTLCrqU7piBbTUbHZeLlPdZaKhCUod7CWBZwL8a
h4Jsegj0aZ4T8EmML/UjnXw79GRd6rhCwYHR+nnT6yklj0NTSPmSoWDPYQi1GsL9
+pRvc2sPFTn6jKzY0EP7k3LzT+WjrJuNVFzNemrEjksgKdrvmPF3vy7Sl5LZMGoR
poefzSPsuOJGo5Y+6ycJVQQgVOS92NAjXtZv6bqWDIM2QI3QhyYNdWb+gPDx6wOs
Q9xLEvnfcAxQq9cSrqqZJV81VY3HAQfXTiaa2SQCUtbFcfadaHr3YgVe6tHtrFz8
WWrYvo/MFb3EfuiXvkVpi9YmfhX6qkISSmjLri4ttv2htR8QjcWMajmHosDlZUwC
6UQYr6yocU7ZORtUGwOtm5WeowI5VVct6x36RbmUfE2O6Kb5nq5+xDyc9qwytW/b
GvM//QDz1Qa2sIWOFyUctihyacakzWgvnr+C3leFsE3XChERA06MSI044pFHFlHq
LUBlKanodcOHF+UpGWTkrFyOtIUv68g9R8uamhVGVSVQTl17o2hyXklYKphcj/Pv
mcgJ67T4IN1be+emKGsOaKPGhlLc7+c6u2Jwtl1IrpD4A0gNpLXEQZ1T5yMrKun0
JeFgReiNGEhQ9V5bwuP2OInkN4gMOBMKxTAp7G6lp5vXpsTiRI2/w9+7xgVOadsp
HVklQEqAZIbBKUyb/z6ctJsznBAdVO1o+I66hA/9PRUSF2oHrOT1zSGmtr9oyqN9
cv4v88N8zLvmy8ljkqCdRG//Z5rz7fYkBTQfqWDwd9RUwFBVBrwvySxFXhJtPuLM
rBa9YgKA1NJTGoWojEwe22Sg3zUW65mK9kCk2Gj7v73Ih/eO667RlhOyfI45/pv3
Xwcq/XHf0YZwPBr7u2a4w3KYiYsOjbwJC8KeTb2u6erNtbWatFRAHDesLvaXeAM5
xhSKPWm153IDB3MvM+ovEsw0HSR6chVKmJQwrlMINYkW0kFRfk4CCaWAmqS6O2V7
Yghy+M0QUis1bTn35j6caD3EEO5UascxiN48bno/e1qWgq+D/k2aTUKfxsxaP0l7
VW2w/+aOpcI7+XZHegQBjA+a6DKTz1vAd5oJ+TPLjbQ84VUczUMYvQnk3TARgmxk
TDIcTWcTl9bFqkuvpxTVBj1DfXoxodj6U/uBeztOntASMrgEK1pe6f5rXPOMDR73
gMIbL78jt5SnJ7eVxTpDL4KoUawDIuh1bw9T50M9CINweubkRtg6ND5SNEwbs+tS
Mx6LcRg3tPPp38L8sOV6rX8WQdAQ78RLTDnhiByaJJ2rBVhxTFEcUnJRwEOmrZyn
BEWnBzl1ObkXjMcT/n4XPmzTJfTm8wHFbuu8UMYQkj4SuxhC06cEQhPDuy9qEuuz
LrDeWkvCJrMDXu2zVAwp2ImpvKU2zHpqokAE2N+Jpmgl3bF8hUaCoI0ipwLydQUR
liVCuNN80/AytO6Al2AmNxUOVVwEcKelZ5f0b36ZRWwWh7xLpXzJR9AtGvjSds/R
S4ia2oqwQAnXnytvNoa1/UM75fGWWnKn4HnD1s86wD84MbLHPln+OYy8SvYNO9N/
TJPEFAwQbLs+0vOTM3WwqfgIItyVHwspCVM5cdxQ15+TRuRbM50KIvqZfm4RZm+G
3j8yVnsZWGN/qM3EAUvo3QL2H+BiRrDe4iYdQMkONmqxDgVL31JKaYNcHhUysy6H
mQmZdq3kZn+LBf/Kbl/JcHo7anX/3GwKBjSDxFtuPQ28laMUske/EQKRW0LUcz2p
5mVXu7JnwmLWZzISxBj7fUztzQHkt+95KC4P5T3x33wKhDjlnjV5WvcY5q9/kC2u
NhG6b42nXKm8EStwEX4Q60c5PFXHWtfy4u5aVH4e4gQsGT5avGYgsdF/HoHKccrX
kBEAdj3uTBOxjweDCykjb2ITNYp3TIAJhC3GfLeTA+d6ml9wx52nIKJgyI3fYG7U
EjJeo28/torCBDpelXfBQ1YWcFbRJqG+yvLa5LBqUu5rrIwpBvDvt8luL6zKM+pd
VnD7wf5ENeBUFw31u8zHn+bS9Xa3HuU40gP6nA+oetuNdtEmDkw87Am8Ash92XfL
0uY0anUta4V9/q9MZmDMQMclIXElUECbiCgUS4ss2xbZSDHY6HWpSIsfNVE8B4SB
93rD1g6VEI4gE8iI59X28185/gh926lxdgEtIwTdJfhjmrRI9qqFHfF4ESzHao8L
FNXhMRqqmuok5XDWFebrbo207nfUaC6R+Y9AVkCbuEfQV4OsbcXrgvyZEGon9bGU
z13KQiyarVJnMbF9y2WBcjefjhxHE2RFJKap1rML2VC2h9rho3ckAfHiXcnhk5mr
2NMn+2n/hYRLgJYJ8Qo+TPmvkvj+NmMlvGm3GKqEawlOQGB59JLinGz6irrDyYQ+
JvkyXYGn85ZigQUolIT39Ggbc/WhrdTvWVFoV00A1gOd+7o3Yn+nUB36NAvggDlV
r1FqaBQbHewI+7GdJ/5kFXw8VBaOAvW8V7t7KTlvnXfWzb35raYSMjKVBfHAe0Wm
tLh34BEG1jk9xx2x8VESeH+yMFUtA3q1g3Rbpza3wDptoXjsRq7ajiQNZsaWUoJ1
2Q7sFRBV03+ZuFgEddDDJv2mdZ3AHJz9qSoPi3j86ghuh2qunOL7mggYvt5XVjlY
KdUNg20FBR4NF9G4qS+k89Ul6wq8vb8upFnDQ6eeeMZAp5O5+bVRlFGaF9V4vz8h
n4amAu+yysdPsySgMymKhResDuY9JWffpRh0vTsd4gDA/p4fxveSwRavP/HqDZ5Q
wCc4nTawp4b4r6LVNSVqSELv27i4NqjSmuChBeFmYEdNVRFMvqgBeBVnxg12ij7l
hXiJVWhhByFjc3z+jBrs+Cuicbm+MGTx781ZAEEMQedkZ+NLStO+YOudOC+PqwaU
WAUf+oulqrkEoQTG5BCASxehP2cFjHFYQ3zGBdd0o8bAd/8eF5h61RTZbjeyzP3Y
6Dqu+0lBup2fyiX0mFpWDvjKZzMkLgNKxF0XteJ526hLwfClh1MGX4cyWt0QJzz9
E4sjBcJd/Iflp2/kVxcY5wJ6oFVdy0ZhAuXNYN5yxK3dA+aQTYkJMK1R2/TahwU5
0Ru2sCMj1S0d2n4ZCvFOa1YhgmL0wm20u4IHg8No2GoIXz/JCfGE0lKeB1xgXerE
lH95R+cjQWE1RFcVOLPpq8MIep8CQfD8WNvP/xt1HNANyw7+TYU5tbJO8KbaLZ+X
BLkSG1izQZvRTglOXItwH1sfGt8nmb6PEeKh7VZoTjRW7EC8/OQIMCM+L52vF5V3
Xa7ixKXYX/tbCFy/iV0PA8GXJVJj6i6fjFamUFup8If52E3Jkh3EY+bXV2MTgSYg
o37xZryZrOEGUG47SBMXOYxbmnwzJvseNn07lyB/uBms8YHIaJc0OOGt8sKbzan/
DOnxEq7JA7qJPwXlr514TpE2Cq6SFK1YcOS+QlFniuRxdyJMZKCKFAu/SecPUbxO
/nr7tBAQ1cP/+bmu3sARNXeO+HQ7uivPJIDUiGaGeMql5EhOML61d4G9fPY3bGgJ
Yhg8wAtuqAFZXqT74A/8xSK9W2i4Sl5Z1asuAxW2fagr7b/3V/MIUleQ8mcP9eUn
vUmLlICMt+hTJWC5Zca6NKVoBogCtMWRO6uKRoQxFIQ93h5Lxh6nvWTVK/c97eLR
xTHshUAfUdS/MnPUOIYrmQIAGzq7p6YCbE8k2Qy/T24srpRFZ5ZsZqST0CrAenOB
y5FmXLozhK30PxQTZbZwpyYD4yP6r1zuFMaFOyq3lCRQTnrPhma68WdSn6MI7SES
JW6+Q9Szun6q0h2SfGrjxlX0VkCxw3fbSbMzMLGjdzMdXmCiF49CiGBZxjmQHlJB
hAKgYmdSN197HQayO6PNe+G7FR0AigpOvY/wiB2E90CbHxO3d2mBnXHN6L7070tn
jx7jTCkUjAaa67s4VjXpn5D64WBfp6kGM1jQ9XSkukAM5PlzEz3n9JvNiHN9xe9O
ZvyvDIOMsOfZbZcRiVyE9UOBQP3qQG4y2atTqSDq6RTDoJ0T3LjvUN5gXwgTaqfv
lH46E4IRcKpkh5w16P6VhNkTOmhb66z07AwPq99rd2s20zD8BoHpsHLNPC3OyBhQ
FqxvOWHsMtUplTYdGfEALCgVP3KsbbQANzDk+giamWHdekGBpa4r6TnWIL9GR7RW
Wb5SMgjWion9yJpv2DEOttD5wCxfgPndtXMDbDQlVkAtrZ3t7gUqsroIGvoOadEH
1mTaZWs6exhQfkgMY2QiJljHk5tH2+L9fwBt94j2N4X4d/wi0QyE+oq/s1Lm8ybH
/Cl8DNdrnlNKX6ojfVwUE8rU9QzbQrGUHyIe1nzvfCBqhaAf05xxAcbyMJS7I8Bm
GbdkbTThPwSjbzW/xu6pcA2BalzICPlgkNgmEcGu4K0xXdH6hbgtrsIhPKkKk0zI
roLFJd+cGkEGpsW+92/6NvucSt10yZ72EuI4ChvN8ABN4wAyISc9suQFNZTwgyzD
aoOz7cW6QhE1mbj5hpmivJ9KTL7Wc9jTaZYwQWstr1azGqg6C0w6BwsbwwFvvN8N
VhDNGCwsfSFk0GQ3g9gIRSdxZiAOkw7wfV85dudK+HejkXqv8gFDLuCm6bGxsNwi
PcnQQbNKrLiha+pKkJDiGpg9Z7mh3unhYYbYU2uCL6eAfMN6XQOzAqGXN+vfenqu
zlD+3GYBZlLJxIZj+XdeK+Hv7QvWI4SofGBqJjdChdZ8q/2/4lNRqo5479ZNL5Hy
wcW99eUvmAcS8FfjV/4/Zz6+Qv8EqDA0RsEw28kgrLBUTjGSmODZXoEBkoa4mizU
aEYvs1hkf95f7G2zcACQtbStoimolgwsD+ZSFfkSEWHXao77Fk+9JB3HQETU7FNl
yq3G/oHmiSbBGNV43C6Qdwk6FweSfwZsdJQuWvvcFx+N2j8INB9HsZEiTSqEY7TT
o2FvCusyBoHOkaS76et1lrepUWuBRMd3+XqREAZAfSAm2Q8eeCfVH0pXgbrNx/rV
g1sr5EgX5iMqKFizgqWBZJUTrAG5NWRWp3h6g1ebpsI8YLmoFOsz4U+Om6OGvkSl
MfS1v72fBg5j7hzYYYpS/YDQIku0PljMpZYgpa+iIFAZZeS5ZsBI79eFPlp27aPU
6YjuRUGXUULK4Dy3zSVhTBryx2QiRkokEjG+fYy3rABhJbsD6RhDpvhVzxfpJ0rK
DM6E+7cxJz2qo8R8AxIPaZ/Kl/qCnkSEM+U3PgZluA1HKbYIbX10q+WqsqI7eWkD
Fnm06ubRS1UcgKX3mZdrbBLgPv3Y5MuGaaND0KoVTeUDmBvFoTc/LSco0o5HYPNz
+bp8itmJ3y1h5NEomp7ajesgJo9HagG80YBEtk5TfXBjrU7Av/RHuhceXke+ij1t
rvj9zZXgl2VdlWk9zmyVVg/hQGcZHJgv9XqiDois3u67SqFjXsqs/ED+RVPY9JZN
H6zj+cyNJtV9qJljTyVvtF7RdxP2h+9k4EAOR9YHA2rwMgCa3MemzQU8SyueIEFh
1GMUgd9qjZsM4i0lSpCqr+adW3SrR+ZBIGLx918Gw6qCvaKVuleetSLJwU1tK896
VtX/YuUGazk9W6c/tYcmoShWGKPanwIc1Kr5dEOS6XQ3ybar852OYMDnXF37DHBO
gl40wx/pmqer86McaJbkG2GtpU44zoNU65Qor+tTKGZHALbIZDOFCUwsMXhLNcbU
9qJzr6Hby3w3GS5kehrFQzPNZaIk11A8PGC1uPsVpcGTvCLwlzz8yhSZn3G9xorl
5Hp7fBCl5dxpMp3hvsjdo0MBVpz4xy3PtA/bGIa0MW3c7luzXTsRX3abbMPchFOI
+RjxG6AlkBZ2Us2+dELwOICAyPU5AHjXUQ5rLD6R8cLzZW2Tad3TPCyOPnovCm0N
fXIFp73sUPDHiRNtkW75TRagqfpjXCsECmLweVAK2SrACtb7Kry6VV8xqKqO7zP4
d251xPVlU9sdAnhEJNJ3Jkj1WjUe9ONZEpDt38cW5/2htvsIdq3+jZvMmSdNzRQy
de4fWHUwjhVEiTPapV/Z7EThF3o1NXd0gcUYSscX489GtYLrP0gYCFzFjCj3GejL
I4hgDWT23HJI4Y0vVNaNcuRdKqhoQNHoQS2sKb1GjO/00GKYlZ5eBgMazHKNnJMd
gVCujBW0QDmnDxLw5YLK9p9IlwrXX59aQm5eOjUCOoE9nf2dem/wUui3yx+0PlT2
UvdH0sjT4pw7/+ku7+7ShOTisVp8zlJVwz4vk3PHUz1Vlm+yHEsXYyrE7W20HPEo
1atfvbsmga11oDCQo0XFdqeF2QcvCO7PPvFvLvo/SYAYzqs+02rmAOcQB8fx7t5W
1zN9PehTCPu03d919bDZhxa0bOAAMhlWrwUlFztDMzEbSejOnvtot470T5U+uIug
52lOi2H5mBzglL6XEx5FdTaaTRIGL5xofkaSXn3Uwcch31CFsCotFZpR7bF8R+4N
aKmdCMIJ6nCl090i6vCMKGuyUopkvJTEIyEmZnTQWdSdOksPDXVmvcewym0h+ToW
S2qsqeXCnkiYBZVM7YiV8GgWRCItK70XMKbiZ5mk7PVCTExE2+SEYn6NDKbLVk5r
FP4PHE15IIBzL18H5SCM6W0ee3tPwKjWeqkKHt7TROwltypgjJ9mRoHMPOYkskSJ
M+H+uLOU2UxMH6e6jubZCzplYgHQDzqHJ9NaTqNXZIW3d+SImmCAEBC+hU1S/jKR
CJtNDg43gcpj6iCf5N9SQ0zJGPJ+4SQSoo0AyFlWRxDGvgZv1jq0h6yR/t9sbH60
ItonPSmmdDlsf6gn3937HDlMX7npc0w3hdGR2FQCN47O01CNkokBs5WoTIcGJdKC
3HRsjT3+tgPUFXJEPXhqkySIM4+EprB/+QIfXtDZtvRvw6dmgKMznJ5ziQ/7pg6a
IpazC5V67wWljZhWLUbhRoR/WnQPrtgiGNz4nCQAIE02BJXNHUKW3+WwctLXxqUL
rWLMLd6ueLwjQrBhUwUDL3JW1b0JLnas0VX7WZ6i4ENA/FuqHZElO6ZHU+7iiFEA
qj3FDwwmR//yY2eCjHYLW1U6db262FIHU/5LhQME1tW0uYwjAngPOg/7CuJnGwOo
PYe2hJ2OxPXfQjSzlgEPS3JE3icnvOKq7RBVLebTauVa2sX7UQK/57JBR29zPJVZ
DHSa6SnaQeGuW0aVPWk1NYqs/uMWdfORypw0o9m+aCremmRJSgz1Sis1hA+j9AFJ
1/SSMUgenprY1g4FX+DS3RxphIvK9+FCGgAIEnUwLsA1XBwqkM44id3Ic/i2r5E1
dE3L2bB4fTEn2RxIFuMnuH8/irmUZiZHa1IHXSvRtt3wdXrh99sQ/zyL6dVRU/tZ
cf497XO3iGmO3WlWtAsL3ZKlR882FRwoGWeAMlhGx9ihBhHG02KUNfC7bzqU2LNH
4mW6tyKUCF6TSEKsh7zQLPM6hyzuSuxwjFiMOH+8rWVHejRDG3XE8ucZzveWZGZa
66WDL3E6ROt0qTLYTgZcCu8pqZ++fPYm3C8/NdFKeRkCW+HLGobsqIk4CN1Dixjj
ACjXzIQzNqQR0T2PljZ8ZeATv1JJQ9tfa7nKSvkkZkxJosiSkSl5NwtLDcJctQWq
TCZ869TGLXrMVnD/zR+2Mae7CJrQBgoX2gQhtU+3ba3y77QAZYWroSHDzPX3J1zV
dSoG9/5OtaK9NmiWZRa0iZ5FuWyBCn4NeLx8RPCqbBtf3Fw9kwnQpjZbSfKlv3Zl
mygEhH32qypEjUTtKVfqhw/ZcmCxmfeXSuYhhZLJN04YkW2e3RQuuIdeHxrN0c1r
G9dsxggfCk/w+1TdQezcuchZFkPPzZg1vZhOtur+eB6CQz4RMi+yRWDtcptrSQ6D
cQI3jUuDokO8FCqZCRCrMEnzj9HESpXJ7JtrUg+/OmyOcBvrs6qdQdNS5NNti8OI
8iD2BLSCSg0xGq5FNjvAwypNsLCNlpa3G9niIDQunCHMImSU5vHTCWZ8/0pVNVyd
BFHC09+7xavVlLfmkUX//EgYE378bPq8s5wH1HQe8vC2JdO7lXQy9rJQhhjildIC
LNIPm9zoZdjpchZP7iNV4WJPCD2k4JgUfgXwINgypthO25IvXsWvOPUdWowYAg79
t0beSvhiVco37d6aSHK+HYvQT5XFN0EKXiNPc1pzRUBg5RfVpbMQsMCOTkjl5n7e
Vxxc5ttldOCWJ6N/nUG0lJkE8R1GXnnZVw0SXoY+8V3okkSUHdZ+QnhRnz9CXpnj
r+7ZOkFq0blBgceABO4GCXjl3Pur9Q8k9JGx1rQOX2alyFgqVaPwJcWSEt8PLoJg
vSaUHl/HZHsurSxfClU3BXtxS4kEEX5Pwge2fUbrcvKq/XCbyT2iFlMlasrVFqwL
VmzBtXR2wi8SUUGtWSgwb2Wvn/imTmfYlkCXRaCvmRaZmzuApgrudlT9qcMcSYUh
yyLhCOajDBjOzXbzkX4ShRIRtbLNdS/dxN4skw7A8sZhqJGKdO1cLF31+R+tJbV7
qUKgdq+QOy+0HhuHCZuqsKMJJxT7Sg1k1444gFEJ2GvHKZ++VH7pzDiaQ5RYQnRs
0Z1o12BovltCTSZ96wGd3euA4dIcX9RP2UJi7UMkGRFGnB8cHHOWrJroXnXkNlsV
+C0PuerYan7SROT9I/VEIZMgnKfyAyD7gkK7JHbbyFlf3RywqxGCTNSlASjWaTZt
t87U3y6sJtnYGu6vecKg6VQa+1dssOtCnhYdoe6FBUHELW8wQsZS8/yBMjz/zGV+
XzVlloa0aGHkynjbpuhRHI7YgtBaXzx+7ZlT3gzPnGoMYHodIkKlQt1zEygrZOo3
qkPSqfTgWnk6XOXzKAIjiMRXERUNDcSLsA5MIxHQBnkvOXGr9EW2ttkMoB+Zub4p
WuUw8BrJa1zW6j/WpLDIuhbbi+2K1BlDhLkAKkYunb/iWNvZRh7ROlh2cs2gZYhA
grBcSnsUsk3i7kgvOODOIFg3mE7lZkSbhxrBnOSX1NrdXYX6Agn4CjCwkzOC7OyR
5V88nCbc/j2OqabORFsI2CqO4cvW+mr4CsmXf8B7DrmfkMwQS0Z98pFmp0lHoTtY
y+4SEaJCU9+imAo+2Ux6lOgcTGRiXvculUlVwgNTNaNnzi4Wx2QLJr9I0eqrmJyv
CT7ptTaCtS7XKZnPNVtWAfjz08a4KDfl2+p+3ZqeVQoWWk6YD82SvF8uveY18Xac
3Lw1z8BURSIYtTug5GzE88ZyGQTtNMMPwdbQE9G5/Ni81tkBvCuRkfydoqBV/CBw
cdlJNezmBgn1c4jSIngCBn4H99jVCbV+GeRXP0cMif9PiwDAASVd6qbgS5TrQcU8
GTsXaACQiLLPPHpOHP2gSnuuorwaqx64tejvqQmzLZduFAAOdjYpP2tc9ekdwtMB
VmQaB+C+qUqtXmfovDZ1kKfvcr4gEcztMRp+7IyzEr9U/vyJt/dbRUJjct/wWZOM
MwHEXaocR2YZB6cGQV7Q5qTvn6b9bzAxHZ1PZLDDbzBTLo5/EH3gNSEb/ESUUpUP
xEciI0AGzcD8VIVAmjntLV4RhGDtCEevZYOjoobfBjG332idLKb2mrBGJkLKqIAQ
gH79WyBP1qXhs+/ywNK5TQlWmZEWFPief23SqKjr43heM5SXOBNuVif/B14qscCa
5nSkACFtdrwCKjyeM8c07RvSmSF8hiKre0DH05ep2vtijTIwK3WloHkzL+9/kmAG
C3iFwHe8HuZpPbZwfRY7RA75APvuBJo20ojrmYdPTnTyJynYih7g5V0Hdvti8bmj
x1zdPLuL5j7D2YcBMhpwKgTHUw0dm06NkPCKP6Fb8dzUV4Mm00CE/cPn9a/Ca7K6
0FzIqMyQXGBbPn2aaLTar5Z5fEH4w3Q0+jUtq/CN3C+tUx5ize5Wi6n4GR30dYuA
5EHyupT/coAmHnsAuryJDZ+OJ3HqeTcBf1ZhGPcOGBGq4LnnIPK/iB0fHv+Zxxrl
53yduB1NEqcg4VX0oOxRRDOkua6qdIpAGzfTx+0j/f+dO/uYFBZDb6OD5/wWhvT6
MAAtTfDnlvZ8cpy9qe1uxEjF+HmTYVqX8F7t/eVttfVEiIDw1Q/U6RDeXH7KCNjD
ZIa20DNQlnRb5vRcMq2h1mOk1245tdOchE2juAKPIhW8ef+ugoaj9R9cugK0FqJN
LuUXXJ/70mOUygqT9XDlETqSksSJYRcx5ckfD4QFNbw3wXy24RV0gcNGXjxhzbN0
M31CdxvspcabPSBXbyRioyEHIfQlcnX/7cGVtwZi2C6tmWRbwO9kNXgtU2vJpu5b
BYRCVfF0nIpqQNpcEazJfLORAkLd7RnVqYNUMZeGip9W5iTRsFEmK28D1jKuubyN
Sjf8pozK/gVV9uM5EVEzvQVPrs1F+PRBVvoHdeg+Ltlac9Ody8Z4TcQRCHYxP1Oj
JyGjEQ4zAWDCvvdLDkpvMJLFRBLLdctrneUOcQ2PEebQL5gNNKCSlXCmDAQUHu+p
aM7MLBTehZQKTWpP7NinhoqNBvk1zuf/MQ7DSMUwFE9V3nu1kEHU2tJOz0QaLmr3
hqWBaF3ZRwmjNQ1Q6OfBy8UcET5axrpyPhp8Z+xL5V4JTuJQjHfpMU48Rlgn/7CP
UTtqFljR0GQs4tWAHiqiWt5Z83w4mWunHaHCsE0fNs51LnVJZpsUVgsOAfVTq1Cx
rZqqHHYaEwNy4VUYEz1jUOjHyPCgZGuuWfZLmF3uaqENImep4UiUPUEhQhcJlSlI
F3zhiaNU41t6V5zOXwbeAUEUmhZkhPkzeIr+F/OZ31z4U6UuYbGU1XiYTBxBfai5
TQhJfl0gG/6z28A+MN7x+4ODRIF9UqrNzim1xmZAGVipwFp80eQIELrHEH4FlJZM
EwtiFOHrDvFh23r2m8Od2OLKcrYnVe/SmwdcHULehedgS/51Bz4Y/ufV33t1iaOs
Aw5rZgIct+6n3KxBc6VVKn7un2Kw31RwxvOTsBTGTcwalH+YrkA4+fCyt6AyxqMC
H2KxfzS54kNXjuNQZtm91hVMKazeBOPD7Y8jF6l/IyHAXM7ooBQ15LtCxGsthKRK
U4mcTcIXsQQeBMGya8CnXpWZsG6mvVhA/x3BiU+ma7Dlvrl2Vl2VvHffvdPcCA/n
26Sf0sNlO7TSq0nXN0AzgqRgonc/lsPb0HYTlipnYZazj85xCOPRNEaJJ11TOhJ7
ZXJ/g4L6ZECae3nFV9M7yJ71CJuADAv9EV6AJ/dcNRkgMVhtg2W7l5WysQPnrRtt
Z2gClaXkG6ltzvYPPaHK9s8BtdbV6j4g4YJ2w8x8CEhlzxfUZRTyTeewS/Hxe0R2
7gY9dIBb/3782A5QjAhRef9jZucWMmB4tV3ZDAu0Jlu0uDPsJ/OW0AnM7FUlYkJE
JWjpsW03ZY+gYA7tMliSK2a0mmGqo2ghXCsRdbZG2sqdWojZlUl5mWkWxm+MKWeu
8Z2A5fMRcCtpVUscGRqrJjPUiN58LRRc7vKRF1GWdTv4oHSZPjUsnjwv2zVBjW6O
gm2j/U21y3WBm3UXA7Siqc9IBtWHHgB3Cf+hq28ky1kYo+qluz/axkZHhdBQqMMA
bdtGtv2oxmVnEhB7q6Y4yt7mQYoCvj4ntR2KfSww52pVWz7z0EuqvRkb+eu9mfkw
wh2qBgoRPtTTUcgSKNqGL7tlTJxzGp6NpUwnWOKw5WooJHbAXbYQ7OZQy6E4xjfF
pLak/yXRw8i/vwGz2zdjZUyk53pogshN3DZR46C047k5yXg7eOfTIHTeq/pgpq4P
nTyyFUPxbHqqVnLK1/hpm1t3HVQHDJ0bllRF2O9ZfzDnmPYTDzwnEw9bCzZd/+8m
khvxXviu18Sc7CMmXk+POU/94BcrzSaZBrbX+h9gGDr42OzoH47Ao5UjRbDPSO4m
jNjxCsl5rHDJ7SLZNIUMsPqWqGqccyRYLBPeoffERYQZZSt3OpNaxX3rYJQVcZB1
GN6VD0wHNINr92mqH/fJ4DKDnFKZrmvgpnVhUNjmffUJuzSTyjOY3ZUdOvPKWRrD
S8QEwcqltF3KSxfOk2ZmuDyKN1iCuSWGKPFvAy36KK15yRwYLl0RR7bEtD9JduTp
uGeH96Ur7lPdehVlVJNgObecUrXanA9x0vJtbsvf/ErNlRLenTT65GQMI/9uq5TJ
dL6OBttHRdrt402RmMI3UuEydYsrUFzIBuI4msudMCEaVLo13LbkDIDBm+5NGxU6
C89y3tO85km5ULynfnyA+ZVFs9A+104tZs2qglU0UolY6C7dSuza1IXPVH/HBP5j
db9rr/3dZPtkNjo84WWoxAMJCENcCosslmv/MgkWtAbbIjyZg/IwsQBQZ9HCuHzv
HLVXGUmeLCq9mgykPIWq/7Ba3TtERG0KYxWTfY2gDC1pOolvrKh+MFfwdOxWn3Zh
k6oAio5QJz3hlj08gCsrQ6VzwRzWUircDbn3mXejG2mkpyS2BWflq/McR2b+U38G
plu7kQY/d4EMHLcwzTFAq1UM9/fw/Wk9lJm/uM8nVQfuLaoRnb/4HpCbZHCkSCxW
+HxnQQXoytXJ1CMzg9rkYKxS1cCf+TbpH8uIdxhDi/aeNKhETGu45Lrlh8qJx2Oj
sCPIezkXZV+5eDO7nw1aq95y/Vrzl4JdTk+KPcNgkvyzjdU9dcl3Sbb/O0WxQ+ZN
cC2HrKxRqqBo8U00jxauFEpGhuerLBfQ+I3piWATj1iDz9EbpGkyoYdZkwvdSqL+
UsP91iQrbDLx744277lmkQ92Hltd0L/UrsY/nlW9IXGZT+t+Dnz9xNvVOu02DEJ1
j7fzy9g/W6HUBLG+3x3+89WMR7uYGUyUjHDB7P7pFtUR2dV1E/pZve8B4Pr2cYbX
Jmy0er60BAbrGvN65/NhYvB5HcYeEI1EEtu48Kpk+Tg/Ds1op2TjZQMMdmI6PKaq
nbZvfX171lbbZMmAZsgKrlu507z2L5wxLmLpAEg1jdaEOp3RBynWKa+eFvYe3ffe
G0hCJRsAwnMR89PBEPiqUjAZtpm9n954PGITlzdp5uyqEMrqiEJ1nBNQhoqwQt5x
j9uRoto3egd4Z+gp7IhzbEis+v9Cv5gUtMTWP0hsstOedMNZfL/tJ/EiA9awAluJ
7wfkg8HqFSaXnDWvDKyUVHdZ4A29HGXSbr97AJu0WeNTFa2N+2Cbh+/MPv20YqMV
eSfaWrhykdrfjoRry8jeiUeoqK1eZzQD15gGinbSVAo5mC1Nawc92neVxcaViaJl
G3jKFb+lF/4dgGIJ/fI3ctmnog4u9AlQZla6sACS9jxNnitSx13XNRKaUGG5EM32
5nr5h2hiLAlojnJwHG9GsFbiytPuNDCIvoq15QjPClSI1Dw+Ac4C96Bfta5QsgnT
P2FhoYvqrguLd3XO0QqhGyaKcplwVIwBN3WskZ0U2tGZVKmIaU9j6CNf1vSuhj/F
nCEvG+8psrHSZhHa5hpH8KA9QHffEm4CYZievqC3RhKD1QZqjAGzfXYwOhrwhaN3
IG5nqz3ATWMaCpAxF20KTX8/w+8a7nbDfHXkR3ZFIYKybMhVuvejkuK2+jFQ4Raq
wTB1mdXlNcpFDRHBTSU4hWn/QOoKFRUapxB2qMFkdXaEJYe66luqbTnJ39KG8C6x
0PgSXFX99XAjd/Uh3h4zEMpnUKwTGBmlCOkie44/3qmajxnPTzmmly2cWFwBpwMZ
h7/Exa4MOgVOoSxwbo14Cte2q4j1iDw7gLrYRlpmRGpRXdrSQwuoptfjHcPdWkiP
ZKVIgK8oFHZ0SIuPXq1CUTo5qrrv/6YYIa0jYrlhW/YIBemQnwCM6aYABij8syeo
lBusKVZZfsIBvGkiGZhdf7eDDjZU+dZoy0SLWNpoU/mthe9p8IRrB2KDDu5TrkL+
VRQ9z6+XjCWyfMDPAjVTi4dGkxXi3IR9bSbCM30cajzHos/JewMM7rRda46j4Gt8
9X3/1FQfZYYJ4ywcsmCKNn7faMmnoSxIZ4rbLSlC59KPssFQmLWCIN1LIU0RBt6v
KwtSB9A3cCqRPfNqGKwBhvB83OotNskPVjKNzsabYQomxHXv7Oo8d5GPs5K8d0Pn
4e00BH1ccBDnXpfipLN76To5i7SSln0hx9HA/Ep8Qpvg9z+559/fv4gTpJAJaUqn
OH/0BY+537zR7++XVngYdcdO22etan/yYSzYbCb28HNQrlDTM5BAajXec+cpkf0q
iNN5j9tMv2NJcKeNET+10PDzKDtN1mYPL6UTpNDlkxqSL7/xm5A8zHIBvk7YSttt
L/agWdzv2k62xBTfE2AXaI303UcQvW0VVH2kt9WubfJty69MemVqu38J4UPgHANh
5j4Xwj2n71LM6/sdK+TxtAVssYJSxLTfyDSFQ9VFUUv+xCm/dEiImlWec2pIqJkK
94m+N9ElmZnOLGKIatM7EmCNlZi7jSmNQgXdyyToevQUrd1E0gefM1rtJ41cepHM
WKL8di+OovCfpGMyo0zWnqMukqPi7+rDPHMnLPVnZE+H/T2CwqYi+oB9TZdhzaL8
9iIBgqPTNRhAzpwKnAT7l8Rkj78CVC8dsM46IJhrmkW29jkBCDWk0XMNindpSdSp
UJaLyVfJ6xxzLERhKGTsPDqvoapTL0Eupn+gbIlmJZhZjfCzhQO3p7xH1PLEFcb0
8CXXIT23xh9UqIJdO1CabT9fDw36YjqXMSdQPwPJmVWsj4j8WbcOx9EmzoXld89I
h0Ze0C9WYqVKSEWndtCYUsWKALR5WEDwbjRnn4/IW0uifgGWigX0xfcN178+SqiK
nAIPbAC7F/EHXdr5UvmvXnVDcfJYM9+1bWMvZgjcEFVSmqsiBozC2zzWiZNoUHV9
sgbjNjWIzf6jw7ea8uNhAHLbLW+ghfaI9FFlhU3YrAUEFteU01RaXCKgiXk2A07r
L2jl0EPL5N47rl8AuK2zi1g4MCRXBxPfkrjR7zt0eOYJKqhgCEpYxh5qBeYSY8+5
nzXYEhH6p2GxLiBrOkJRt4K5JGR2+0BQx9GFuwpqj2HqFRHoHW8Xj35gyNlcjhP1
gud6mYP18oWOYvbwAwnUQXkDKLEPnuDf+ZZ+iYaOGoTpgAHa4VAngO2crIbFh8RS
nzCTizUjDO6CeM4J1LGoh9Wf3KP/6spXTkvMfw42wGIq+2Y4lynsUYekZgZnyBIj
6f0hVCLMwkytdoeCJQDHCm9HVO2d/emAVCROIAfR3G61StTBQIb8mGiGUEJ5PQAi
7KHUDD3qKEes8HZqbwu4VElOiJjRxxpcPfmT8Kfn0T2N3rDWcSEcCxaBT/wMx5vb
RZJR+6dshO6v5Ua2fxXSE6zYINjjlecgDJ0cr995ztqJDV3JgUdnuZ+vSsKQPz4z
7sKVAB5owSgGrarQqVSfwtwWQYYpOfpQpD449zCdctEoo152/J3pjJZjt9CXeN30
XejFK7Q40USj4YMlrtb1GaNal2fNP0xpfIadT70XwlagzYGoYHCl6KecBlhXV9hH
X6KsdewjY6s16EQLBSoZ3VFHr2ITftvq8CR8q12xk/nfC4EoQGiEsmJP7qX4wy8Q
vjpvIRG0ZUmKO+R7EQChLR3Ju65Qftn98t6Or7vaNNf3+qwL/GNYt+XhLdmAEw3F
ZsX+L6QydQvOY8CBdf8QjXgdPh8HYvjCfKc04i+EGj+w2sDvpKyx+88NI+Wy3bwH
NuadW3jfjRrw67BsBzFnpjyCdfG9y0M1w5ohpo0UWteki3LH/ODAyfecUA/bFQtN
mxlpaOtOQVDRzTjk+MQq9xUI9l+R+UlrI9ZXdHBMIFlNCGOfyqEijvAkyXA4P9xd
y+21Kav6+ol37VMga53SqB2hGdinmVCdHnHJsGMWDg/uz783Ab25IGxIZStb1XHJ
CfrS8r4pEhw+sZ8LwYTQgfru2YKFoDYvcsufKz3sRjQIwGXDfsWxgO8mEVdS6tVd
+QPJnVD7DnyiXawgVKm27ZLTdvtZeXcpjZJQ+A3mdYWLwCMlI/QQwuvW/UzBxE23
qtQydxFXVohlgGnzNYmHyUzbGDQeo3fTdzODRFK/dsIrRn/Mi/hRS9ByzUWUQITk
lca4TaV38g9BSr+OZJdO9EMWknqLGoWmLPPJbjiGgLy1vDT9NtulP/7K7vNEku7n
nFWYbeCLyPCC4lln7eGbgusf8Bg5Dmh6h6+4LwrnUviAKK8rBLgRBM2GS+ZgCikF
Z6mhlcF/2abw1MYPWSy5mXwZnhXVxjFeWhOnwknVf8Mi3hefzUC8JrRGVkDeCxZN
yEGWeis6LWpuAcnNxwEPymSDu7Slm3Q/Fi9AeejJIje2IrLJazb1FvSZSBHuDJUp
CJil0baXTiqDiSKUe9i+V7iTl1jL079n747tJwWG9Oq/g17n0Ih5GXJtL7R+Ik4o
8WcsnTSmLNJJL2h/PS61ULTVWkxtuWgyN5j4cyt8pgXJAX4GWiQQzq0RyaUeP4B9
6LDzGY19xA1ZqfsqF9ackM8HU9FF7aOaaVtopKjDMxtdepmE5dqDLdsWnDgomniB
czsNJ5omVaqWMthIHYF1oq6IgsCQq7MLECmrtMM1zvyMGheFywtfQEvtR7Q1Rxga
LfIkrOpXPvNsXAS1Xkt0p/9PlRVwxRMD7QWbyazhmyiC4jwdli0G4pGDk/OX8oEe
MmY5rq0EVBRW3BpB/T1I5n8cpfg/82QFSUv0Ce01E+QQs/afd2F35Hk7rOItaOER
fEx2v4Hl9RcdwIrgbgIUR7niEcgz7zwclDB7VjfZUfZnWCW0gbNm5aMUzaX1SvKg
Qb66kXDKZuZe/iX27xlrOCfldnjKVa8/QNg9rceznjYgPOp9oWX6G6aEcPDXAZbZ
hc4ojok+Wm8WgLc/DTaz52pnU+8v1+sQefSVRAcxRcEUnK+lRVAM65NyBPE/pLLF
DkzL0CKbUnyi0hHp0N1pO9UtteSgu6QtY8SJvhhHls/b78C8+FjPO9T7hJZ3bzEk
G5MNv7Vb57g2Xw4G2j7nY2X9qPZXMQe0RrrCV+R6BE0POtTVlg4dekpy3puiKAMY
PnD68f4N7wXS/VBh+ncCXvj+OCVgVpcIjyasDa4bWLvgiQzh33kUPtmFG+TrI9oJ
J6FZxBBaK+Dse6AUYKsGPyFWC7Gks4/uFhEvpUdIISwBYkY8RShFDpJR9ImTZ58j
moqgE+cs4eoZ3jWAs/5iyf4B4A9iOStsBHdxQvEQOwoYzn/ziuVxlRfQa0kCvcBW
MAAgchT6cCnzP8vGSg0pmstdpBvDpA1oiWY6yVlDSefsS47FTYd6bjbKJ4VKkJtZ
i11hsEBefmZfxMWpYqQL2DSDKTP2dwEBGVkHd25wwtEKI5aj+CveOtcU7Ivg9SXN
/4X0sU/keIOHX80eCT4EgbNmDY3AQ6jAauFmlodPJ8RFMU+pUDz4p9kIEaTaSKJk
eX+mAPLXeiRWon1w316oO8IGpzEqLwVMJIum3ZSqyFzIlYOrunHhu4Iv6MXqMYWB
4M/APXSl9TCAzoHSip5/jeNKQzc+Vw2O7L1SLTSnRX0ZxXzCLQAetSnsG3EYfk+k
Zg0SCIusoDmTTSaB4BfvzaF6rKUTLI6MMUg5B5h4lyR/atGU0C2Gao3d+9sBKJOM
K2yJQ89EKxJuZInEsKWF6/1GAmWgCNYgpG0tUpaRnMsUMuhqguhGlhYUuU8yjNf2
Xke23i9myTyznTpu9Si/wARwh7fPY334BjceCG4ZU1mtC45A0cyBm4cOXfqiSGIm
IO9k44MWwjE+tT99eGw5xhR2VFnuU5ki1ORG9qAtMM+iPQINksH/nDSsHD8hCPp6
GkSsqwZJG+nnh3m18ayKCta3tpN7PtDTAFChQQy6qzFdpbmJSgHEGNkdzu4Nby2S
5DuApYzt4xWI5BkJ51sHg+cAivwvNbFBdjxUvx20EJQcFTGhhLBmhaxRRKcpvPNh
YvqCVIadtYRYqEYzsy6j5w1hJWBaeVDfBG6ninWG3xuR4GmPan9GrvBV9Bb4Xh8M
VSU4FJw3xBNQZ6780fsI00qY+6/+CwNAyuElJ3bE/NeFJ2fKJXtcMjlQ2eL3u9xU
u0br8lgX+eN3C/ROFztWRgaoPSzpoFkR8T/9VY0Ajy9v2mqV5F7K7Nmk/kcNdqwm
uRWo777uZ1TlSQiEhWk9JnzgVlfD5eY9YpZXofJagToOYALFVhZNglM/ONdTZK/q
c53kK1+tABINKB/oChK52X8+4CfWvRxjpjLRO0z7AY/CjEhZUJNeMFq9v1C5ClDy
2XyzOu893Cc+xdSisjlZ0RzNsBchtzyI1gIF0uWiwh0i+5wic966clGrwbXh43nW
N6tKzBrsWNoOKCNpcdxfWhByPS4K01yocoIdMONxr0yzd1IZ49kl0lZLNHBguZp6
PFEMKvkQMvWzpuocJTPnci9iZGe2kY/8dWBb5B70TQsxn4Z/aLgPGSMSx1nr6rRo
GKDtRw7fBgArCWvywq7gF3L6OdutesTHp/SaHDnlpE+jRGqSRftuqjaLDVc7bi2L
Ty85npbnR4FH0gH4EOJXsIcH1+XZehw3I1SXzq1oqVzgp/+SVub3aVkzkiYR/V0E
cB20DS87JUrlA6Mna0fTvvboS4NyknYJrHC8qmx7QBU8+UDFD8qXXWyqYG/0DDPy
33rwtZxLAOMqqEiHvyhAnfMBUp8nhI/Vm4GlEgspMhGHpqc6WeybHS1VZblD+OhA
hzETkn27qjC+D+UYNYkzgcfAL06S3cHFB/D9W5yqTu3C3aLxdhq2WHxI7hsckBnt
8PZrUdDBQyt7/o3/2cxjjQ4NthtctwGvMvJqMjiGNVuG7NAN1RBMH5x1otfkju3Q
zm6QIhfjS0q8JuZlljrwPw70ZdjECqccybalkF9/gSYzsycEnNZ+LDolnNWfT/oU
E49WeodsCV+aYdaJs6iJX1kTCfjl5HaNQK+t/WvX1rtsvPPlH+kby4J2F4hd4QwK
ZQv2Y8MmJ9EiaaygAs0S64yDcmiXAF8uKd/VfDYcmfvYwCeRCc1Zb/tZs5q3k1r9
UcKdVz6f8R2jRKnCa3b3ZM6Hfit97xQlRfi+rKaB/gygrJqb/jyrnYPALsgEuJCQ
Ab47SCXJgwCChLvygb1V1Z64AM5xeBpIz0/eUABf3RGs9jnxb5yNCSTgbJYX0GJ2
BngNsXHXoWOlB+oQRlFiHDd6ddobFfxQdyrKwzxwKu4nMaVk+hR489yZ4ATe5Sjy
zTh6l60u8fEzAqOVAeTXEW2NajpiCtlEgp9tJTqYzhV+IAu36y6djKE/VVStUZJQ
MykiyKJh5JOfAfHh7b16fWNjhHHsKnPOglfMZBLcrbntBVAWPXsy5nJQ82bDiEsq
X1u4OidYprVPNE/eTx2k8lb3mvnknuFar45mOTYarkYXbWNQQwtBSyVFucn1Rddp
q6YWCKr8wwWBjxqKh1IM1Bu+roO0Gli6UYrU+sJyS7SC3ZmnyBQ5dj6la8vF55oe
dF4Glg0L8qplWYEhdbSvp/Xi+86ZAKqw4jPW3L+v1LV1UqRLVUpdtoUYXoRkFrbn
Nz11F3W80uvdydBVZmtEVvjsI/on3g3r6LjCqT+9MX3B23f/3hAPkqeeD6WMi1JB
6yQfldfRFJhSLB/eNr/NH+03yawa+5R5ezFlGBUJQRUOM/FSkZh0Xa3OWITLhZtx
YUTfQ34YhXuwVAggliVGVd/ViXbPvgxGBKNHxRNNVIKYwD6NDf/iq9h31pP9TFJV
x28j/gLqjt4WWDcCNhbuZPSZbDfzzCEtidED78EJTsfbqlPEv6bnR2YyoGSet3kd
KFiz0vIwSzpOWvH4nifeWGh+/3tuX5ek7LqgbBFIxmhohDNL/bjBJRTTgFiBijKm
G85d08p/Jtah8XNDPIS13GfY8Qk+iCJNCQ2+KqNcCQDLCiks7E97T+YkjmVZcpXx
80HSqGwGuigWdlIn9CvgyX+3PPqGw0V+UTuSRAURn5KEOckUkWF0vjRby7tktqy/
LcnU/qbv2lgMQsIbi4RkNVF+0oGMdmbwrGCIefzCwk99ej+U7fNrNiK3cga+eJpA
+iEDCCnXtc1SNj4DHiAmbpoAzGA2hi8E5+jqP3lU5A0FXsZvbgSFKUNenL5sN18Q
RudUu9ymjXqgvfQjdMD+fyVZ84JyTtS85rpQ4Qs4J7Qon00OrNkxH4FyAfcJ/eGN
cP6qPYm0I2cmywrtSIxvam2uRtzB7DkZ7IWbzPbQZ+NIMkdwaAtnVXEsUcD/qqbS
rutlTuEXTxf+AB3f47dcCH2JOXnsIDJj29mTBTDt5uVPJU9SEQTxAw+EFwrw85Q9
TK5S1E0nai1BsXvpF40qSC4251XSj9lYXBDNS7ar6xNdrGg+JbnyM2rtR7oZ2h/k
uKWtxOsPcQC9OdGHSJwMdtAwGmZPKfKPyDZrpf8NecC5L/ugiYx+esMVt4zZwSvH
i86v/pdcSBfjyqJN8lAdlW0k90iiEghzPc9Pgs0gUIW2Cjgq9QSxtz4sQXVwrQhr
5fxUHKC7/m7LJ2PhIIBq7g1YzJT651SfF0qTsoNWegEK19c2oqaEQsoySllY0H2s
whzfWcd+68z3j6KplFTR8b4oxQf3v7k+XgyID+2vl/9SrHZukJ/go1RwSpFiRmtM
LuTi+5DXuLcBZlrjPj5ZKZFBVTH5WnkzFt0aAyirN5PXOKsRIkrkF893WHnlp4DR
wbxUUIe4DrWvBdmuloeGstZr5DhqGX6oYkGMpuNMONi2Sk/kK4kLFe5MFh3OAXw7
U7G2Mq1T1tlRrAixgRAZdg9Wn2/EbYOc6uSPG/5ISl5n25X2R+GImqOddaiESuzR
Q99Jrv8vJMendENQVbdbpRZ760ZCgvYw9tBVeoPTLmvPzKSbHNKTheBDyIKeY8/u
CDC94z2cypOcBnmVYMWosFhiR0FP3qDg9dGPbxZBgsZwa9h1nYvgIFzr5btFiZRB
ONwhkM/5TE7mUsqTA7HIcr/ZPQArabpTjVxaZDuS89Fo++971cLuIMdKkZcdJpjD
6q9Iqf7AWJKj/vOk/7eEXGZV9wx/BNUaTxmG8udoku0mAlGwEzrLskam8W1OwlBs
ZY7U7s/PS+I6K+J72kPrZGa5aLVTb5fQ2v9qpaki6LzER/861HI9i1dXbqQd+tpp
HA1LC0XDTFE1qSKBqvWWIKei5xcaAqnSfkCUCEpZbjOjZNiLdY5M56ZABX/R+EB8
tmHO3RtbzhcqwzsyM+61gNRblXiexWQyW2165D+ikWg4YAoTYkJN6KV4EkX/PTKj
vV44TI+lmW9gCqeZQTFBqPYxEOAphsC4zvZ3R6clY62bFUMwy6QXg/sGXoSJVWfL
vJpsT1zjCuSHsJn9YPR+E8Vs2Ea7JgnmyK2aewoB3oy/xWxLXeH+ggSfiH//XLY7
vNLTfpaEj3WpNJGchiGHgNxRNL38Xpp8//k3R5PQs8kO2yzrh7bbU+OjU3IRyGIQ
Yt0OfNE7x2o4VM64mZuHkbfkbBm42vXEfGwZ7fgYu6luX49d0plfg26KcEVkiE8o
K3sO5kBORWF4Ag1LPNZ0gsk9naTs+5uK/UQIPipleUmNOBdhM262vAgtCUDbtvLG
xKRloqrzc2o/NonLLZwzGRbshGpAPcdw3YHky6x10+w+MD1r9v7CTLj4Cp7EjO9c
ab/MppAWuo4lj4/hsxgyVT1dBgEB7NLgybRGiqeeN9zG0TLZoEP/NdYWaNzAaTc7
WEqiSYI2ImAtFYbh5Hv2OtiUXJyyAgflGF+fOF58Fu4XEzN0QffPAXJJtLJpPNu2
Myx2ASwcxmePQ9XIO0ZMQt9FrDyrRvNgEWptOG478nThuwbNRjhKWiT2jInriUbn
vWUUCG8U8ufZ1H13CtWP1zQUUYCDaB7KHidPGznxfM6UiR32127PhglW4NnG5lRa
qzWj+2TzZ19SgOeZR+DEg0pGnbOKPs9e0oFmbTLbsjdu+ozpBHHA4Asa+y56OYfh
vFkvOLAsSkIIJzs+8VuVZCa5/4Ne4zYrPy7xDheVGrwgLG4O0YrWqdmQ1yKX007Q
jO5Cy+mqKpAB+UFEI7NIODqUtxO/K1zLGttcwShAAFD+Py18VYNvEfHegPAzh49j
tzGcs+C/MqJb5ZcLiE/Vqho1fxMmPwVHKFfMm+dXpGkGHdA7pVCSK5GISqnqXPKz
2ZAmQ2gxnokvGi4BLa/qugCHJmCrPmmL13NUohgp0i135d5vPzQ1ZNFm00GIp6uI
AT/EcB4DBB3vcnvKqecl2KtozvgT7mIL69kfa7XX07UtzKxFmVF5M9avAdbbrMja
rihJjac/XUSZR2dXwglhkuPW7WBSEzYFCNMtSec98zbHkHnvHpfVqTMLRpQVtoCJ
BaVYItrDh0Ho2cw+BUVTUXaPiFzmJ5pFZDXyYTtphFsRSKYd2c1EiZDt3IWXSWSd
CWiAhkMF6RtOHgTGsa+531ZF4ywUvk147VArEhGf5aZHIajc/suE4yMv+9ZIZ2oI
Sxpk4O5ZRcE1VWFN0dAN5350zLUwoK+fM+GarXJhfT39zKRGilf14URL4kBMWonT
seBXbWftMlPoBlAVlJsJw5JItPd6FWnq/9U6isIs3/2kOL92JEYe0/3f/uAyVuqR
iaqqkTH/wcAJmndixX22puquGx72N9bfCOzi3y4llDfgWGBSjID87bXVPbxGw5wK
lRFlh2lI/pJ/0u7hdhXas/vzyhWDrWMSlYWzNUb8fSD0PsJAVxl0aIjG2m5ysvLD
xYjdud7xRFYiJxl2LQpuoj65fgYoH0qzd6xU5s7zeYHKjpyhAhC+w3XAVU8Z7QK0
lJTDcPi+8Mgic0k6Wiex9ONBodsYjaCbtB+RiKLmGnVT62hiOMBibt4aHpfZiuS5
Wb1EI+yNrk2f/gqmR1A2+S9RWWj1Xb2bi9gOw6f/zcJukGue7KSoIo3NTmc96meh
aCQPqvQXKhUY+cxydKYU8sjzd1bgmkzIdtcKbpHsw2BNPf9SzTPkcnUFGJzMgoFE
7HP1B7AiqjFEU6KP2lq0nGsYgrGKsGMT1BCJ/Igzanrg8aeJqN9NmlcVxX3UPkv+
d0yq03x/r2Os9gM4bQIHlMHRKOMx5luIOzCXsZNzm2jp5SUvZv5pHByL/TK5BzqP
nsT3Ml2K6Q+TZT+1L2fCbBNOJzn7cp91WBB6luz3hvyOBVEskSpM3M6dJZi8McGp
eryUrQAWOV8m7kKXsrD7F9bpMEdv4M9ClIDijYkBBvjk95yJse5rH4GhoIKi3GmK
WocTFMaGTzr2MgFRxEZH97GAY6C3zZ4RbWapA8qSaQzvhTXQXpHd+RJVp4nuaFpB
GeQ6h2T8bfF9iMyg4FLm672UZwyHUV0UstdEc4lB11I8BIY8sKPEL6V+wpBFLpKQ
xGdQuqZaQO0dwxJQItBgMX8k4dm+a2lQnHitlB++n9fbodR58SaSq1yOBdy/tM5v
KsYiUhV1f41zoIqT3wcDVJFF9+qmNvXWT13hqHyA2s44KL00et0TmJWpddoPuOdr
58Xgf74Mms345EKN2ayPpy+Cj8WMEPXyaknJFHQug1DQQjMPdaN6AH0oSmXKy26/
WgU/of7COqLs2RW8mt34F3JQq3YDynFMfQYWz/6mvymgAcQKHb2BPXB/A27xLhRi
g9eEnO9n9BjyZhfg4mpLHqBjx2MPY1z+mPf5hc2xlFUz4El6y+x2lJVGm80vHTYl
khozt+1G55lufkzEf0rvTIdNBa1VuXBCSyZOJx9AT/173/cDYECgu6DPnddJEzYA
3DBtn6TU27LF+05/nbU1vpdFmqv7dd8gdFKjIVpo1iiNZ7hnK2ZIuea4+K1KLOTO
LkCsoy5KzOLQz+OAdaS0bVXZHpOfHUtTltCCLoHYx0gl7KKKfNd4A2QFYQDOEmgq
DMt8mj0id5MO3uWIw1KhQk6RupV8bMYCBz7XfVMJ6HguTmskf8ZW3awogSmb11sO
oEc6JMezVkgIBhiE3DnxzpjyEnuQAIO7xRXo/h4BNNCJlwcgsBzg6p6QXPXfjVry
cYRwX8eDOO3EVJDv1OwgkXxJw0G+aCujwG3ZENBJoxRvWqac4Xgwc1ETc+SxFNYP
ERJt+Z2MSCDnulW4iIsidIhet4oIJXJB6PlATmvu9DK44nA5fL5Z3OrIvksoWJKf
v4F1qguUR0Ce4psi7MFleEJwMHevTRabw07sPlMGWO7vcfCigtGBihqjBC54/4iR
+uN3SvTxa43clze8A5BvxnLdRS19VK/PQnWOp2sMEFSFJmMKJvmRMn4WMUN/kuW9
VyOo0qMjwlEktH5Mii3tNv0+z3bcEYG2bdbkuqOPnGv4PZCCxzkVBMJL0kBVDuf/
AZlrB75JTa3fXHAqPOcBdVkN7DpndO9o9yf7fxoe8mIOvVyE4M0ZfA7fsXon9hnt
R2Dt/94y7Dcnp0VNjpU1iHPPPYfnzIctIpEb2GlOBwJmjMby8t4xbQKBrbJ+kMwL
fdQvtrpodAkve++c9wDgvQbqnUa1LCUURnBwYx3nuWCgzJPNcfHx79u6nFEFms0e
/qwVLqp6mrMaOCcz+61E6wU3XOGVEDuc5sX3FqthnuvoyMNB26WNNJCsE+xsydgH
FHk9kv5nlLAPMaSMvdqBRW7n3wI3KBsvysnbpkLfsaM1Gq0TRBflVIqp9nTDlb5J
QuKgOWMYN+tmDCUzVwrZcpQN9PWPgXlKT4dUVYWng4BfmU/WXCdixv1GRROcu2CF
TTDkctRtNFLGLCs+meBUHticdHRURISDTLAgM0/sULWJhVxXqpZTmi79zL+m1nl3
SiUOKZS9k3TFB/40vIECusMSfUvjpnAmc3lzVm6nUA2S6OSGvxmfoxHfloLg+2l9
NS5IyDwLg1G/+SwH8wnHexhqS/KkfEkiwopBDULlhYQsIAi0Ki6MfWG5/KNeyTUf
o8J7g0xA7svKoPPXHCvd+NcAO1vdBxm2YC8dmtq4J7vzmvtOiAodERlRBOF69JaL
Yin48tCjh79Iat/TYkKluCGLQPNFqA1ZVijUhsJ5+lZkt7zFV9nIKpSOgvKlaPBx
pWHQuhY5/9/KYY7QOUrIsZth0wqfYY0KC2W24rp8h/JmkWdoXzRpRG/DXG07bEIU
HFNIkAHnbeTjfeQiDMqEZOAXfo+FuUZo5exjGeCBe39Lim3LfO9pKzffwYoUlZqI
SPb72KftdSQlICVHz74oGYUeBbG8ecfbaD4B6WiHOzOZO42tlZ4v6PFHbZPs26Uz
nfa4/NPumxvU0bjycco2Q3vGsXJriFXMYCXYv/+U/RJwB9R83LktmWiGV8HzvZiY
U03OByQsslSR12o2btxl27hLd6SNr+OvZSYNmPc+7JICN48RF6pGlZSrFmTEnDzo
UVpv9hgJjYv1GNQwuIhD9fdYY5fm47dQDJ5IpjSNOfwizMXsf5glcFNyKoFv1iAP
2pdGEKAyjQ+q2rOuDfOhN33tIyAYHvsi0r7W31KP/UbJ5CDY44DnXavSdT/Pr2Cz
GFJ2T2XHj+7Ed8ABGTf1E03jsUC2EeZgqKyw0L6ik6gQ3gCKxRyjwtaMyBonyxKH
OXXpLBBopTNJwt7RLSfbaSZkCB+1Lidn/eAoU+xhXJoLlPGjCitaqYZHd1Lg2N5l
bM3TRmFnsfc3EJjbcjiy14Pqw1bh7jZrsIR6EU08Ljl75eFq2ns4bWo6/OW03YqE
i3l+KWwCarYfEg7skfbq5JwgDZztaFxRxqWMA2pG9TxxHynbdI6e5JjTM7HABSmv
lQTmpTNQstpU5VHojEQCl72olBrwaTPatLlzsP2egpZ+Or2SVIqRFxfUzOZxFCxJ
Aihu9fs6twTDYOVvCGUYQm0bJ3xOcbRiPx7dDLL8V9jvzNj3rWXzen+OYdpy1dNV
fK9Z/7bwP6hA/w0zZ5oyySduvfReq393c4pj1LSuiQzEk6lTBmOsOi6aWHMF4pW8
+0WfemOD/sY95dz1/V/gYkHE731wbJYGsWSjjfwyukM1hY3GFbYz5T1tIQe/QD49
ZCvuRRTd1Jf7ZIYZhAnUXCTqgpvZ5nPj7oXsFWGqEsNlZ+NFqTx6e2PKJbpDh8h1
aQSXvZeDTcJj0xyzOi73ZgyLvjg4ShT+EnJOB2sgmxo4At7LWUjUkGrXcQPhsgLG
JA/QZgHLcko3Aw/fDm2G5ViL94eSK2kT5a7Xb9OGdv8pPqEcfkGgogKFlUu+TWS3
5X5u70VHa5O6bU4tLqy/hhJg5hd/McTk21cIOUQlf/PeyjF2a2DuLoYs94ehD1H1
DjbBe92Ek7uhri6q8HCibZWJefunjqhw5jFSjwudZHawRQB0lV72D+Ivf7gRade3
dd+nMfWiYKBt1XsieqbhSkrlXZdtj+NCg7VqZOjCAP+ozDDWptEsN7334BdpYX6B
lYqtvcypZ8I1NfBOPVfbMAyjdRLiGtndf1EndYWLuz/1XWclfRU+VO6nZngNTp/+
0ljHBsKSqnlOuJgy1J8sqnsMErNolaPRBDHfEvODRCKcQYM0Y2Fa5JyTf3gQvMk1
bcJTnNTot2+8g23sEnbJxYSLX5LZOJ2MJP5OynLKRB5w05T0pHd0dusizv+7ZXMG
pNfkV27xUZ24CVj+JXM37H1ZghjOaLuekTsEYwjjv6k9pmGhIOphnMoWgrfWVH+0
OtEOHGOKEuu8DmewzgrecZPG7TKIyc9JIZOSjNiNaY66Sr1vlM0OFzEEk9vkAG9v
RvmbXOQp4erjVia5n9nbqUsyy1YfL27dCbDwTqKanqSOTLamMv0ofel5vbyVRKns
yb1ciVPQT+R+ci133sRzzJF9ASINao39HxuIaQiHzslh5xbGIvbMv8hR1IPr+uwv
CJO+GyR0gy6go+FIFfnPzeOsNfhMohv5HvVQhKifMW32TmjM6XMcGgTZfBr+l8Rh
3IeCFfXlHqdpiNAALeeqorTUsMxghYmnUypzSS9TaN0V7fSBERALBjnwTSD1N3Rr
tC7pIw1pM5faOLjLIPZBCFo5r+2L0saZt0dImuV8pjn+RMTe87rwlD7w133RQrKP
T1ZTnOzaHwYTqiFSlBpHmhPzbMm5+i/apsQhSLn0ty5nK5Mt1+4G8vRfn0GwB44i
0LwUzFuBvsldox8Ie7J7EiQdq+tI5XTQQuBLIJRcRluXoXWj7udu8a+noxLCOot2
t8wrXSUMiNZM8NkHjH1KzqZeY+ek7UJvE+ZCHOFoUXRgbK4Yj2DeL7+ngK9/cxcy
KaViDq7KnAPAPy2kfXYGDUz/2AneOvg/nV/T+hZNKD7BBBu+90PQVc6JM332pO+E
l6WBfwTD3vCLWhPwnRlSOEHMsG5lRF93qhdOituyIfaVyiQeiBXotOLsg/IzHbIc
1L5C4+hbQwtwfwCvor9Px+xqz5l+s8uLStOyEMLOowvq93J/5WWzX41GE/TLGnm8
w9viybCrYqYk56BZYwuYOoGSUZ9x0Oq6u8mrQ1fGYEl37qzC7pc/T4EEYCGB31lh
MgMCRfP1ricuGIojQjQsqJMG2RC0usGLf9RApm3ABMqsWK0bioL1krGxIb/0gKCv
+CdHuXE++eP8EnBa9RU/jDDXQ7bThouRl9OsSlgQUMxljBjInkKRYm4FiKeJJhDD
iGKuyV/JjeXuJzPuM5deuzkBKfxE19wqj3pISmwLR3gSiM3gmLwn6BxgUD7vowri
Mr8Gsk+kHBDurayZJpPCIt3lzF3WVIJY8sAkUftP3FoaDKFjuWQEhglCb3uVA1/v
ibmUhPxdbaHdg2FQbCL6FFmuQQ/PbiP547F9NPM23F4QOohyckIRuxzLCTlz+63t
JJJaWY8NTxSDPB469YAJd7UaMUNsdu2kl+/PGJKMjuRUXubh0xG85Wt8igStUSoa
gkdREUDnkLijpU1MODAIeUjnwJnMHkj2m8AaV64veh/H60EgJkII9d6IRmM6nEMM
KT66b3YvVQiJZWgvPXA3OUt66YH9ncYLyWbv3Cn9IVcmkNxGrCKvi7E6GqEk1f77
RsAWCoYyTwcsNpD2xCrinXfHEwnIm0sNTlVU/Xbjc2PPeVg0bXuleBZVQP5sEDo3
T7wSCKBWfMs5myTm9vEbWm19V183OoW+xyJsHtPqtSpgoSPG/EiobKvkg/qyoFJ1
H4qdJUlpBJHZvc5uxrzH/bh/3edcCI+et1VafQC7BEIZIM/GvCF3lumdIt7EmWfR
MJ82ONohxQWLuF/PiKdY91gFMxaPrxWta+y6tzfLv1mqICb1JAJJIpwdqjVguL3s
U5NSCy4ZRzP3zSmfvXWaXQ8ty3fpLzr94cMVsalUV+1RqGwVxrLPQ4a9lr5gldp4
GkbN0I57VkirwGgCqlQnaMRjpiaec5td6bJj7/c9lHupNIc7iwbs/p/T79EmQRe3
kO+GfDgSghKq4Ah3HOVxEHeiVEcIYabH6wlWBihOlyjclN/VJdErjaSYMJs9hT5k
oj+Nkniu8y1PZJUBOSbkLkNEZnrcs+zwAygiAjlct2XHIIx1DxcNw7pAQ9kICT0e
EviyBqtHpurfpmfO2Gd8XJ0AZwqTMkY+pNNF5TCivTaSHjt5X7jSynEOmvjjTeHf
NxxlJxS9nRpx4s+WKbkNicKc0flmshGeu7Rj1XUCukfZkBKMtEqzSBEI+VsK6ALQ
AfirV5FobFbxrKDdxduRKPQ3CNMG0LPmlKuRKMuZO/0B3Dpy/p+VfudnUlBYzPHn
+YcWL63cRsSZnV1TPxhVmTHpjgntxjeIYGtHVTN/WlHfA36T/nMbrW4ErwW36LKD
qAAzyPD+C8zPEzSmO1NiCBmDeOkGAPcAqGsgKO+Ki2uP22xEYyAUhacUKe/I6iKN
VgMhpDXn1zHr6z/sMNoVovs2PyL6p7M3mA/pStnZx369DBiAWesjFaiGqCM8jfGU
lStAMaAQJnbCwrC/3gNc7mJMMb1sJ0qj8BzZ096IpQv4Jy/1H/4AuOBmgggxc1kk
rCGsePJj5Xrvlvr3Ud74ANZ+s7TbpN4nZyi51rdkzBpIjBGIv2lvufaJSkWTkJoA
KbT2iagCSsvi0aBfOtrEIyZsukYSte3m7AaPEq5tcGadi7NP3PI6T2KhpfgJGiFF
DI6CUCjcTgU4eeT+ysJr9mc/AHR1XFYBH+2ijS7IEVn9i1vD6BX0rMG+OXXMe1Cf
c0Hllq/x+titDWwoz1/JZ34USgGhECjOo3nGf2sbk/PP+Rh4RSR5R3jkaS3OtzYD
1Vqfxk/V/y8Pq/e5KQp8KoA7oUBAlvQRfC6vyYEPhEgeIKRzy4Xv1ZpXb0/LePP8
rySv5jT5imXV92slTe/ssqEaYaygXpPiUkEdOQ9tPNe+j7PnbI6NjBYQaNOov730
zXIGkNhmfJrOSzf/jzTzzQ8k9ykBhpm/p0phHl2bavS81CfiCG5BGxAv+1cT1BKm
G7e8n9jwFC8Di3/7GKqVeei2NjLlBH51xVJ7Dsk/690DgPotc5u1mUnc+GtGesPN
IUURQy5DKXhLD8T8swi2GucODw2JVZU8P5Tjtin0DFXgzavPDRKBEGO9pCpTauFC
CGxBi0ktO9Q/b70KEm5+CmxqsIgQbOQ9n/AqGZ7+Q7steaYGVMMFVyZft/iOGQNY
Yoz+zyfx8ecXkSniBOcjyjlHDnRMyI+y7nPO/43AiCgTegkiO3C42bvVnBMJZurN
Fux2SCEBH2L2bKCcdg69eTc2mz/gIIObxb3ANHuQ0oTNkZshSp0e0nHTVMbglqgO
SU/MPxGmPy9fgccLbkVcJ/terUHgX7Jz9MGqFYvO8eNrInB24hFf59uG/Hl16GVJ
tNDymZ6LMtd7lCbm4wjFPZqFK9qDryep8sFbd9z4yH4bvAeeZSfxfmV+n0nR4YKJ
3wCAFqR9J729iWKj70EU9/kcYqK/rrbyNTZ7GEqJoDQ2b/83uChPh5SsZgVb8lQ5
LgzCQqB+xgMjB6gucLpXLLPa8Z7FImOHlrcpCS1YesNjkl4MWUeal/8jqGSuWbQx
wlcGDxAC4dO/hXneJTwwd1YwuWxb3pnXBr2mJdDKM/JCvQUwOtVis9k1cwrX+1HX
zjSzJtceiVOK23r5hDCXujzfCY5Avs2LVeOVTB1JyfZ+xBMnjS4fBJx0B6TJhSOF
GoCjwoJ8F8F29NO5saz3Z0NaqHHuGg6opp42B/JA7tCAiOZowE5lr94hHEIUHmD4
fSreCU5mqre9XzdT5HXuFyQ0Smt0KA3tYoc/xHTNyd3ODgIoHxf1t+EGYZiV2Ptl
PaJSUkbfiqwV0YMV/RfOXo9/HLG+a3tmj8SUFo+ihJkgC/StuB7OVGQ8/eA2SXzD
ROVICqKaNJ81appsdQ9WQ7ChOg2g4knYTI/f9lAPXqqqDoSS6Xe+XkbJ7PSt3lQX
TfTuIWGKnnnxZ8+U9+7acdgDGweuaio8AhlIgsZocd9UBxPPtNQ//3BQ8LZ20Vdg
t+3dNZ/XGz/nG/dFBWZ88isAfYiQweYbeQPF9t+mg1v+7+vvvggwpmh6EubL7I3R
nYX0YoNjCQGRGGhmWLW1AGh5uDap92Opz4o2tflbjxS1ydgzBF4LCszuWNU4wG2N
sDV6uLs+9VCkAhjTsTBDCwMlafUcAnYEAZrrQMElrB5oyYGDF5aaIMyaodVbnka2
iktHZMbLWUR7WIVtSik0CcfbnL/l10iw2IFM0kcewvpkM/KYZCoG4XK1i8OzXH7X
KSsBtvhzHo1zfW5ri1YsYugyA4x2Jcm/8U9f8V7dyjdf9u/ZE5xLxPVjIcQeL0hO
A9Zer08ereJxaj9MkmI9KQ9HDYvw+SdE7UkMPJMZPcpe0T4/mO/UeD+uJ/nS5eAh
BYrhYeP1P34a0Sc6tik3dM6ub6Vo9gPegjzZtLVRoGJbx9OxUiKaJ/5AiPpJa725
sAmmpn7anq62Or20c0d6C4lOZb/E19VfThFvWsSvjibvjD5oFRvxQWSg34ao+iMr
yZlfPbi7JTTerL3tASt4HR5eMuMMnIsV5KPblwAvXFtCY3I4wPrLUj5IAvu6jXnc
GaAQAv6jQNsfESC4iqPY2k+ygcYWk7WrqfXm6XewEdIgz7FQeIyX5nOF3edyPzn/
g4fsdtmf5W+naMIMlpYCZqflxZpJydcsaL/qUpe5k+ApgdO8/dxO+X/+qb5T77Wo
Kuf4hueH6a9eL/py2TEelEgxlBqW7I58ly6tw65E28+G4belmiqRUWups2nZK852
YryNlNGvpOH0NzR/GcpQjdaVun9gKXdnB7isgTGBtqUroPs/DxcJWxfBZ6Bwhd8H
eA2M8P7H1buWPs5SALAn2pB0UL6/LEYxaDc15P+8Zjq6XhpEjUmGHyyYaqJrm0nE
A58zu5mDm0saGvtyvYlAh7E1KhP/2PFaS5xyg3mvNyxPBDMoZVhDLxAq4nX0q31V
4qMUKFNMATi2bGtFgsQdS4+gMi6BXG0/kP57pA1zfKMKnM6Bt4WalbKMbIW47gi0
qQ51qLlpuYdaicI1a7t89bBX5y5ZqXmMCJRi4dnyaSoNZJ+DCM6t6cJD+gFNjSj2
xhyKW7Vy1dOnbhFxCEEGzu7VTmR7ZIl8Mn8EmSNcgFyKrkf/q8ZStwaaOTua5etX
tgOwqCqy6vtu3teTIGu+1ppGfHMTjOQy6y8cMmtyM1oBY+j3EEgErlJxgKl9b0K+
nMuetEN6FTrrohfwRgLavd29zH4xvOA2vpcZelU5ygEBwzkcOM2Z9U51owY5M8ky
C5p1KoMi/7K7K9fiKo8SSt/cFhgkVIqW4dH8e4E+2AT1E3ZCHwNUhwwrfmygSNv9
tXtRxUB8Owx1q9Flu3MxZQGOfbfz+7SviuMvxEXD/jQ/8shfIbF1+T+z2igliHeY
n1/GDHaWz5mGc+PfRiRcnJHiiFdJIjv2juSsCJQDDVbwWrgc6GmtBsFq1AqyGrHs
Cd+H4kIYLqZFfuBGIKnkS4IQe4vUtLcStDedCzqzbmh5v7aAmm+SP3o3RnbIYjKG
H+/x5ZfQkpU2lsS3KPSej/8fq6KuTXOPxA6BDR3JHP2Zs0MQ9r6bfCap/2T3/+PI
UjqQKiBxhsbF+cvngu1zeUIRIJQocHTqoLiifIRxrOVz8lyWjJQC/4bulC8vg2UE
fwwuNisyzh0lyKAlhrVvt3jOd/dCt52owj9DmbgzLKT+ZcSsa/Tet4gD93OrKF4G
JC4x6BSpLj5UYIQCrqwj2sCaPSvTdJwXzLXgNrJ/mhq9bm2wxChlYp1MWGTpkQkL
B0hxEXOkCVc1v7hGrk8TK9bghyPZaEA6/Yo0uDYOQ4TMpj2t30QEm6oC0qQ1ZnTM
oxuKD5yVZud6SxBMQ2af0vzJKgcajsl4zBukTup9vM6ChkvAcd5w3+orTv1lq7hG
54WpLgcs5MxGbAjTP/aEhl/QQ2xjSX4ghrCEAhJrmVAgS/aBUmB1hD28zdiV4ZbI
zC6bEe4EV5US+ZQfsihk7Xjur+Votnt8F4QHy/l5sW1kRIEcEQYo80G6KCwYnav+
sFs7TbtqyeycTexGlWp+pkVgYPNGMee8OuXBEx160rJySIWIJX0dVNQpie+rywEN
Og5zU4Eh9eRjHgLTGD/pO2OPpX0vRJRahYpDxhV8xTypfcN2tuwjXoqDmZtak/LT
3FPgaLIliqH4W01Sl0Te1/jKgqvAx3LyBdmKe8CtG8E++MgpKFEylCtlwM8DWfMO
g3qT/Lz/J+cr1Nkb9KkRNMKHDLe0MFbWl+CDcMOi+tVG6GujorKeHJCDgQ7jg6nD
C/LESEA5oCql9hnzaZslyNAErnDBroEmYhv/bh4cfe6mAV73EXlByzI1UQWQo/04
imrb1FDD5DpsfqGsMHo4rhJc5DpbsGx2Xv6WiLKdj+p84mID/vNqF3BWza9/ha3k
Ql/AAFNplNleUOjAeYZ01lat0iUJn6586xnvOH22ETqX0tOjpO4jz/lIRxtu3rOB
Svlr6rDWz1fXFYqBsPIqcKRAoN5UAWz0U25NI4KNfLxJBjq+VZxQkphCX2SjUBG1
S3WOVZf5TqUpp/5r3adk84qcXcbOGY7emccIyARclFlHnxltmsMYttU0V0zkBqHY
ZG2c11/9+LVhpWoItwQOGgjC25PFPdlXeE/l1jGQtwFp89SLc5YakLBzU2nF7V7y
B8Dq+H007apXp6b2yCnVBPrYdSKLXu3r5kV2QQxO4f000DR227RaQioS7LE/m47+
pPbhU2hstuii44hAqd5Xo5o2baQeA7gvV981eIqRc5/8vX/X4Y/Xv8P0Alwr/Yfi
Ws+PqPVLKabTGZd/AiFHc+GgfYpqsL10oYVqhBi4AJlfTTm1p5bm+ZjiFnqMqA1h
50GS2Nu6QBR5nyOXujOW1LfBgTskDgObXtN0OQlCy1I1Qp3Jh/3frMopvXrZE3Hl
Q836SEmF9/NSra3sUWxP7RMxnnbg9tovF7ySvjm6Ea3cZJIow2H7Tvuln5CJnX14
4/Htk+bY9Dskyp1ASC5hEJ5xbkdV0DPB++vOqNC0X5w+h13Rzp433I8XtJvEsa0z
xtpxtGd+2yfKwOVAU3pF8SBTapNwdMHmki+kF5EHShuRXQI8YYJUbzdWxosRxe2e
g8VaY5Ucg29/k3WklLa+VPq+S1xYY0KZ2cDti8w3U9RWvlhHGIkZMPk9sVwsPS2M
fLEc//Ai+snbObvEQAmKmp1vwezJnTf8+ZMW6SIoQq3/7ppjoPiQtLxL1VygpVGf
7ULsOxMSUCpd6NwvaM+CQxP8gLWi88pIAPjcKqC/I2YssOzeryyC9y+LgRALkr3B
TByj/b0zP+iypinU42u28v+zfKTIYsTz7NWk27Uk11oXYQQ8XjqOJ2uXvDqeUyAR
W8KKWQuHqqu4hIJngacer+uxa0BSiJzjdfzZMCWnOesDQHK0/X/ppdkabf/m+tCl
obZnfAt5kYjsVlDUKW2/NiLnl/+SAYI8pX2qNaXrISR9dSxqX5HiT1ay+fDRbhpz
7e9UMrF4OmCVu5BkMD6zsglUBrZL3PU5HbfYOa2mVSNMF3C0Ni7k0nvgnxrtR2rq
GgzwlJYrPHrlrID6FmdnP2iepw48vPHVkNoTnzX8K5BAZXn15r3UhKgTMMK1kOAs
RMro7qdNWhvjA7c3DW1fnL8x1vCSwJFG7023PfdOmdQTuWQ83Yz3E3JVsUeOGy/R
sTEI//E9+P8KS8nJmBxFmq9JrqV9hnLLtKNWgQGRvSqMm1ke17+lXtCVPzX9pZKD
PXYTzkkF83TyuuvSTz3u260jeeESUBXGURaMMvDhcKwuoibm/6yHwYytKYcFoKv+
lJp2IO90N50YAUv7JxpTNV2pSvdHPnHqaHfWL1mrciAIwtR+NEKbgBDDgbFOMTzB
CGa+jJcNjJXCs207ufuWjPxW84W5Q1QGxxcb0TCb1anq9shzG/HR9ZMohzxeAQzT
ZViolGWH9JGWzOhkYzkdUim9RxUZnG4L969FJMGNcMVTxe6X8/9i5IiouDlbKTfo
IbOL0hghkFJaslDSFcPKt58x2RBdDYjzeSVWD87H1gnVs2R0iPp923iGBmLgL+7S
qhJjprbA5I6Q0HOghkoFyXJiZvs09cZvqT6c4mQvHKhsNbrATWJNxuf1lMjkzMQt
6Ij+eW82YjoD4O0ADlYVyl63EfjYDIZ80lYb4JDn3fJAZ8Tl9Wp2Q3kd+/ac+p9p
ddgCCfy+TX/bR5JL34Nktk7kJ4vNxcTjtFdmEtX7mhDXQKy3opKidUnS4M+aQVtU
3+Lt0Bq3/qG2vOf2dQ0Ogq5M9vEQIRsPOHPwIPFAlmIucho0pw6ajLko9hrMFGh4
YJIc8P2I/+xNauoAM1XUas/VbYFb+r7J1TvbyzaExm/4kxtbwV5IMrZTUyui52lS
rSBEHC/rvHDDWtsP3S4WVes+vu+q6yJPINXN34xRGTalLSIqIjiqAOtRW4zgeoTY
RWT0D2QuqM8rId52hFk6Ck+HYrTzi8o7HWpLJ8B12jmCwj7qVHCAEjni79gPAO3L
frYzVUBOAXLBJS6Hi/lfwT8BHE8QhsgvZTyqRJKUSRHPxNu5AcIkd+No/oVxljky
vSr9hUHfeKg+9czwnYZXvwvNLu+OJ8xldlAhpsu6STLGTVgD7cdZLMNrvXNVy8r3
CQ0gDadDLX4u84EKJU59LQE1lLpwD25i7SfDyWSiPGzRwUMXjMj8OIzQcR1gANWh
lsTgGhSFoDNc7DDbKmHEsMMlLe35piJI/PiagjooZG7ogtJQVG3DFURobxDi1tLJ
r7phaHG7BZsMJ/T4e+hu64uYc4cF+6a5UZR3e63Gx94GBYEK2vXCgCcqY5d+bOgL
lh8sHGH8xrWUz5gBBtoFJpxsd63Px1wMPyqNVHD/PSCBswTlYpZGwEbz6wiZ55B9
WX9+YxPQ8Uc3v7WN5gWTy9A/LQ5n/m20dv5jN8wXRQpsywgV7909y2qPHaAERU48
0zr6WILKnobcF9OpzQQ5EiOtNml9rqZbKj1z9iW9aI4KC/LfY5tqzqjll3eKqs1H
7r4FlWCkMjaU2HVDroSb3MOnMaRz9jodvPza+NthOL6DOAddocp59T1xm3XyY982
i89ouNPRhNhO4wujZDOQLcY49sKOMTKJtjYNn1g4W3Gw6lblD4jJ9sFoAdKK8q0M
9tTuCa1JWaCQUHTR+jAM6C0+w/LeSw+XMxb0ZCTI6UObFO7ytleaSZ9wQmuYRdoA
ow5XAhybYnis9zG0t9vLAvYs8mMng/cqnFdert6xV7xLNYo8Jus0ajl8/b+4VU6y
g75qGp+p+QEH7oNfxKVzbFTCCDJ5pnpT4c1zD8JqWJf+l5Tsjusk3VBGcSNJOF1y
kBQDtQIl28Cj19XfmvaJp7AQxD1QGP09ETeKhqD/eCCjWyKuHFwfLTPjuBblpAbh
C8VS/8kKX7BGOGSNqWjQjwqkNj8WcL0cCPLJMvGNyED4ru2zRqmVvqO6OBG2bxX5
7oR0zoYnBD/1NMHqlWfFoTfyUGrZcK5bIcpqYSrFfHNckOq7P8peZZALt/cZ0nhk
UdlIdi1wL2UVxQrerHTn7Ug1jdPwvFVtrcO/gaxuJ/wbmBIEZV1VMXvgYOnL/gzi
k5XeILUTyCMe9B+xpsj+5m/yFR4PmVmBRUYiS36MYoXc54/enpGHORmF7+MuD1lb
leloZWKlqssw87Bibid730qA4t4xSmRmk8YrOivSk7DApUpVGDU8xZouSyb40i8i
lMnrrJnG2vs2qUkTBag5PH56+xw+wAcBXXZcp4bv74Cj3qNKsKaF/NNy1qlZ7mX8
iV2FVYMYIF53NUvTbHbhBR8YxnIj+J0lvYFpJeY8Iqp+CYBv1VK0rYMHk5EwboW2
9OLU9BroWYHu1I72wT8T+x1O2TtOVBtRncHb+hLJNyyZil+1PBQH5Rz8D7N+nfIM
1K+1X+HTsxlWX96xPvde3QAjNuKU44zxBxu1J2vhZY6p4hCVaRO3XbVa+6U6UdI6
3g0sUN4R9L1Eq7ce6BgSzicD0HhyGY6IZkp6MCK6qj+lMO/H6YtOfu7bTt3m31pa
zxIjlqKhOJPnyVnHs1ik+r4uqndx4QOhEWhg9DedkFcnLQTHqtKhjcdZ5lk0wWHW
M4FTP172Zrd2OwlFcq/YtC3rexEA+R2BYa0pvIZcjFDP65lCg5298mIGsJ85CtpV
jlPCu88RVc6kug34Awlh4OoVMw7dGCraRiGUleglY439uC749KvyPH7sCvet6aFD
8tVqnVhMyjuxcN+DpDbuGMQ0tYPSX3jbc0PdTBdzBWfXRcZZhPxANPnfIzIb5psF
ZxEl3X92r1Op5dyO+Wcte1Y4xT/dftLzhCARCT54tmc+f0/if8O7PlTejh/0ci0y
Ih6IYI/6gNFVW23i7NabMrqUi10Q6vbhPiSA8tz/E67gKM642UsvjtMhZgX5ZESS
ODiy00QR2LxWBVZxxdLwjYE55QNLKvGxzCr98snrCNQfZSL0u0Lfi1izdvtdCQZx
wbVIlBXKfNenaaq0G1GzF15VAB78m3wR1v5TPEhqBU0gqmdE9ffce8fKY5f1qjB4
jfhOG7EHENRgYnScpm7ZVDPXB4WALEddJFB19BZ9990BD/PPWZs2xKqTBrRBlC7A
eanJfR8+mxZElLzQcRVPWYGta3NKY42naPRxPUBXHHFzPbqn3YFohGqnKfVmVxj8
bs5XAG1lKhuG1SbA7xLMsNxjShL4peVzQOiGiQAxU0mqpFQxwheeM8oILjYDbhQJ
5mS6V9X7Ezh8hjD1hmZGAa9gVLqHoe7kUp18jhi0SmhzIa0C+jHG/WldGksh7fzS
f8STio/x1RStazIJ2DnZG14Jka4s8aNfSgN6g8zAC+PteOp6tOraMtXUkbWAG0By
OzyyRy5qGs9kUGix55pLPlK2asEcHVVjWdVLFHGUYYR232X0JsgTTI0OVzpPUuE5
mQEspvoYUuWytkkucBWSAjSlVnOuA/8XXHca5zec75XXc3ReJFXmc2MNhYMeq1wy
yx0QCMNzOjRlfFRXAT4m8qc4UQ9Gw0DCYwlv3N6qZA+c/vLhyBbbKEmGZJZKwg4m
Jbr6eYXGQujJ3Gnp0wvK4Vf8SDiPHxWqZe4jBw94p6VEiLTDhCkPu/B7S+d3+RuR
yFHBHb8OG8u0lF5LFDz4nTeCgOg9br3XcXjaQaf/3qrCWKYhpj6whWDw0TOIYIhE
ezO91YE37yyczqQ2Nn+UbLxyVVChcavPXIe6RRtHoiTSr3z/IXxN4Xg6/Dt6y4Fu
T/QSAmBJl1MAC7USJSOTUHIC0Kvypc13ke2tZnVhBQQopHvcdXgoWAd3Lnt7BJmx
fPD1FDXxoF5JfUFOltH1QMDalWy1czfsRye8f5Sc/vX9zU4Qy1G4obOWnKzcfxIg
jobtUh8xnVlJAPtkEYKuPGpvA5go7ZXD14vq3juy9S8gdAKCT1a4VyWCqTAmKHc2
VUmjb4qk7SraYCDFuLusCgWbthLp1auewIM6Tm73k4WiZe4ltxL2bEi1JnAoVngD
f12zkBd3nUEliSqpqa4RRenivccQ2aD0YfMEBEc9icAZnjBK5NeKVsohJ/ms1TXb
uHoPlIdUJb8YMrhzIMytksAHjGVKJWf2yVKr9yMb4OXu4ALGg0kYMhxRgrMA0Suf
J/oWs5nZvjRPaN5OODc1LNa8zkAy54FMlw+rQ4hX1C/yFptMl9/VDlJhDwReySym
UGtLJ/gRkHFvSDkL66vMp+we6s10xos3NrCZplB3fdEwdTfgiAkO0cvGSagQISJs
pGVzuMQuS+bX+wYpHoeFZlp7XTvZVdixW13CwGieUmWxpmOvSSn14xfsDUCNeLeo
jJPWx0lnvBvCyLZ+dkp/uYBg/SS7iE4RRw5gIbm+4H6SXmLEBS0lXM2cmeFq+jpZ
uaDOvK51WRRn3VwDFZagKhPdza8WmTPzg9C5JSmGuHM1eWyXAViXJM9nVCHwTqAw
GoYEiOMX/2BN3oIRS5IFQT1NGXV0XZgpFi7m/3R4p13VED36/qk+Kk00qofjMqBf
TY7Sn9Coe8sCRJkqcK/jJxjZW6ZOCPjCT450LwsVwXMo/mbenO7cF+6yEvtaQ+7x
atOnhwr0sNteunjOtPt+MbwmmMat14u1gqzliFv9sH6MZYp2n5cFd/lpW1aVdToa
x9/L3pTxKphaPh0shNshEOsLO9Ud0wSKFSiDA5RNax0eJd+swy7hWQSAi/6qKYAn
ZAmKJ1pljtnqLu/ZgIMNaR2Cpii7cdqmfqJDuAWU1BIDmNrab9+pB9DCHuaCIBCB
4kGOQGrjIYhN8PDZ2q244wJL1iwKwxExjd3BuT8Pw3mF4qEtD/Q8/QV4IEsJtL46
SUA2CRneLUgPJy8ip16vuuJvxmZEae5wzynBmyjhFZliCN9EQYGSIl7u96qrMXmo
6XRAiBs4xPsnIe7ndD7S5VtLjNrCMICpIh7a6BlMZ3Enw/dVCgnBR9NWppMNbJth
6AFRFMXGDqHpJj+MEHc4WtFIfoMM2V/f3mdxp+oeCCojbzkYOuvSKTjP6Em9SCPY
ItMHDp8jlPso817RKUTz4Hz+3IWOO1iV2G+yKIhh2BzBGdHS/4dQ/t5h8GczFdbM
TdAWrPOFWm8DKxmPAvuqdQpGZjtOwZizUnwGosR34fDfZc4iTaBJyZEiYR78kPTm
4G9+HkhB5Xqm/fyXMaGZVxxmXPIfeZ3OxMT3GGThSK78VJhdVIhvXYsZr8jBpPbU
iQ0L7EcMkBAelZGfrM2KdyB9xDMz7cmJ2QoxO43y+EOC9B30FdngdyVaemym5Sw9
YVOZJqWeEbINUcgMWJ+ccAezbYUDMxTLO9fivEdl4FTp1dtYlHVUPTW9ItQROFUQ
sPgPjmMK0NvoQPRRMOYJqma/fpEbeVxdYhlZwBfq2rVq4C4b+R2PEY/FHrpKlwGx
uI+zMHuxDv7Wh2yextd8ZjYgu5Rx11LxPtFCb2Ww9t9mQR2RZGbKk6b0CEWMlhrk
DOIyHnha31vITnKxL4QXz8HvdjODfl4BDLWZljz3NxEwzsGBd9kdmbKRGz+TVizj
OnIf5W/GbODg+vNH0C8K9bSyIwlUMaMv79d0ol0agl8hAbp/j977zOZdDxodsvZV
rdibj5PC7BSpqA7PCWSvB8q/otQ4sPNx/ae9dzZNBLKc7SRkLvj3zC7yHvu3hDHV
M0okpOdezj7BaDOPDm8Ig9d4wWO+BdA/ybcI+y4GUTDJ4CUmMHiDjNqphNuV5MIQ
LyRmu5jZwcdAxGNq4eEMgGy30uANqosbTT/TMJdPt9/I6VoD6pDuuhdQEiE09QeW
dagmzoYSlLIoOZI9v/0gpih/VjlGP415/CafNFLw6sPj4bS7idubVLXsAOxY9J3j
N6rY6ntwL5wENervfSznfr29EmiMw19Tc6laJVNv0RfQqFtfkjAIkhJEaVZOXcE0
yoyRnYKm6aY2qxtshY7AEko2WlBlICr4y0Erwcszh1QPxhE+F8F9YS6bCu5Q7ZDC
LjCTup2wLnwdvmrOQfOKIoxwWpkDUx7ZnnZyecqQdiF2yTQEYcSthxdQvYt0qh0L
uiKzOWWf4mMRDj2Zpty1ZHqAbHYC4YbqNYZqgOiigvnA2seumDQAdaEnRa08HQvo
0pXgd85h3oiuhTtRHPAltSXsFBkGf913eHoRP4tug9GQ+gu9zlWyheJ5ygoFOKdk
rjb2qUke+thMJVdfmFwjlptTHQengACVXecsdOHgMvq8Hcp7HNWWeLby9OHvvjwF
tfdAMF7IrFZiJwEfgC4wv6+eNHBT0xg4KJ7JdcQ86WqgmZyxx5ntCuwr3RDsEea0
kJho37lPoxfWcDkrOl9J2/Z+WDWZ0ueEr7a66mB7ReOP8AJl45dGMSeUgOPty3/k
flr20vveGc7h/lVk2iboPSe5HTjZnkp+LLdLn6yTpEB+d+R9CXc+gWJKYg87yQMl
A9tiXe58ls+Ms4CZZAj5tJKNPysbbNgSNFBB94hC0DQZyJzLanJYpmfHPOURfPiK
WIx3yBYNLwWwSI7yRjlkVNvDjP3buzShjS6XEiTdV+pJ6cXfyLfGaKWYjc9gF/Uf
vMtphoAX97gKDBU70Jp1ZtVDwnmymRdKcixnQ+DF0VkdydFJz7KJv2tXFikSelVF
PhdC8GWRVIHRfN/vp1wl9fOfPz5NkcxXxtP59veRXBX+hXsEyl5g96cZRvXsH0EA
0agmMSij4Ld8vnJYuoZVqRPRLDtSbbr/pX5aLL43ugFnfRE3adrReF8e3+W1Irj+
MurqcHnt9hIKV9W4kPiTFImEiydmmPxRhHkzzTLTrrwpw+Gne9VmznehaTZFeX7t
/bnAPys+s5F+nqPtOpvfa4uc7CofkTFtELAOJMOGrEDboUkgQfTF/zwwf2IAzc2d
tVIl7NnY+uxPHpRTyLXEm++4INAY5xYRVNIvDUwxzBa7QvJIXywZKJzY4ewlDAsn
wqYUuL5pouDNiAUgrkjLqi2TIm83c+oATZQWMaw4OuKgL+AcAnRWPD+LUyJvsaNB
icL0rw9tstjs1j4UMamBX7qXfi9rJuxF4xbqRuyn5v+WlpJTj8HVmysUb6bfoJFD
EmuBMcUJCO5qnqeT24boVRAawx/lRLcBeeYc91hKg6dmuElYBY8txsFExD1rzJE1
G9p3pTzFhP6TmcPsyOPVAMeuP0Q/I5lfhkPQDteXG2fp9eDLiQqbFq4nYsfMaZ+a
Qu71/+pNscE2QYtcQ2XtcvoYApxAktAPr3Ir8XGBprtH9TUrz3UGaijDamrQL+i0
mFxebyfhioF4reOjmiKzA7coszs/Puc0Dv2oL6X6O//2b5qVpYLfX5o198kZvhMT
TqSOdqj4wXhpZh1CiWr2wC89kM02cBpoWvYtw6eFOiCd2J5YIT7MoiSgKAKOvnX3
BF1mN6lFdf+mk0QPgdY1KwZdSS25Pcoi7cb8KWs2/6nL/jeeUQL5vJPBuFmJtUhl
LJEZKWFbx+g8UMryRByk4bDls28VNqDJg8tN2GjRP/FEA9qdGq7gP7ivWw9ByPft
SHRrQXzH7lbmELQZ42DScnp6Cl6xK038HtotOzSVs9RmhxiJa03CH8RMf/gPEFrT
ikh+69FTQQTQjGH+8XZ2KDy0tJaXaXOVT9JZnKE16EX5JcEtSpnU4q9RDDfnUSsF
YkrfeuMK1TGUo+V12eYxbJnjve/FdwSmq/Lb3ltgql+5/LCyNsyfIWLNxJ2ndazw
EtkjGlCiJtBgL/02x3r/XUOvFQdGxdXC8Qtf0+b8YSPjgqa3VemqnVMltQL0xmOU
2f+nGsRWu5wERUplE+hd9DeMWE7j30iNXmM1VP9wAoh71tdF0DlRA6iDCmMxQT+7
kvqYMxXohYGsLHpwnvkV8pfMCtkUjtm51MAH2TVF1xBRqQBCRQ7pI7Pm+7MSXspF
foiEgUsJyxre1tKqWzBhUDjwrL6yei4n0TT/JVgFvYPH9VUaWUdJN5bd/Z3jpOaL
8eZuB5ip72oBT3I5lpAr+ByQoMttVNISCIqy5YKXBTQR8x05lzTkrRrvfe0FsH45
Fkhw85Gag7SNIx6C4nriwS+wsSrAyDNQZK1PQYHSgTN/1v4M3ag2ZBuaHp6VTeUA
x1KYzPH215zsnfqLt0lYQ3gWECZhktsvCRzcU5GRfMPFQQwnNsmI5R6lZi+SYGmZ
kBE13J/IQJGGpKk7p3+e9itcu16DJmZ8J9BiI/gjJvcJfXZBzWX+x5KrXSsgEPv5
XOfCOX79hBuRE1qBOTH1m/mZVgQt9PyJF/5y+Jzbju4Hg8Y998WwQxixcKX8F7Ru
0gc7eJdu8VR6c10jymfPTQo3phJVsmhoxRpEfK5HjYZdCOa7JkvA57JPBUMe3jWq
+RoLVcj9dKJxQhnaCn8dDUom8PinP1+MyXNq6t8f4TDgNQ83rVq1Q8jEG/htM2uB
rdFwjNNB59txwHNq9l2Cf2OzLavfp3z052NNjn/6sVcHDcelfrMpnAJ4x7jvX7Ur
BBJ9qXWmWedrbK4G1kk8cC4z1snxdWh0QRue7ghkdyp2PgxqEHs3P09jRxVAHKIr
KxcergG+zMg10x/AIfVWuOsls/HGhNedi5ngrNDItXCDloJ+vLd8+8fzrUIJWVj9
wUpjWmdBkOjR/SKCCNr20rfKufDXKHzHzCwyh+LuP+9Zx0D78IypLxi9+VC2DdaY
Rup8B00MVUasBBd9aVYDHZXkNfaJy6ebtMGhM/fNGfmIUMmmgA52E22DzncwxyQq
E+/fa4AbPbEo0ZUx8TyUK6eJdcKnuM1BsB7Cu+mXGJU7HCw6SXZg0zdhWi0CmSkH
HaJdhhLqiWpD3URrqEtBZMT0BLBKcvedZHDiX4thNsj0ej8ightAziPPZNG4M4Xx
z1D849KLNH8g9kOXasaytFaj5YabFs+IRd7sGFqzrRsvMDwCKtvXy48OxksewxLV
BqFx5eKGB0QdC4nJWI2cAA0dxXBJfu9JFPz2Lt/ocW0q+1Ch4Jt6V2FJG9+uje/o
mgALhn5SvxwjxFxVqWgB4W+gtPKlL4RY+Fu10RHUpatok4zYctslKFpFZShaflCf
dkXCWsR2kfysOdONXvyRVVzFG/Y9y/1E3VA5S6XAWrFXYpwSmW3xxMDhTE7Gs/wz
OfG3QymIlkfaNjm34Y78bfmIe+8/XjhXIA4557VuXPEPOKE8kG1JRoNCtVdTsbZa
KRHc8vK93ew/xc/mITjHIr7b/jYXdB1C1qtxfrFTfteUqgbC00n79Pvd7JvCqhB+
LWbohWM06IcxOuoFWTr+C56kol44uYadmliFlW2nYFzF0iO9fp89Gf0fbErjSWxn
Mbuq3WmSS27OK6nQLvb8f3SLWQMkXb8s0N95UfXdJqziE0JCuN0J0D5LPD2BfURH
FNibdKL8auFAvuFWxCXtM1kZKf6OmL/ny+Ft30TCACt93I5CQ+IJO075CgqPrBC9
b3u9ZUiLYDpUKJKTKF4F+gfLQukQWp3904YQUnkSpURqapC0z7IKVKr+BAoYLMYE
jx3H8mTnItWL5K4+k17EhsXek6LgVmylOhEKo4ZUvHRNywOd/rCJo6ys0hQvTK/6
GwPDPV8gj+FpUsed93quOdnYHdo1VVAT79251Qv1jz1rphSFyduA2g9ua5t7m89y
UgQn8Mg4UGSiJzxHRgfwDnnSI1O3Sp4fPVgh/nCrX1jYlhABjvKhpQFG5blsbgre
u6flqCEy1BiIyDEZv6zMXXSNcA/Z6WF90UiaA2rdPwPM/Kq1OiZgbQB/RsjzWwX6
uWpSeG/D/tI/R1P0Ggzitzzsxz2cJ7CvT74s8mbJ16y7vS6nC8OS5QM66Wi8R8rq
cO0irEOfafo2XdRyf/q09qp81xPrQESzNmzaUfFM+00+Ge2ipWszgwCe+H518LgX
AvKDZko2v5/vmBnII2Rt0lEX7gRJC/GwC8kIrvgSNAotorb9V2fCaynCnDVPFvF5
0UYoz1/mRlNh/SmoCY9rtZRjo+l7RTFSQPqw8A64OGrcX/RnyJA2wGMUc1g5OErs
8OUzbi5xKDB7p4HWi+yWA4boLSLtXHSq3xDNQaCFodKkcu9kVBQbVITaR+Yo2sK5
moH4EbUoE6Z/LA158IepYCji/Ed4TzkbprU+ue97aGnIfkoRDAhh5fCDrx/nncaZ
cvNHUKAtrcrO/7DqzfpbbLmA1ceYo3oNgBSWqEq5YphrI0GV9rw1Ci+xkhbCk8SP
Q5lsbJA8T7fh+ai9ggljlnsLWFSQWLCxWVS72fBGxhArdmMezaTrRQW+pUUFIPLn
C+SfmhQEVY6+jJLETHuIjfA3s6Y2bfSly0xWoliwNxuje0R25sKu6uuu1fowHNEq
0eQZBhDy07h+KTEb71c+kZ7tbdCbxALkKkQhUQ1sTISBdRxQ68AvhT/8WvmjYf+W
3GnxfaEoGR0teJlY35q/FPTlpwaR24n5XbMI+XzrkOH2X7E/s/AwRxbnfjLooFkK
5s1jQ4T2BUEagWKxxD0dUSdhV+u7IxbrndcA4T0Jl7XNYPUBfYJUGYa3+L3s4Uyk
ed6usHKuhKi9hnFy22wtA4oorhldJxiaZlX8q5MQpvH+TFZUZ7rgaLlI8MTg+n9g
KlJ5XBTviWeX6DnSx33zhl05/IDOZM0cuzPZLiDgG7Znc5SeZK8h6F9xUhYlCTLy
ivlE8tUkArlMsnEBhJNlBp5frYeeGM73obwg2GsHSo8BqfIuF9/wNIwKdTPDRckc
DaoFG6w12ONRExvDLuEphTvCf4TBpcDFfRYtic//0xSqyX+zblw2AMZhaakbgsdf
UCLAk1gBx4scMrIOeuij7cAhxmdhoIdYuR4IV8lcYq+2VC09XbAdFmKAOFMYq+iz
vi5VXeLRkoQdY3Hh2QlTgVk5YtvNfUAcybqOUcaZhts4p5pKGu+AFURWZ76NHZZy
0h7Fr4UQ8/mC6llp5CllvsrV5n+Ih54g/Pyg1Zgib6nhIbTPfMQ9fAUkKfBQGUHU
ATtMovJOre45PzABwFSLNh2vvlkGun+vz5Qpr2k4HUzkCkGjwTCMIkGUWwmO2gFF
p5t+oWI34Al2F8Q4ZYsopqK3pvEBqXzhWiC2DTjUi4w/TZleOQWJHRsAbbOuP49t
534XQ/75hi7kzsp0F7BOUGTBldUn7jNijRl91FrnPterS7Gneq813gXjXkjUg08a
xY7p0pLZSzQ0VtU99GGfPVe00K/kRb9mYbRUE1WiKe/dpCJarypKUyHd5Jy0Ybyx
veEJ93AKxf8/D7vp9p5DFXh2sIW9izXvVncY4xCPnQ4juoImXfEzZEzjfaQsevNx
TUSfBjyMp3/fddzprPzEOWcteMykHaTGuA48blnNMCFH3HVhS3oSKpBGyWou3mBe
+Dl3Nnt81gW95ZQI/wTgeToXW9P8LqaKraiJnwXoAC6xkKn3S5ZtdAHvvfILcJXz
rHohMol5ire/2RxWp/J71xeoNnmTBWDFa6T/th80Se1MPw9nEFJDbpyW2G1H/E1x
UqXGtY/4pSxCvHEJ406rWA0llyJp8M3kqNCqrNBteccGtqQhIdSN8nHkZCv2Pq6R
talY8wlOcXhfW2RBf4yR3up/nEg0XU9ZC+fqxGTSHQxcvtEP6grsx8enQNfmWQVT
cOw48nC0NI8u4AP3IA1K5ZivtRArBpccYeSIpME6c0kIDLC/WaQoS/Dh2rRdmp1w
PPct51Z2FCrkz1u38t+mcrNE0aMXsFC+Qor6y6aV9pLRJBtla6MJQY0qcNiMDcZh
qmHZviRaGfPkayedmKnNUALBhQC2b4zCfKVT4s+8QlDwD87DizmR89v634B0l7TQ
5pGwt/NdZKNIa850y5uNfjPFbS+cUQtVPbH8yjyTyUWJMa8xgJi/GN9cZmmymMGP
4/ey+8J2cFYe3B5QmY2vKdd3YZ+MmSpvrnPdT9Eg9tvEO8ub9mo4Cm7JMAo55+2P
fNsqf1AggBAQQ1LjKozUqEK1n7VxDCsrD1gXSfMl+YoC9/6xbxQaBI7A1AjPb2Lp
mJIuOUEweMVquXQjv6ZZdz50XOsa5jJjxO2am70xxFNuT4RhnDeoqRl5oUD4Nezt
9uXvjKQaYXkXBPuXnl1lVv+epfMUJjOFHu0jk/ZdPUyVIMmCw+QdtHZ6y1jjAQoh
fS2ft1khWzvFzljkUuGiCSw+xK8v2NbK/iYSdnnxefAiMQDlc6RybRHnsz4YZo0f
MAmcjEV1R5JfdepF86t5NNlfI+AUGAa0ECQcSRyhJoSIGvkpLBtrZo6yDlVE+5F2
5hFudZ9eUMtvU6eFIpoc5QMwn+SkzJNgw16LsRJVfFHO/UHIIV7chEjXYcltan/F
YankiRlP5/ChYiwZwXk0z2cN1LUDwBt3e9N0XplGzXW076mkbDLzd2345Y1ETOyZ
W//tuwCPgaTQPhoOhk6QMUtSFn7+Y8r2AqITGcqC03EKbYDsgvnrRoAi2IJ1s6uP
owTl0zPUtd70BH8cyOTMudebR8W3xgpVCn2qei4vcSi1D2hF45CS7hDV7U3c6/C+
bMf+nHo57Y47lCFlJrnjxqF2qAxJ55itvUl2kCeV7Vruj9r2cewGQL55QQrE+kKU
LIRb5aAYrjqJzv63+EqsaWlEkLjZiVtK0UklxADRxIxHPBzk+OB1tSwgkcdTzkxB
bZIVKHSdgcCNMgE90J25PjOQqSkUlw1LlvecBZA/GJzMWKEAcfvvlgDtAF7hGmLJ
MVj15gOIMqZmqegIypz7cJkDr8I6KgQi7q9tMewSAgjKBQlAhNNtILwxO+9Vp320
sByIRsPgoqT+4zbruQkLP+T5rfTZ55k0bd/ljutsP/MWMLbqwVaxrvnCoMqsBWYt
sFsX81WA3r67U0sWhcVHmI2gqvS+0LARrLBQ3nb2dpftfn+ZkXeUGnhCnK0lFyj0
ocOaqs71RanFb8EpSJKePvMc4MsbRDJsxOtNleojyQ7Eb1w9VzsAg14ap3Fy95HR
bivsr0f1qdua0clBNu6lhFWIof7aDDxiqSuXfYu5xlu+1xMrSYfzNuvIo+MjNAvI
lRLc9CyXmanh/+xLmZv4WvioxTjM+xZd3MbdS5k0c6qcY0Ja3fLFrvtFQOS+cYJC
WdpJXICm3UqfHqmMs4Epfym50m4AndeFdzU9hTsprlJEd6lNw4TJGAUZHpC9PRta
dsQR6jpQ7f/gyu1/0X4uj0o0RTKKEIwfEIkwIgXdi2oHNKc3/KuCYPdqCPRIkoON
uyl4b0gAZkVieVxp6XL5bKrLPKNwKbeIz4H/2A2IqVlsuyQHu8mIzmfELeY4ntS/
u+/YV/wBw5T2b+YiMznPmtvpeUwxRrB1yvTmzivcXTIKYtg1K0TEefzdHc0kZgAS
Pr+xljdCHjg79/umdm1pyo26Oki8skPq89rH85GyBTZTZezcnG7XETqB1igKnwpU
J98jb9vWjWoqV/AK/atBlIWWOjfOCPJTxRWXZ4uZnwrFWAZCztQiZaLNydNgguV3
WG8VLmtK9PxNciXiOA75DwmeDS6PZZ9/PTtk43bxRMjIpTA+B7UOV3PECI45oqSA
JIXwUsGikme+9o4YnQ2WiHqlRkbI191SLQtTaXOWchkb2UAr4iPNe01sUHka/QcR
FGVUiuVdmMiu/+znrFa6UPK9obA9FGUT6S3LqA9HeDc+uSXL5ttVLrQ6T8mr3jTX
6hkQg/tfF01688T3QpMV2s70H6FinWoO/NPbXFkntux4PU3vCqWLkitz9I+yDe8M
omBTp/jlXKXWBB891gBAfFXJDpWPpeAAdFH8anxvbY09wDIxuIQ3hlKLed2ThkMH
rk7PPrMZ/Ca5tCNycXwx9RgVR0Sbz4HcdFiO7304ih4XF6Rc/l2xPHBsR6xGy/v7
vg4hPWOtggmy6V+aPCyM1BGc1UXJITbHG+/03+60EyFQuy1VcDS38TPHkp7b2kmg
23PHfWForrRdadgHh7tyGZ1Yd0O1415gBfarHT+AObugWodouejgg2re5JbARki4
U1lbHPVEAdUxAPjMcdU7CC/jCi7AwdDEEVdAYpq2wlTtTws719zTohRQsG/BFmg9
gihkUVlCQMyDomjtpPcmisp6cVh4wNXfhT3w+Pnp7ZQqSXMrL6YuGQtw/wLqLxw9
K3e7Xpd8IgqN9rCBOzmC5/MfAbl0qId+IsEfaQf63DSuHhUaZ5QJJcD7sZOLKM9u
U294bwZNT+K50aUMTejaMdnev9HjTgotmrzX78Q8BYmxiRruLy5rt93Sl0gSZI/w
bsipe+5QIpd//qvHm8CISVf+ohbyFaiYE21bqW1AA5fsSi6BZHKXbxZQ/YWTlYV+
od0GP3GJ/JU/9AAZQNBUATycCtBpuKXk09+3Io3BBhKzJJqPp5Iz4/ikkYQDL/iQ
KcuvqQw+MiQYvTW2+yMvp5omF51KQVyzZ+wBLa9VmzHQIf1CxwootcyVmhB1mBu6
6/C2q6rYyE3wQFRx2mtFGtCXczIiP+/e8D4Run0KX6X7/8x0DC+h1S32KwoVo7jm
5e9d5Icg15miHLtVf3LwUxJnWdnNtSJxLMgA6mkHtuhu/srutn7jceInunOxP0wv
iGqNEMqsoDYyKldcTTp8piCwSy5S02870cvFw0qa6hOEUi6vFcJBZj1w9fuc3BR1
F4GVcFXJVEsAf/9TQ+6agIV+/x+QOQGbPB4WZWMANsYXgEpf4cFURQYA0tVmr3n1
KlAPjG2jeUXl+eSmicVxGXrB0b2QfAlJOaYVTz9Td2QwqUTUMVdVlxJPl/syqdOM
I4Rmk0vACtFsD8akRORxHIe7cdLeX7fTwfS/gPVtsfM+Z0Usgmz88CmVTDdbh8Vz
+jJbhH+Ln3gWavNXUT6ySQIQHDXQ8N755q+MC20Fik5GYEKmry9qcFMmKMlntFTQ
M/I2DCHryTEzgVIhztg5F02nZqCWoejzHe82Aw3ti0pQKmDcv5dQvwoTq8g47Vs7
0Lyktbryb5pnYpQMukGOY+8inGfc1lDnMnOn42gexgHMLWOOJIqXUqvXFwfHdQXO
usIzI2D9miNXF+kgNA4QVpylgPpY2Ok3Mz/4xb+JM9EvbrdfrE8v/qDDrBljakM6
yvzvMwzoRDXXFkrBhbwqwz0aWHL6UdVhlY/HsgNda2lO/XUvfUgnAKrwdARKgWwt
Xb8M0eaYlIRmiAXUdZMm8AP20sxQ1y6kfALgxEaba5alYgUINwGIxBGI5jM1FqrM
ToO7hS3QFYQqtqT2KLdLnRIXT8UTHJFhjJrgupcqgM8W6GD+/Z6KT5R8fo4zcY99
O33xlMNhwpNTshkbeVdvhG+TWPF9jxcdapPZ0BQ76azJU+DSKNBMu6NvLPM6hBWZ
HH01ok07DlpKN/Te2loc7YMkoGa85C9HFD8wYjn0dAXjKRIiBlaI2fqA4VhC0nEa
0omMGhbgdT77p/LHpJvKLJXfprXARbEd7rLROSIz3wTqHluMJk5zGQno8/mWTOKw
RbCNM2nJ8KOTEYnkg4clr/sd7dLspzMLZs44sp01wbKchLf9EJvI6SOgy7mCefL5
dOVUmIqdpO0qFFq/4kDJT1FTyjDcZzd7wCIyBkyWulJBmjscu+SV86XiZNjYtTJO
bmd/HFUQ1mO7EJD6BkLxsG9hF9ng3EVELVurkbY8nkltLcg36+pNj08v2avp7M9N
ku4WKtHH8bdxg6DemEuog2eDZFlmbKlQOOgokFh+4UxaytObSXOcL7a093o59xvp
ItWHjO9+1XE/ZPu/1qBavsKGuYY+w6M8uj9TxVzr2DoeUVo9HSowjEctuprd5GUa
GFJPZG06oibB0/ZG1laTFf0Sp1IBDWrAL4UFuVhOZcGi0+aWZhQBZldLvu91H2jw
PenRpGm2PVxOCWdoGUKLMBGxz7ALssH9TxKBgNjurjdLAAUlTWhNxl1qhHvJn2nI
cXRAOTG511D0chWn+uNIDVmBl3VKKhi+d0Kh5unhZwhGU04VbolncUk/hahs/h1l
io6wcD81zENK6uRmVaqcfnXnKDNJOr4osnZTkAvQFK8t54ZYu2LO40hXMSRzJUoE
Abg+JUgavXBt5jbWR1QAEvWqMoPZZSoWHiikUPnjb5SINXszypURa7GUG21zSMgg
mV5T8xVTzHtRRSY112Zh9d7Uu/fEETqQqNwWdgK8OTEkIppsfC4n4He8rI9hv+J0
LPY9HDuBesBfLs6KeyAvVfpjTVvUmP2W2cRKBwVDZadfWdoPpKLWk4G/0Z+lOOtY
tHyv12Oosxuv7aZgi+gY68Inn1vB+8Axh1rOTYBUJwWlwwa1QOb9oPsPZFMWQFVP
3VhDZFHDqopUDAovaoWRPP6XxlxsBUydxbnJ4p57+7XaV3AXWlKorBHH4qN8LHB6
nECBkAGgXxu1dczOWr7Sd6pPgj1u5P3bRAvjCshj2/5KJhr9T5pfWB41xnmXE9p9
XiLPqF1NJXPmwnFr2BoPuW3guEWW19YxoRzj91Ee/cxSDfHVl9bpXe/fWQX9FA5E
Qejj9z4W5caKt3gjem332gW73UqaewU8fFlLEe6fHgqhUFMytBRcX4YRJFUiyWyg
CLMMFcl83h/HaiAgXC1wtyGZd5srAVwiq/syWpzb9Aq+20wVx6ColxhzJ1cX8oSI
ysI6cXgn8BIS4cRlLIzEWxRg+sRglyoVE3jJSZ/2sa3ml7/rTdYBI7/0trqcTR09
DzWBfdp586hYJ8MpZ3E7M1QdVyvUl7MDrT8mzSJYtPnKSQcsTZvrInRV7MYI+OmA
BAkKgk/Iv8Hfi4uOp8x6dBl6TdHCfIWw1HtF4DD8jFSH/v3PPKm6fpU4nHKV4aA/
2cL3JpRlbCbBP+VTmjuQ2llgcF2sZTEbEmg++xSoKjN5BJJRZ6TZJygd7Xv3HTgH
MF1I2TCvX4MA9iSmqwJxOQoI3YQGqMnZgoVYjnqy6BuzerM6Qh2PX8kgJEecHe09
WlxWkEo94mlA5q6l3n78/s/rKS0cOl5J7sQThK+dz2t5LCMh5oUEZwDfyCH79j9u
o7d4JI7kT8lViSLfAsziZHxBYPCyZIlf/yRVvvtMcfejSL2vyfgSXUoInRonjZKc
+cpMnHa8eOegUdfFzJUnZexeAzZf98IHUCr6QyFjsa8//DJa2ahqjj1sx2lLOtqT
rG9MKngjJMXgZhB3GqRMopeZe1G4XhAaDsbAGEva9gsCdf2ytrgi6WlkOlOdieb2
snFO03gsRla9ifEIQRMV8lKwlpTe62ppAcZm56k17+YUSToCyzetaBxDP2ZZMIk1
GXU8llaAF/9S1BBI+m2CjoTdpW8ySAX06XVhcpY/qpe1fwntYn2D5Fqr0qN6QCYs
iC4jE2KgX14EW1CCrTxW39mc5K8Rd2aW1TLjANHZiZxe/5SNDlf4w4KnBvyRcPJp
rZbnHQkB8K6T7qBf20HWBu7KzU0gVLKINU95kebN0ZjuTL7DTwhVEIbQEvge9fiq
G6h0ghTy4crm8x6MdNmECxo2HEkQkSnmvxVo/PqtXHiwh2Hbn7Z9Z10tZvqK6Idr
XpcIMXFVfBYfVM67PDKl714pYN2i4D8Q5ItBS6g8NKCUz9qJEnSqjGSt+3+RvXHK
90qhGVJpXnGuMeIQzKEpA4ZLHl5K37yjAFi0oczNljjw4tL9ENpj7CRSgm77vYkQ
tubPXSJ7C9J6pN5pS6CSz8cnm6CI7vNyXVZXqir3rBjftz8ck1J6+cB0A5ZV+K4j
bprg/Jl7axiw6sI6yYRtxx9T8+g3JLcDjYDMLinwChlMx/wmfUQLnxJ9BUW98kSF
M0NPXCnQ4n81aahl7lRDpNO2vGiMOl5sYWw3wUFcv/VrYthBZtaQetoLvChNoFZ8
b/7CGnCm1vc7lgGl6zK0alJa/xnedkVkwH8atxRjo6YqsCVqkGUbOTKImIdqLWqN
XZPVCF7QDYPQyiqeIUMYZxLFY70aWvbLzknndkwRrV0j0vx1n16SvTLteXTu5UAy
gicBzrXUmCvKz72rQzClo1250vCHvryXepwnJ2rwCg1m+2g8ELZ9YFBdzjkgn12D
Fk1xhYba1+UGezpc+Gw9x1XFTlC0+khUGu8XUCXbYUzdqqW7tMBdG0kJcsFAWrcT
8Y5Pyq8fhNcp/GsrUsq1uYO6DhuUXWne+boavk8ZalAICg+kgrJ975egYC/o44Pb
+u8HnOYTKWoHfTdSvUtgX49GyTqSy8NS0/74ovTuLPGUZsKvvqj4fGKn/PxVivsL
T4+tu+O/bv/41jIw07cQHv/42SVA1gow6avVrohvz7iI4MT3bNZoSsjFApLxzCoJ
4kxZkzTBkR/VaTBF442+xBK4ngf40JTXTNDhKH76OBiY1wseRItnlJV41ZZrBI4Z
QUesBTVo/OArBvdggrBDuSqezwRib6sTrmuN5gXg4jvpLESuIkgnpsO51yx7oX/I
X2YmxXRAYrLeQyWXOW8SS1FYbubsYA9YPAIh+Eu3jNqarqM27QIn6ZmkqQzbZZY2
rOD7rI0IV5nbrcD7rLSRlA0+hm1Q19NcScU+LND/Zwy/DTu+iruVam06TkFPhvne
29es63/S6prkaXs0FVdapOcJWfAjDjf0x9nYhPvOADUa2d0NEkO0vXDCWDfzGahy
/Hrkze0RGu3W7Hezp9W8/YFGJYbtE+7DQFniByyuOjRNs/QhLUupFUXFTN1Tr9ah
EXHAETTE+AptZNqYbaZq/ptIpKEhaQVcQ8V6kyw8g0qfEGBCQ/CUbqGDYy8Nx1e5
mAz/6pLzap9U2Ys3QFDU/ySFlTFfyodKpyMBonNXghwkesXotnYyb+madTJZITAZ
dWzXPti3kCC1KIFNmySVSjvX5cimF4sMacFOo7aeivZCne9Nm+yZ5GzT6U1ePf6g
ifbX61NBIgtLuXKpoTi98ZRLN1SHe/GIytTy7SJdG/Nnrg+M8tST4GivSGA4g8iF
vIlspHHcudqJdY0yUrnJ91mRBbV7dQ9yGDf/Q09AnFt6GqVlOhGVdiGZ1Zb4BlMg
R90iaOG+2EEjSGWF6XjZHybj9T/n2RAXlf/BjD3Z05kIfjT/1n2yJ9KAnnpH2zhi
qoCFKpO9BkMheNkq5PBKTfUfUHPlgacKm4BaX8HBqwhFj2WMjQZJ630XAZmCbr6I
3R4z1bIQXFE1wKZ85Rd2+oq+9OdHjq6F7IuohKC8FUC8Cazyk2pM8Xgtlr/F3PDz
LWzCFUZFRNelsSRsOcmXZg41KPBvmp5Th53ec1C2doPA4V+jCj1+b4hLS2Pc1Evs
mm1TmgvTiXrqLCyxGGJ04EvF9/Bjjyvna8x9UjUlwD2Mi2rJ/hXlTzWxCZPFMi3h
szi16ewrDuWKsk+08BT6JZCITNZzw1aH61Ih0HQS3rAbc+ArPiTd4VtThdodtuyO
nfY4HX9bfybs8yYozQwv9h+j4Cox0YjsTRmHHfnzHHCpquoQGM76GD2qP4AbKsHE
AYaLpfXqWuC9eh5nGLyKvV6OTf+ttAD5xRR4NmZg0HR3odbG/f7jLVKeHAHv7hTl
GmhE7Z6b6L2Jw1yTbsKYcVxX8FXOg9HrySMvDQttEx1CXagYOnibHlwn8wIIEpqR
ZAZIebBWzZy8ApethmNC601I3G0kpRfiEQsZx6/7WueniO2PGtz5glzAFWVQt77X
P3VNlhkIu9/hhEBNmXAIEJ7tFn91vd/z0X4VwYE/6M3ska3tYlFV9/YyDcz9fSsK
pq7jkjYc0SaNKCaM6HLfAVfnbsPeZO6rJw+jt8Liygjk8mjk+gpMZdwYPCBcelv9
M0L3/x+3xy7b0O6ELeUu7Y9kgQ4LxL9Q3bUbV8jL/rqOGdMhRqitDou0aRLXjtud
90pS58ouR+EP36hpLeVc5cV31LPXU7kFTf77qrkF/5Bfr//qXRmgKDU7uRvaUORo
aNF7Mfsl4dbJ8KTM8++1Jt71mD5Pqdb0XcY3bYdqU2JBWqO/MiuEc26lAJhzHfy9
og4sKfnkbOpLz2CVV2IjXlqpPrKbBj7Db6cLqfAac8FqJqsPv3nwyFroVBhFLx5h
6s8QEfr8qajYekYAm3QO6HAJXVdrxn7Y+mLfhqCHKrxs+n7r4SunuHMfMHm0sCSC
MjD/5317H1iW2hW0OShSJYjjAtrvgOWKyf0vK478ZtPM5LbWBwc5LbHpTLcEOUoZ
ZcD7DE58Bc+elzVtbjFaKAkY3zVR0K9P7NRU2jTYysj9r+nuzjSm7gAv060IeyLq
aBAKgaFhvwQYmahBLbRVBGgtSWat/tgZOaxzvEzAv7Yy2fHnmDnjTwHO/dL30eQA
MY2BtI5uee2pcQK3IrQs4OHZusy80AaPHy/LMkxEEaf82m5NALP2JQU2bjvG19Vh
qvbMnaanx/xe3lWO0LROrcFFVdYXz8F7QGuO+mNCH1HpBJ8ElHEKj2XntYA0WZBJ
iVH41b48xcu5v8pDJn5GvhNjcVL6ydBCdWdCw/uJGtE6ScdX7CsRaNDD37qlsq3S
kw68iOlwwkk0J7uU7ib/ffk3Ag8bI9pIfUO2+Xmi4+Hes68tNI9hNeG4M83/9Vuu
B8QMeA+ZQWh2NOLOXpzGXnx2wRRTOavKZfP3XHJDxA1Ggb518zqFYAKoN1feNFoC
pln300/uvKvZ14Nt70/tZJZbtwaZ+pR2hYbr88lSLdKIuB6AwtRRzjdy+HQgK8wR
J/sAg1ODuOEfopbJysAqzegxOs0TeMOwXZYZwGF1IvMMVF2pI9q3/3KVnbp0MpPw
GrszuWd7eo+KqoO2Q61wpfcfUxB9Q689EnvEJoR90XLXSrFsIFR2j6jWukjQj5fG
6tB0D5dcTDnaYH4q9tz0TWaIEhve3WdqDfqGseLCqgfk7YP4jjAp1Kr9X7STddpE
ATe/OZp6M/mmFB0TEedyPDSCZhOM115Wcwi5UL6Ba4PorCiW32ZxVMuEbYbt6nEc
JaWrtJt96AjG4TNl/EuCdoyh0qBOnX+SD0CovLhKGb0B0sC7yk0qFiQfgazC6ako
aCl1djE8n7am1wba/uNSdjVGDz1qkN4ZckXj4u0SdkDMpPU4sHz8NcSogQp70BW2
2mVXDW+3frAvaNDnYZZu1dbV1lJyDOHWa8KR4fX2cCWeGbvhJYrWhFXHYPTs7hKT
fsnjeDflxIXWby+NmULZXCMrZHPtn91LAsWTxLxrRYuTVIArJwfPS6eFLiPeLJOL
zAanndDIJdPrqhNgnbe+khZsAddqUIAbhxLZ4jUW5kVJcLSBkH31sSaESEvpAMsE
KKRaCvxfQIC4YOw71FTk4aNJza8aMttZrtDT3dvZ+7lStLdP8yQVGBapwY1hydQp
TDcmbUUC0cE/eVzWTyaAGm1dhyEZKuSs5mgJtA/zUApiFDlv1nTd3ezzRkqWijoG
695gyrRZHcjYpY67kzEhGUvx21BDt666cRCBiZ33hQwDiEwXA8HhRALQE+tYTV5H
dPvtk4WQNJmETAOHhC1+zjE/Sn4hxGglNGxIXlyxTWiEJ1vQ0VesBqtpZF8tvfPP
5bNWuMWgbv6pnLHA1ULBGydVqoepvdy8EvGRivD1D9h+zC/wASK+KUBC8l5ClAWw
SHpqXFerWMDfGZHEYwGYqA9Hf1CmrjVv52nlp8aYZiHdqH1iVmGoQIxTdMVxMpvi
/iA3Z4fzh45Xo1ZGfGRJg9Qo9+ClZFPUr5i9FvuEug28b/Fr8abCQNInUcZOQAp0
/CjvzyT66OMtr/AqdHIw2bLBh82RUFyW6zmdweMuEW/YJ+9bjgADjHsmVbU86hxS
MQvUv4N76hbpafB099f4HM7uNgCJuzkFioykfjwM9fUvB3XRfqMmMYVDs1zlpxJ3
ZTW1ROZlR4fHst2nZWc1t920Dvyt2Ha120HSpT8+H2FlBjzc51WMhlyf5YAC8lzv
9LbSqxZDLUHsdY8qYpq+NCdsY/hA+jMIMqHS/dlnMxbVEZRaGGS6Xp5mGabjQyCY
PY+P62o+XUJzlr7GaH1SgdY9AzEKUK0+WUr4XzwYLiN2tS1dMqvC3ItlLdnQuxaX
vgtAaaEAGJb1Tw4znUkc/OHJsQUosKvO2lsqb6f/RT4WNpjJAPOuHwkvnGT8RnTU
ETaK9/Oa8b6Smrrihi2LNsR2aZiv47XvOUdO+KvbFbLtgBgH4QvCe0wAQXBAMSTO
SUkrr2IihVxjVeTPDndfYVT5V1Xdrx6/53wtkekZ7ey5K1M9sQqSEatjnus+Sm2N
e7KzCzDAwW6GOvoYltKvI4cflVh8GJiSTZgKzO42ePlyDItjRXsKmEUJlc6wHapD
EaIqJbb+yF54Yv+TlLtvjoXnQ4NFte8Wc6RmW+XaImUfBMAeu+L6QeK1lMNuaEwI
J1XUHJfQxofWrgH/j8wBQWOa7U26v/Ya4qyTu7ja1LD3XKvj1iQHFbLM+pQ0HkaB
VdAVGV2Il0x8ZOdOI3sj3sXD5E2OgyivyAGS3ECh1Sbtazvuot5rFIO9e22ufl/M
9k47hLqCk/KpWeHhtXmhjmtfE5KT554s2Vos4HGvqW/imWs44LydhcINA84ENpKh
yFjSbP1IVdE+UMKda9pOJiWIXPpEgoCZIfPLeNyskhcF7OcNGLI4Lz3EUyLfW36e
50wMZcukBMZSVMYDltPJymwpWQYB2DhwE4L8b4xcazAJi+JY8XUtarUPq+7SBNEY
oKzZ2HiWyPSdoplCW1r2+gc2SFzcvdDh+z+7ivxwaw7COUQeyjNKSGl68POFTkb8
mns/XAnqGI3lthM8PJuiPBKenITyNa2d1Ae1HetiUiXnVceYZ7cYijzsw6sKjqW4
kI1ex6i1xlcdQc7Xuujdhxw/d27YHN8eDCXTgpI26c6P99PpzaTNKs+4UILrOJWQ
g64zs3ymw2tTx4He8lu2rSOdhth9kxjBOaDyxaYiXrgvMY0pPH8TMLylEkw/4dFs
JwubEd1qiCMXcWUTvWQ2Ak6WV1KqKLzMo8CVIxjggsSIO8CGMDhyaVAE2sPSt6Ck
6YZUORdSjy98jyHB6/0dYBJEWQ0Z788s2h8wEB6flYVeeJyg/RpuZcSx0s7vwsOP
c3K661gIQm9iMjWM+C4t3Yax3FPfa0BVjXZv9dlC5I/dMyhQg49KbPi2QNoNCH82
S7MrtT0cbbcpC4XKYvCIK3twSkJ1fCltsGo9UnSbGGuvfocRp6NbVHABhXTjSA2q
StGtxAp4Pavc64FHIJlu3Fi7DIpM2wpT2zw+akb8nuK04vEMWqzVr9nKXF3/gpsC
I5HHVv1qAkFSLdHs0R2ikcQdJv4TZuCPCD5ygDKLTCsnft2uomre2xRukFW948OB
lRxseKG/zhzNz5WtO8LDdmiZC9NpkwXA7bJSdFrrcq1/SC5rYwGaYFLcUHdaUIWr
3iVf2mjQITq9GxpBeHm8vijFi4wTtsonQjDumqPFyuNc5dAr8FXnQBmqxynEZoV/
y8i33KrGE3UE6jiR9XxI/s8u+STmPNyziiEYdkPJtqkm2WaTWItBLPo5LMjHYnOO
ztipm7CUi2n7Oz5NQdeqjz1Rh7BSc/8vqLEZ3L02ChS4KBa2GydO+zG7f/WOdgEY
3tlR9mlx2kn7K1TiGM1xrBwRV322oyJYmVINqGtiHKCF4eviY3loNnHAAVLtKAj/
0mJv9XcTshPUAfNxVeF/6RqaPDd4IqzcbbEK2dC28GTWU39c/L+IWYN16gKtpda4
JWKxpmj3YEg9hvy6BM7lm0+57sUtScnnYjqK/OGCUVqo6PwM/Tr7FrhIHgwvGyTk
uCJ1dHx8wcHTAxfqlLIpmhfDD/SgICA8L92EIbVtjpCuvA9KVPuOBqr5I1hiTPkU
gsvwN1KiWMbHKrXlNWImC6+gz18L2zijjkgSY2593UIokgcdkqeKYWDqHpx21ERk
RlftE4ylzEZqBFRE9/W/JlARVpET9FGkmo3OzTKpOMiFca0WQQxh7+bEvKRerQ7H
tFmoI5lT37CYHManSrJsfwytq9cZqqDhmmiyvF+rLBFgA9RZqCnZ64QrNO1Bapd9
x37l5LISpxlDvshdrpz53n8J2a7QHoNh5zsgJdtOxVfCbKxU0GPrXTQDKmmH9Gu+
ekJESfhAFlqHq6KvPSL3h6ra4+LoPYgZet/2gzE+4DrVlrt8rPwZBc93Hg/iCgMY
s6A5fN4c4ANdqizLWsOe1ugLAk9xdKULk0iDnMKkNEq92ySYKLj2jj9l7To+OuvV
YeoIUxEgariT1rUOfMAS6NYFCpR7JPDWB7Va7A+mosuLRFcXRlsJibnTE0TEnqon
elKGnjSUjnNiaCUn1PYRx7ntcdfUI3SKpCyWCvDdF07tCkRdwEfPu746fWpHyBQL
LoZOIEtJGW94QF9xdv73ZX785hQXFa2ANVsgkBVqcwzVDD3b72KNWpkc+f9b/5CA
M3mz2N2slt4J7DMmC1xAbmKzUzFUSgIHqWpHdAM+DeNUIWtuL13P7+v9kyi/ePNv
tMRvbyyc6AqIfqgSCMp4lvhgF1eMCJcd4iBHgIiPWhlETcG5KuGN4LG5EOnTNxSm
f4Rx3UnqoBfis2e+tmwIwYU3wlCq82KUOvHO9YAo0mGKvInjenu//CIz9DOIJTWn
v1mOR5zFDOWwWhIbZYhfNDqtixdhE2sxYKeYAhFSxC5KasALfqDtXiAe7f7QjYtT
/cxp5Aoe93Wk1skFExgHyDNy5vg5yo9LKbsiFj5W78L7aze0RaH4NPTUp/1HszVt
OE8FACS0BLMPbFpxLPLqFrmZyAex0DufRz07M8Znn4OKUAedsqPF6nYbcddg///s
3TjYz6F18578chCqskE2sH7SthB4rQojXxHylsLLpvyEDxjLsd+9kN/HcaR/HOG3
MtLFUcT0WaAHc5qsygiotu77o0mCJqTBaFS1QNqWI0A5z1zjCXfEvYNoms7YrQs7
o4cCrx4Gme6bIm4+sUfu4kT0iIKvzl2xQYApsr/Y/agymYozEvuZPXtehgxcx5Fz
ZdZOsPbeQh7ngQ9OlWsYJsky9I40GMOf+38ZNE5zmWtBPZ/wyohfdBVeAUqJ1z00
WeUQuyKBftN1oBrCCIENvtb8RPsflMQhkmt7DFtdvwXOtBLloOiC7CxfCV0VT0kW
yDAHKBQCGFEX7Dj/UCbqo4hPvu1kuztcmnzDHuf7yc/x4DFn1iauudHhFaHs/qZC
NCbp8LFO4Z2Crlu4EodQDCNpHn5fLHOpaFfU0v76Chv2Cgs+kTgzZBoVTOOhhL1E
G7hQwU5m7KVSWKoF+cOydFGJ7u+utxhvToMJg7zq7kUBmilE+cuHv/qG2IoBPUtw
p2duFg3aGkDFA7QqduoAdQpqqpuRImto17xfF+U1SdNlNQyl8M5SJzq492PlG3C5
fohmSZWrNMO2OeGF4zMQaVJJWzkCLHu+hkAhuflLJM0JXK9kFi2M1OUv4UIk5OAG
ZY8EtfW42stfpTHYCc0wxn0DiYoAN2ksg1HtQdOX0qcMxYiyaYe+TdTbFDS01+Hf
TLa3XwOJvhjtpZjpaZhcaIRK/TAHWtsmCrbsFHgJN9lVcdY3VAQKetWEp2swN41U
MVjIGeScWOoi+j9xae4L39jmI2sxIeIphUO2+L3edqnMBIacOVL65cNe7U/PKwq2
87K/lsVT0r27HiOqGNH0uk4+Y/LasCR4nGl+BKj8a64FXuomOCBhQcyc8ZWzamdS
+ibtMPYPaX4Z7zoWgmstvMqkFJRohJ0RVPxbTXITgfJkeBuvAmUTwjrGe53ghoaa
hf6QFuiT5vxPJQVodGdNohxO5Ie9fQ1rYu2YhFZj1EThyN0nWnxezJFSVAXspvKo
LnwOKVmIBLQAhwdeLHEYto1cN5m1QFJJSHmjtsfk02bVwuk9pQNR6iKUsibE2DOI
ZmrgWLd5XrJnUXFLPT3xkQQ/q3t4D2CsptqDcWixfIV07MOPxtreaEvIkXOg6X6y
sSyH6wX5kacKCk6pPRd1buz2kuyPhdJrRcIt1VzpsBa8wQU5vduVSjiAXpPPsccD
IRWNZ7Xz6j5bCR2BUz9Zb2QeQ8mS2geoMIP+f5vwF1hPOfCRvrRQLiQMG5Q39RZu
dyyDiyk8eG2tBYGIHYbbHhSQKaohzIiELil/eMnEgWOkxVqbosqAaVYlxSA7HGbf
WG7e0+oD82AzFlqz9LRpZqZ2tdvdpIrlwzl4erCiPqcxjvC6FdgF+TQMw/TKxRsP
8oYOuGhSW/+hIWa8uKJc59bmwrrTQ4o/+9x8H4GFie2jhy596715FIsXRrhXZnzf
SNPHs1A1pb5pmfb02CAMQe5rvdi5rLN0ezgSeDZqo9vTaUafmuPWjadpc7xdHTLQ
JiCaewyXFCa2xsZVIGiA4h2T42yQS6ItlGPfUqFOYjCCkhraNF8TY+7g8p3nx0xY
wo1vjVMVrrgcl+bUbBPsqOKTbzc4B4sgw2m/xYTuoT9JyQTN/yTIDGP0vGFJh22e
+u0W0ncbUXCc0NDntW+uQrv28S9eByvR8hEig0AP3azmEYlG3ssOIuRYasxJzW+O
SFcsSf7jDGgO6ncWSLHsOxIb0mgQA2TJGLkSOjz3qfd8jdEUbRMkd6bTKPMP6IQo
V8gWrYsy3949NE3kJcLCuTF97qnKysyBJnBjqCcSpbpmGo5y7ApNFXW/wi0gFFJK
pKom7X+mMd7ayh2v9vbA+iJx16xZvudjFayexqzSPe0LHNAr+p5t5HHxFIEurprj
VRFX+aS0jVn24djcLLD38vWJgw+WyUtm8cOO6mkrrELVFHaaiuENzflvLQjH0oSh
rWDkYm38u5KeD6eNx7hwW1jeYoWi2pRIWtcvcMf3iUypS7lUwKEaYUMIQYYFC/Ye
3NKeQwkgI83aITdJ4NLCMKDFyi4jQfnRt/lHd4TrwABLWA/n1eCm/P09PkNad28l
WmoQR3Q5FfW8p237AUvvVAGrCeeYqgVpWeOGVCyvm7yuicDy8G/l3LC3LrHU2jGc
Eg2hH2GACXJtoTPhUYeFo8SRZ2U+HGRdqZQ1/wGwMmRhEKi35jl6lTJkAgfyGjXO
t5VMc22yi728eaCG9ylWCz2NeaTx1B/Im25MDdApt8FrnfyWYa90CQdMyvb4QnjF
qbIah9apZXz29tI3Dt6pWbyXxTOS54lqzN2ADrwAp0hCBPoDmcYUsYVrgdG8kDlM
Dh72m+ePKeQq5IS9Vz/E0IZqDN3ugO2SWAnN+Bqlx930OUD4tavHAaNjY/PjvRcX
6CoAHkEenmMXmUtBroGbbsDV8iglc0FkORLxQ72P0nEeBi1TiIes0jR9u28MLBYf
/AatGLxd6ZFl6o1aQ0WMs6P2hO2+XBJni/E1EsdABZuj6yAKZC2JfBi9Osjeiylm
fjDDfyIz8DDuJOUcXByUUEkYWYzl/FcwbQ7nfj2zGxJdxMGLraxUCN584mJ1jgKL
/BOpGIuDMjIZ0bCVSSZJQnV7KLxrT9cpfMHXc/KtOUcsVMm+BjL3HpsncCQk1NHi
oJiMe2dI55YnN/98arN9/lSz4mGB34nGRLr/zo3qehYvkUzOjW60OhhoerVRXoz8
9wy7/MeVd0xk8JpPbtsDKHGYAF/rDj564+PQTexX844Q8MbSukCjI4UnzQQH9Dix
pUP3cDWiPD6DTIF1pbR5wAGCnzXJc+ZG6DSyKYLHpeAgm/7NWfPdJGM/DG7iOhZk
n2B53eiEUgwu+/Ftjc94mYhWEzjjb5XuCs5Y8pweJpdIQtsmBTRbLEFZTcuPoNNM
Q190Uc4/w6nzXefDZBcU0g+YtLtIO6kdOU/rdAUopwcZWz3tIYjm1ztFggOvOByQ
eaK/4YZIfYJu/FjXPLDB6zzl9ZWwOnBzdTNNuOvo4kRNyj7zZbGM8asghYKVTUi4
wrr8L7Fbd3wD8moKi7vxRnZKwHhGWKd7tTai68/eTP/79K8g68/hjS942akPoIgN
GAOXJS4KQ2WU0z+RGav1tZemypqBSAXYelohXcOdtnvTqM/QPiJXIRVZS/wMc8PJ
fjlr01X9jrhv7tsn2HLwCqKu5ii6VfLA22nQ2S/ptn3YTfKvcOwborqhzIvdzVX/
E567/hiwKxqv+8PDzkBULN+t6pHD7kyh2VD6jrYQsBPUr/yZOJ/w9l5+/OBS0HHG
8FZdoBb6qocjL0L9GwLCcX3UdqM2tJml5d0KCPT15nAShoNWvWdmabD1fOHYkDMS
KhM7q5+l+uuvDfftpfa8GrNgfD8/md0NXXMm3hYy+EtmDyWxXIPzFIsV38awkBBD
hPzWoyGPEple5a4EutsAUg0pY9ZyafDiENFwZvGZaeAX110AHzPLo4VYhEH1F4wk
NhMUXqbhe/YzoF0WfhAYxTN9/4pthH8Q4PID5rtR56RSdVztpsnjK2yVxLDykp55
OEOmRABBuU81zfN02LTqzzBoPRD2YkVXtU1cGHrddI1Iek3BS4EQhtjiMNvreiAM
agh/1F8ikweFt7sWHrps7TKdtiGEwi4k5yIDXBAIJ5JNTC04wdW+WoL8JdbPk3hl
U2P10x/UPnt9MxFqTDuf+3griYdIQuNGSdENIXwRnwwYsE/rmJyGinTJwfxUHOO4
Ippsnrpqujf5Gl44RV8YO0sWGJzHpBrfFNqdG06pycbkZztb1hubhyoIqF5xEQUj
9QuavKADXiMEDrVBOHxgBPuJvQ5AxxSvSXp2TRNom4xKBKCqdzZkecYr+kQ/Ieo7
DNp2xG2TpQQfNi7rFLq8nOy8M5HTitjZOg3hMsYt6CCr45Uf0gnRx31A2VMu9gK/
NtsRkVwAyg/VZeUdGr1RA0JJEX+WJCTiWAReO36b4DoGm5EVNjMYYi8UukhDgTwW
O2unfTkd59ctjU8rYn4nnbJnVrxZsi341+LBOKroqzHRjWujHrMyoucF81cl7SOy
orhaxv9jY5eobzHK/jmSGaNx7UOZz39VkJhFN+7px7GzIQjWQULfTxb4vwVZpuDQ
kswTpoCdsHw8VR01d3hZCSQlvBhKC15Xq+MhCuII8uxuUChfKpNTtOmv+JIu3mLi
oPpVNm8zW7NOR72r//vsHAS5rS2dvZxj3yCNZwWvrdH80nui+/wVX/hG0HHslxoS
vZb+3ny8bgSUbNRd0McQkLCsXWlESu2+adbOekObnQx1xmZFmBdH9B9Vwu0VU5ZS
NZX+aatKRrxgDx3KW8Az577hq3QVBtZN4pMOVkKkEFvHh6Zz7Jbrur80yv8SdSxt
sdVzF/fTv1pf0AyUIFsBz0++x9OXAmGTGgZ9UGQ3KgtCwid/HitCMh5KX3ich6CC
IdI6GZV6HCxkjElVcD+QUjSkuy5++KF3od2WJug0xGSHEo79t5506P8sqIM8eA53
2PeE6aBddQa9qGY77yApnhTOnpp0UP32s5TmNukIhBvs0eXfjbXCJCLYQ4Q6I3aj
dSYyVeweAVM2Py8XW4axdnH0Zm4rSCG4/m06X/nUzx1K6RNlvsfEMnoKz4c6ST2r
dBc+HqB0rQv8cKiwn6cDmilRa2TRxeWXuD2yGQlbD7IuLzJuZD1cL4QDlb2JqMft
reJkI+R329qdKDzmzeCYksdghDk924ge58M5f34Ffbyq843+mDT096JAjgn5HfPH
x59o2XC1CJZ7+7YZty5mjBVxQMl58WNu4cVvJtF+7ij6xGyPEIf1rtwUF89jZWG7
G4lVU6xYB5l9g0Ls0IMit3HE6fw5OyK76skEgOySBBvqEHbsadeQloUC5XEzqdWI
Xt8yTPm/PKGdW8H0Br5TSu838JFBtzE8wy36ohqkQwOkvc6K6WbaP7gYWft7ReCX
H5ezYdj1PjgGN+jYjDutuTSlXAIMStxg9MR6ULnZxsmI/jWozUWcFfkjQEkNSvyj
LInsWhz5TRPTQBxI9Z91ZAa3/kbhop5bSuM85YerOFy9hM7AI6k8Qn73eljPVqyS
1cJOq2t4vKu7oSgLsp3kghPJs0ksTEt/lE19gmx3+5Aw0d4o9Tz11+gFCRibA5TZ
pJ4U9Ln1BhL7yTt4BbsOmHfckqfkEEbyblzJ4QX17eUdEJ35yCURcf2FO0NyTlEb
Tzql/xlnjLzdu8BYQ4IkeGSQWSJa2QF6LP4SS9B/6lyG4d745v91QI5+fiRBAGc4
u9oMJefOyKtLplEYtiYDvK79CmJ3EybZFRGM/1cBTXgGVmb5fZ/FPDh6x28AacCD
ji83GcOiXP6ESw22Ua4WbfrKRWtAguV/zUfeERthb/3v2ceN7RY4bd+nnU4VE4Dk
NnWzy8CXenFSJwcVyY6LswX4G5lCYK1LToDeS5JdukIaoX3Fa1i6cuaKDkiiPp2k
nBVIqKm/02SXgvKg35EerR1vZaCxSsb0x1ygjU4WlB1iAmQgXmBb4DK/OjE4lxMY
zBiEu3hG/jTa3fmHgRlK8lik1ozXPPbq7oH1E4h3KYRKAbedE+9c+DbSB32HQVVS
sNJ0ep0ks/iD4US5F8L9+MdJMJSDpyWYEp9BRlf/cG6sLzhqrkY/LcgN+FZDZ1Rw
kRYbTiD+tyfahag9DiXcfg4PjrxX2Fwx3jjfu3U+mGfC7i+1RcoJerJeJ4IXIXD7
wkltSVnx6DNWIN2jv/VMc0RA1y7uy1eiP6cBIoSBFYbPKl6ljsvov6yIJt6GfY9y
SDIQwgBzS/Xm+ZWCXAn4MvzZ5RxMDq4VFVSxV8Kkyi5Pz9wwZkBeINnZoYmYYuDM
ByFR8m5etrt7pHKNDSqU9Z7nO4xYwE5yWDC83Oc1nBZo2aTLpJgL1VL3SFcV3MaG
5Qj6ZymHNSibLQYfgmwABfPXhB1LoQSTRHpqkC7gpDLDcoy9pKk2JiIqY/WU6TSn
18on1dSOV7hIuDSEkt3Cy/9xAqrP+cvzTFMikekYo7VtvKB60xoCnmds1p43rziy
jgBZ5HjmNefV6c6AbS7xBlW82ojRKTawHWQQrqeKvp9ZE9ix8Vp90ve1/6bt8aMg
8kC7blpu1p6q7myT1MV+imZsSWdYrIzGMq9DoyE6YY7gCkXpDk+CF2b9XF41/GAm
MvPglHhuxs37vUnasvLgtjdQV/aPG16PVQLrotKoB6PrORi2n1mfRSBicq2LVccQ
csD1KD54mhOvHWcs+WchYtDPQn2YUB6mi7LRQJxv3CouMrl1jrs1Vkripsb4SR82
0LqkstODDJPYrD1QKjGXvtpAANbiXPCUpVDNK/qcXUT0YK74bBCXkmDPhA+oGzbA
IfZbfcp+m+sUJzla56mTYvSJQh3FBE6cT2+4QL84TCrPhwfNvGH/B4kgMNT8+g/D
msog+3XNobVL1gdxV+ONS/j9liQagg5PqZEEDgU7VYlkt/LATncJnjCNJIhoTx0e
n0DWiRsh+ukGbUQF/uZIhMV/3kKtF3QujSnFs8qOKnio/Xod2szYBXP+ySg3Kyry
h0HmX1L+w+nPsB9em6Jsn1uFJnZb2WN6pKFq0d0WJthTbrUQ6Q90Li0zmGq8Nwrc
kIE/SyrXyvjheeuF0OPILB7xLsdYsdTsXJF7hntgA/tRHQEu9XlShR/QHqeALSTA
3FoRKFdsq5t0/f42urrK8t0jS5UxG99JHzKFPYx6CtRoxnaXFgGqyiNFxvVRvGPd
iH+13aWsstTK2eFARJ7MbfHJBdSk5JJ7yyLpnTGzU0pOcMtEYLBjJ5nSZJO9T+jW
k0fr3Mxm83djQ2Zeqk8HM8+HNaR5P5ND6fBDxlFF+B1PsiGK2BHmwmzaGZ/SXo7i
eYFql00CjnZNKA/fRurk6xjlvothJIveQeHsVvzzUkpLtKrZNnCWFQldr7RbkViT
szhNDO2Tl1fwNBJQdGcFOaHx2faUHTxlXzGAdU3ibKn4k8ZE2GHRWTiiYQDuNK0H
J5Xv6X4sx8K2pRd8pdNPhvxB093m/gq+iLmulKB06oPgPg9kWwEtqqzHcirNw489
l8ch1hlWviJDjJPvi0kl9jajdIjhbHk2WoR13RMYURgs6D8LBE8Qz/Cgu722S3ej
F1HGhdxjCw8rpIG6sD7gXObKcUBpQPEMP2bauW8G+AmgAeNZd3FgTpN0Fj9HilZT
E3nwwjBpoFrE777v3LcV+XiaUFVMq9iHUSEbnsOD4lkVzD94akvYpG3d4l9kfcL0
rFpzNEkEDYvXkR0O+2O3BiG029e+GCF93b4nJqN+loMBAiiF1ZLMylsr+AVu3eW+
2qh8zteU0kq5DBwMOJxdq0ToG8E/ltmF4unPOYAgECmKpPCCvJEoQtAssgxn53RR
P7y4Nb9xYLOgGmCrV3ZQY+rvz9iIGMEgE0y6hxxydMdi83TSTmccvR/7boTouVvN
BAvsRkuajhf3YrqBoaXjUaDGKPknHBHe75XIZlc+fSYESO+TY/zFz9JxiYfohvhQ
8PQpWsx1aMydHtLLy0V6fub8ieY0mhJRy+ZUsm64sWMM3SCHdSOhmHPjorpmZOQl
ha0QPmj/uRJifRCMr4LNmL+3svvqhC/VgxlnQj0C1kdPkQ+g8fw5Javp7d5/YCd4
eP/JX3PbepM8gxV0skb8nFTczAiWO1QGWrc0wZv0rnUkkFqcHAa/jqe2MYIgj2Ck
WRB8hS6wIeLacqrEHMqshDCRXTwvwovO60T3wGANAmXDsrolhDOP5pGkKOunHFAb
hZGEOlVqQDxtP/AaoLhifeYvZ27ohWzcCrvAIiciNEHN+XcmWZJMVD/yuj2WvwhE
NQWaRrHlD6UZJfZpUy6zAyn0JyhLYy/WicahpwLJ6wQz85mw8j3XAhEOKkYFyfOO
tnkBGKNNDKF/J1GCFUq/Dp1B/YtwwsiZaloNpoja6CW930GKBq6QbrwSAMtq81aK
y9ivbD93thQFstDIlsVcsDgA5TU2a9SABs1JWJ+FYcajLIhvW9tV7pkjWYPyRmlG
wdswqHu384xCzqYGT9UMYkoGkPdB1krqrTGxcwsO6/W02EGQywkctj0LLgEVivxL
ScZx30uK+24sjYtiaLZQl2fagjm9AbeyCV4oJDZJauUiUPjGK5guda3U+SafaCUq
wcMJXLDA7DKuAXnehcObcHamiAvGbXNjPT7RwBS8CieFZTLGHwm53n2widAw8bdu
GKr0eR3hXngoaVaeea1rZZ9FA1wUVESs9tbMQFALNPlkZ5hO7PJ3NouyMdFiOpQS
yuh5eEI6Sl3rOmzslzRwmfBg533wXthC3fvRCUlKuoGNdr9grNF2IGez8ICzAOJ7
0J4QXzcSzkq+MJ6axDPJc8sZaDqvxlUQ2rnSOdwt2wwljn7Ts0gyAwsxIVS+gVq5
7ArNZwbIiJcR/mJro32c6/k4TyJZQGuCe0uij161/Ix388KpJP+M9W82ZUvzLR/p
Om3WFGBK3Q7gDGd12YISoO6Edz3L3uJ42rpLdHLulqfO0buRDVxH/eu0gMhjtizh
cA9Ln/mZ9RIxzF7M8rBTaRVvOTP3cp9zb+X6+esXJz7xDO9XpyyZD95a+rBaUyVm
Kmmd+MaOEA0k6pM3Nw8AlxQBRd9/7EVPzGkp6xd/wARV+gP1fHGcDPclpdywrt0g
pMip2/5UzwKx5PZ9BheRx5GqGBi8/m9DVkN0HO+y1Fmyb/ut6h6AZ9ocH/OAF3Sl
CtzdTzl24n85Y07aAGGQ0pEaHUCZMRcGEI078M0Pb+9lTzOJh0267wZ1KT2RaEqT
Opr3+fYbFX/1E1WyIwKMdHIRaG5kKDKu3QBmR8h8/yAhwgFH7wgG0Mck0ASzwjKh
FfU9BUm7kuVgp9rSfC1H6T/FwzCS5D6JQS4LOmc9WMjTtN2JyCEgLEWO0cDM7oE2
jS4D6vht5TYkhzBf/nlomAGH281mUzHzewaYPMdcMPM6SrsN8GvEVDS0igbv+3W1
0+/HJfYkGFwgPpOPPO3doBoPZ5TCE7YKGtu1T3mvhzrwCqgHKWBImM8s4PRsel4B
fHt3odNhszpNRQKf8ALeiFLoPAepyl5rUGuMcl8brb8wrwzxOwyhn1ydJBv8IpNs
rinCMbGVGuLhf9xvp/OWjq185YoWp4whT9FPWr8zu2Rv+uBgKDJ3aBsUfwBY3b11
UFjbQKaFm69P4Gy9cV9qiFShD/o2IYQ35yeMd/epQsNEtHJtofMUnlo/s2r+RRhp
vMLXbndA85aKhQWwtsShwgsiDWmPseVqUcjaykrSnpnKoypOkU1c513RG6qLy8W7
EqmjVnuG0LgIdEczdKKYFvxP1qMf9tqqB+4iFSaBGUvDG3uwXsJzA38ThjgGHMxZ
1DSy/esx1hFkM3c9t1VFW0LzdVG+9nRMcu36Ed8Qd777jvVqwg1WpIOa4YdSSLBr
8CMqAKtvSOc6878bBAY3Niep78O4FDjzcZriLGxmXURC11YqT5VL1MZG9w8QbX0H
rZBQCjjg8nX1jNerfxGxa/aNayTaUDIkA5mVZy8z+mXPO3b7ha7/mW2MGF1SvnGv
2VCZv2uHUD2TOfEpqA4i41qPh/UcPcL+ohxkP+AlT2tfdZ/ESPTWb3d4RNu/HqNX
Y+K0kZ+cuePA1GRuOPRm2IYLsZo/8qj+D4erKdxV5sRNz+IJaR7YnH7Djlx5Ds4p
M1NP8/oICKgOxNGT4E3rbPRNVYNVtqds8Cs5U2Kd+ChVv1lwzFeaQMW3Z/+PmXpG
JndNI7LSgLS+qBEMymmytVJj8x4F3HHwFuuYhpdCPeXI6UgxpfIpxDfDQ2k3jJC9
q8dCi6w98fSSLTIrJhHbsm7/sj1HaESV37mcGOA0Pq1v8rskLXA+3F3LC9HfNjVz
AXtWRRWxcuNze94VTsDYs1r734MXCqn1Wh27pgCMWL6fyvNi9B9cFuny+l6/JPgY
dVi0Iv6pFfbbPixE2MiBsAXNG0mqCFNnd5COZvx6kFhNEoqILzBtS/djDTLY22/B
Th0euT4S8nXluRGy6PJvTTQQljDgX5DCV8Ql/dGVA6jJV/UgxEVM9PcgjJ+rNshe
K28+E7pbJcG1qh+v6rc44n07W7PtjlfyR55GPNoMxDzlFCEOWoC0jj7QG/ObOZUI
/+qANefLowsQxkH+K6Bc3EjPXTztOgLDWnir0ryGMdztK42M1MuZ4Gc/UOlasuKZ
CJchRouNVroC+6W8ahAmvpwnhrkfzc1N7j+67kbwVuPzvB1nalfuNvdqdBQ9Of+4
8jlvNCPymgZj2FZXxh5BUy3LnVmavF28+JQT9VHRFmYOW8vqbXHGBzac0h4q2cOa
9LlH04QdJRbxGO+2S+pn0AZT4NEkmsijFKMJnkkzKHoHFiClRwL74YTpnqLaGIOz
bDiKduX63JFoNGzGGOc550gBUNgYgwAvMbF56iVOeer8BTDy3T9FQefqVI0snwNy
nvDZEa7krUY4rDRXpNRcBOSByVVFo2kSZJ1dj1k15LJKQRS/b46UGg/0CHglyqdI
G73G3EIiBgJwVIYu+8flMKiqmWCq6I1bQYNzKUAeI8Ibl8DBtq6pl720+2eRe4Eh
WnBUgI8Z1QnzDkdAkChozj8G8AeNphDFaJNRz2lc52wgPXpt4iB+tMAgeXMishrd
kG4vlLDEbcJA5HAvFZ+lFQYKtRGtTz4VdU0lMiFeJSXrXo6i+xToiRpqVK2ts1yy
rLYZLy+drQ7PCY1qLLCC7NDrgy2TcxSg9IEQK9fZRPs14Z86cZzt4vS7LKI9hFBp
jeSe0DDC2tliotxtxIFzmR07Ciu8ulGNSC3y4jI0YN5TJ05s6ARFPxbOQHi8WTLi
phC1D9Vl/hb9ZX5SVhjdeMHnYIyN3t3W8FjHid8/xuZyJuIAfDqtQj4G2DeGAiZP
cfGjpUWa/yUZs9S0CSoM0biJMCMFaHwa1KnL4+88tMH7Yy9Cg4qi5LLuFMqlFwza
2VR2USs6a5L2e2ED1LzIfG7kxZkF6GiLXDOEUuPDyuHwoAY9SiGjvaPiXGKv+Otg
TwDPQQ5lzUdokg3NAQyajLM3F3U276kK21Tx4drEeLb6dkaIF987n9V3qC+U9zkI
lf9WMpRWb4FhIIjUUxXFdMvAWzgGGXoEG78J6TtFETUEY5nMbWvqk/ntxzNN1uEV
oB7wdd+P2vIdFrbMs5wHUAdxyQwFo/QyahKPY4+rmSTnL9AxOxgn8TJYoWM50mIc
/EjqdM6Bnhn0u/0uH3ueVuROe6NvDu097g1ybyR9ojchYHKrq2hRTAfS7eeO5gI9
FaLVKE89LgGAntaasX5pPzliIZGqjtb951y2WjZcwO7iq3a/l+qjXbKmOrNDbdnz
HA24dM1suLn47G7Y9wfifTGrNubLOzAorfyzidz6xwcF5IAaMrzaPJiHANCH6wDu
jWtTe93lvjx2fwCbJ/ihOQ87uJa2MWM7/gHkVv1C5Q0bAJCN/Sd4+g5fPIdMbZv6
tQEvBCE0FarWv4hbnNA4Q7lfCPlQizFlwM8MfXpmtTH9FB8bbfWjJqy4pfEBKERZ
xVSXp8KyoQf7YONianeDs7WXx3qkk1CT8L5jaQyd1bIbddiSQqxHJgZrnZM/s9kj
fjYznsl4emtx7EHAVOF6JkFI5hcoKyPxoWv4h4nwRDc15TXW5CHGjbffhLN2+qeT
GHd/boGWSQ4Nf0FYkVpwe4SVEIvLV24GRkfyLg/OPLvTDX/9ZpPUC9eurady0U3g
4DymxrJBw6/e4N8x+qYBbRx/reJ+6dVLLNNzRLEjLWauT2VLG8FY3tTxt29N5t/E
UpXV9bQs1LJ8Vo0l8JtKV1Bg/Kd0T37djEW8lE7eK2vGKQTrXCZ0SRYlBrageOJG
7HOcjIdtrgsudsNyjhD3RofGWq39/ZVQgackKJ3Tx2J1RwYdaUwvC1thzpIKVlAH
TSQHjQToZQu99SpjHsFHwsEXDHAwi3y7d+gLmNvHgdh0z4UkOnpxY1172zzFI3yO
bpE5WHmkSPvvo3FmzHlLAd4PQDrWKayGxa5IyeodS+BG2mOPnAChTIwv7Ak2F4Rg
NWPok/RHgbM7FaPlaTaZ/gXiQuUa78dPQZv6bMVGNg8rpudXSN0a32PmhFwEhnZb
73CZ8e57uhWECWtO/C9bHnNs0aBzlpiKgpyPBM6o9c6aKpLEpSfbp6mqrWGB/Xax
PnFD59kRG59W1Kl/fDXVjgCbXTc5hv6ruTvGawIkt6RpBgtrvRs7Hc5PGdWPS261
qr1a/TfMy6J9QDuDEAq36Ggy7Xje2LiFPv0Z6ZI/bT8mX59jzSzSHx3vTE/0L9DG
rxYDVz/e06qbhAvuOEYpQZDmbULIq+BVA9RiHNIYc/dqwgBZHBksXPJnUsY0ai2s
KnEYIxvmNsD92ecLAqEIb+stKgOZ8WNqiGF96myIm8fMvvbIImlk0BdroRcZljqR
SS+OYuFc8cVrH45c7mEHDKVfkAyzP90bDelqZ9CGJpaEfa7wNJ6a/yC0T8fktN0v
gnMecxAz1yB226mErVZ+YZeboU9lWwTSQqda2lMPZpKy8k/Hb3URdBCtgHHQMa/J
17l1kZGo5UrFu1UpVjJFZURwh5kfyGPgplesyuuDPQ6yeWwfpgnv1j/DwEyyg5PU
TA7zKKG2a91bvQ7rG4lH5ozKJucLxb8ygX4gnH3wZGOphDSnj1a26xBJsXS6BkwY
8X9SSEz3MXUc1KKziBAPXYljoqc/F/Vq7VJRYXP5krGDF2qraf7Gd74QZJ/T/x7S
/VBxOy1770NboWI7lo3pwsihKzVDZKPptFwKnhz70InhxiOg/OsjRrWbCDN4U5tc
BWCSxvRHVSqSFE+XX9Z6Hj+SyKOjdwvRoKYiygxe8ZucbgSOETwDOQKYxTeu1Yk4
SJrrATKtMn99sDOgkess59mKmmix5n6/UGDyMCCk2Rc2BxZAIiX2EOb99t4XTjP9
3jNAz+3abXnBfcnsSxykn+LWKl3iY2luluFD08a+sT0qejyMp+QI1laG3/RJQWiA
MTmxxEJYvG3d74DKkPP32I0NzbXD9O3HQ8dxQk/8izQRz+uiU5RGKCplwb63MU53
w4jAGJkdVxp4om54ufe/HeoDp1s6mC2yix9bf5EkUa9SQMRglgblI1NawZA1GdcE
9B5A+oj68JZiUFH8qZldPWUn/LC9tevmiv4fTjv+ge+TPgsoZwpmblmFTXET/U4T
dS7PxigJeMaRAKfo76JHfac7aAeONg29MzByAL6Agf/e8J4cBUMmkrXL3l+pw8Da
UVV30GjkM92Jmj6scDW2uFM0GF0cUt6aYgJeKMWZslHP6JvUQqIiv7Ld8mXwj5OU
xChcEbVmCLIriCzAODOFH9TXINeaBa236RPLvq1rpVl3nIN7DRnhSTyjHj+XFh1v
DRX/Srls0G7NLxZDHPCioX98cXijaKK2p4DIa7eoqRsgQKGfw5oAKXfXoxtuVcvP
hdfpO+5ZGaSNM8aciXITfu3z3Vu+sfBQwZtjnxJ9IOHrgIFHc5EN4+hxaeVCGETn
vmS6tl6TY0mOiJuDFpNJyyzWY4hPHUtVqZM0Tk4J7DNoUUsAH1TDPOXyO8poI2u3
5ZzJXa6ipJ5tclAbaddAOm2kOjNYAAOUyvHJ07OorfNICdnRzFKfHcFXKPUrnpfb
ZLs7yz7fJf5S2rFeyThh4bzt9RhLQRcPZaK8ZGgv0AX4KGEXd8k8ONdJyZ8inlHi
Yqlv5YMGmNnyB4OZlUZfnHfeQFEkNI7uS286rZSj2/T7SStGPpk/df2EnYl0C3qh
D7GFhSbehQFspHkISRl3bGG10c42KOV9+WpeGMVhNSZJELEQ9P/q1m4oCTgrYT4L
MyaNrDWu+k+w48+2SgNFzyH6E5UPHLlA2qe4YRIINDJXpr+3lzPLMXdcXOuT8GGB
hRsdG/bdnjDNNRwZ5EqzcOex0uYlk0ejt/z1HKeuPKU2wGC/9NmskOP4TTHqOuhx
6jNMRCpv0028U55Mgj1XdXSZksT7Zzar4S30ChGY7KHafwmAtAXpRsS64iSE09l8
TF69kv4DEMjq9U0mIRHY59IZpmG5Bxy6IYNBtBuhlEGdlfKA4Qb8RKmLwOFjFDLz
d7FCyBth3yiKlTXDqYpX0EyiO6ojjCfLxsLjl40omiPEa+u4wURUwaolCwb4pBeM
JxMjaroBx8GDS5W/COZxzFXn3wUQcd+nEQRIYQbAZRJdFA1dAzA1+IC5Dm4cumye
qPDLbsONDiFTG3s4+GsiFoUJS3Ou3mk7f//eCH7RKG/M1wf9522nce16U3vh4ipo
KRtB94zuVgLuqvpfSEjFGPeQd+0XnnjIUzFhDmaXCWq3bAs50LZDexp8V1Dliv7T
nRJBOVZ4T4QcPcl3XzkcrUjzqZbZxVnojIl0y5HJtPVLuCj2GayRoV1U6gOQENMh
3wxy4hO/of3tLaRY3OeUZ43YvSy8SMZKo8eS/X6USzpDioph2cXAgOQ74BHomb3p
ROAullUTLv9dag8sT4zUJfkO2XPGNsQxsOZSUiiOY7S27IJZRz2PGozEgdXwEy09
bg/FaGXm8wQIrR+ehs/TunAa+Rqhy4vNPKVE875udyl+Poqz/8qleuULtCt9IR8Z
g1XtST6+WqzS5QToJc1pxURkwXBYsPOV4g9FGU5C6v9AKesXrTl8dyjltCCP8fRR
VddSHcSIXB334jCCoUcLmr/7lZtce7zS/OnUtE6V9XZLponE/pQocWEwXnMvK1+G
rQLKHXyl3TbSwN8MNKX8ORydbhF/O1PR+kxzVnGqULeTT2viAo6DTpiSz9C1G8Zl
c236lZdlQGpkRo/2DPRvb58NV3+Qjgds8ZlEhovm4GVEhSu2vuMlJaVetKmWy8f0
9vi2O+ZGVWSER+8v3dcTGzQMnzsDa6kws6KpOENoKlpb7BGARtIAt3fVrhyxrD1T
FKLlY2MvoTk8snqwkhie7rt3vTQcG4JH3tPGX43hsElpOq/ELJjCHDWjvScNX6pj
JdCKFQw05NK0qvj2yrHNJXOOZpnUAyuCMPs/o9mBYfwEn1E9q2yEgWpyTM+KXdn8
AbVURrfZ7I9ua3NSpK+5TqgxgxISqiBB54WgtA7J/Z4smKLF53631nYIeVALO9P9
+dbr2QZCyeSJD6FxquGoPHYV8rapArGvWGDsi3fdQl8AHOzXkxE5pdUx6j2Qik2c
gD70iRTKluvbGhtLBnRE4g6gLjHQTNA4n7GbE+cKnXYmmLoiWVl6quUKcMhMR+1t
rxyj5kmmmxwN2rd3hLW3PJxPEupP7oX+nii6nDDt359LVqpOcKFbvPLWyOnGRvGR
vYnY3qzykozTVjK1KBWHhdjQhETWD+pTX87MVDqHnoaICq08Da/c7a6XaqH4SL8W
156ow2ZN9roOvKCkjJlhDWzjd1Tsl/sP2vaHIzXNhgq59ejeBvNmYR0qBFRDDjLh
HQWGbaXeaT4pCLAE5UdNOEZrj69K6CCbAxgNbaRt5UVpm44GqyR1L72TlNM4sBzn
UHhQbbbQ3jp6ySKGuTOqiDQXH65vYGVkCI7O/UAP7J2uyknlTFKB81Ab2oJ3z00o
LHL/3sXrP+Tp5pmYKWNKaTmS7te5nk+p6RsHKELLLRV36jlAaEm3KCjVuQe7LxKO
nDnoDZukZCHiU9rE+acf/vRn671ydHzQU+GKiBi07QU84+5J/aaVohLVuIrTyr/S
piCO/hzGkOqt/ayscnE16R4PTMi5PqyMlvOBuesvZgBlpx/DrHb3cmv5JDETXs+Q
9UPne/dJy+EOgKBm856WjkSxIiKE8/xOencj7GCD6bZUw3beLv6Gq0PHxKE2UELx
GtGivg3OqRwwj6MVcotGHhsgK80f4TB7ss9Q6CK1G7e/9H/AUB8e8yrpWTDpky2C
+JoatzriQAP0KrJBFzGiygllRyJrnyDhJv6kItTf4Aeq2wkkgQ637IFzrz5n0rfJ
YYwBH0kiizuVIfYv7AAPpKSzDwUL29gFjZA/s4q2fOjM+vNfObSfxsyXnQdqcyq3
15uMRz8gnH4x9DqdNSbh/1mIagle3lMvwSDv7lfn1/9UT+3A8hACf16eGEL7S6iP
EOM6lFjCC71p4JdiVilLtihYPiI0EybN4boz8FUPACotS9+LVExHvYlQV6cahhBJ
oySxIQ2CC9AScCxRggS3zajvSnSk/eXWEHmcPKYA5UIFQvjLri4zG/2dWkhTPp5J
OBE4z8d9YTsP+SN3w9XO0bR4OA/Y36BsgRGglBxlO6xU8do5ZbJXgqqZOvhMmOtn
bLMDvI+g29bbXlQ2BZCb5A0VdU+zbPMu4vOP0YJrTE4qomz6zWr3weMDfLivWCnk
qdwDpDgPYG1JLyY9eK69lYg0/d/62Z0SyGnrV3NSBKzWaE1CP3YbsdRGpXMKzNKr
TFoexOnN9YX45BhyE4Z2WdBJuWJSYoeCUIKJkkMIONUqnBoEO1A0hazRFcQxyTPX
6EMvEFkmXhlNHVfEmAlZx6iCI21FuiUSrWyD6HA/Ey6+UNglN5HBqxFpi40Nu1kH
RPz62DnTS5iT51SEsF2C+cCHJrBOUdYh9+xPM7hNkXu846SGGIFflsawj6A8+Gv2
8e962cZk5XJmeNBfFAh1xEeitMhZYZMAQ1oZnwUwTu3jZTxTcacu3gATtj2SLV7y
Oe92EAdIWC4Glb7hBn7ioRHIHgA3RnzodZZNBaTVh42oviAyA/GgatTxe5rRujV7
dXUqpEurbGFzLLd5jJaYJpQs7Eor/L5sa/B/Kcio7Ord9DjywMqmMt2JjrbsNju8
KSXCuHC55qWiy7U6e/srb5wSP0m3gcgkmxy/uDkGkMpfwcwv3JIbfHdospH+HA/U
ByBVjuvg0EM0XmKfPEH0UE3dv15xiMW6F0QmEoi73WaLzBgaeQZJLSRHg0eUsKuc
032Nf946dq2G32CpYkAiO7wVqX/2ysc/lEpsqmR2M9qhwF6lZIqAzwrNtZ1d7k4b
d5oM5+8hwPOlnJAwDgIy8ffS6YwQHG8MNOUdPcPn+KjiCaUddWZjJpgydSgQpvXt
WiSINvv0LobgJJww7PRx8p4vzMNCwD9HUkXZ8pdSnV4ohMyFXcPaUMScjW9uMb/C
c1rC/65JB9FpXJBHhs8ZU3Eg0it82bSZJ2owRoIMFNmNER1vFms/yoIWXWDfXZxT
45lmt+8DQhWOibFvBcosK2lUrcL98qKK7KRmfI3alqFqRFhUtP3eIwSLpbc93Dv8
4EnagS142613J9J/GTtD4eCw/LHPJIL0sDuSkFjtRvg08pyKLxAzpmVX4a8wYT5F
w0/6raJQhjezLY9xOgxlqdS/mjLp1OvyckFd+Xo8cnaBLyUwVk83RV6BG23d7aSm
NZrTQXNXOf5G61UjWiowDhCtLeKLzdIiQw2c6nUB0K11pP0YPfmCz2oMfNDEp/lw
WNNA6wtbKdDFBOiU0C9rdbMuiq8zMR0fpAnn1WpBHYfbE/fSdLbspX0P64mZKiIh
iYxRBX1pouE5QZzELtEI+82ZuMzWippbjJJUyu480TOZT+OxBVTFUnCkAh2ar1uD
LZsGpa0JCdW6aRvkuogksz6e77AiNkn2QVRUldCN4TsUXVCDPhhHvD5Ec1Ktw4c1
Y4sKPzK18lXUr1u1MVAbcOW49iVXCkoP4y18CQyvLXUx5iFIYBAIuMA3SEjCwOyN
eN53odgrId6Fqa98W+f/vnL0ItXXUHkBLooHvFt3ABuGUjJmXsvvf6fLQsH1aP2M
wtgyQWOCP7C4XVUumQLEOTKp5aJsPiwohsKWQrJinndWL4WaW/A27RYVhiAVw97X
Sg9CMhM+iukw/Iogv7Di/TVrfLslzVYCVV8gBjASThQ7rsrlUXvmAleWrGexPygG
nf+tTZbcOsTTLS0RkUHFeHmhUY7jjuXGNWYdMs5/8R1HtB/t975QebgVtd1FdDta
3c0pK/1GDX6YpSxx4mZXSzPZgbYGVRqy2FLMXezqekhXRDOoWGeEqXwTjo6kdXZg
0QrcJnXmUa/kzGUyY+y+wzhsyUvP9iOQF5yid5k1GQvr6HHyjVsAbYFHPSZYL6lX
QlPcVpPC+eq4OFz+Km2U1npegy5LhIZbHS8F1th//49HzSOLtFNNrruTl8FcGtCI
oP2/lxwQbcfcaP3eVwKDxQDOlelo5ylx2RWQwI6kGYYna0vdXseGoa/TJr685oNX
h6y/Tijjm8ubDsQcB9RJSZdwGEDrR8Y6BKMUpTOoGdh0tpC4CEiLKOCPId59U1la
V1/QP2hnp2Nk+XItm6q8nFtgqtw8+JEbbBcnL3r3+fre9k3lOG3HhNU7HPTW4k08
07lFLAO/FG85RA6+SWUQUzEAf58lUeOzdBpIabr3OcugGkjFsQG3wPyP8yYY5is4
I8IpPayM5qo58CI4rUa7mN5pZpbNyKvSE4WzXsAssUk6vhegMptvK6wu1CP+9FSx
zsEkxfcXQgkmSCcZeDgLG00/XSKhQZMlXMo2nAk0TM5LWoZcERRzojzQGHmRd02z
YJGbYHnIzBPOBmVHybimoVwAVfXbWo/L0hy3PBfuUzbhoOmk5CuQoXkZW0g9jjTm
u4TRXyJph17M393sVur3ntAJdIbfC2tcfWc8AuAvXAWfJgu9222hKbdFLPuMbwvb
XCHqPHuk7uoWZ9ToxvwnDszSbzERDFwVZgRO6Y3rxV4QvBFall5eIivyNK8Goxl3
qv3a1yt98AbfVfGyTIEd+QDeFA8zKCKG80nNk9dlOltyvmh7r4/vUyYrA//27SgZ
Cfq0l0EEkYz2c5SRTfmzwyRswyoYcDHyCW18WjINkFTKe+F9Sw1XTj+eM7JW2dck
GZFyVX7CKjjnGmizPLlb9Q0nWWIbioMT7tox7Yh9NF0N3qE1bRx8mO2jYBkNQ+8z
G+KCTAsS/dTdSyqqYSEJLKKZld7rc1FXO+npSUniKUiaPmdUiJpnTqOBM5/2s2HA
KQH8m8+0NH8zGtgBbD7AmSukLldKG8u7z1cRdqPNYusvRSy1B5V5H97384nx5Wyx
aQxd+5lIYLb5O0tZf7loofMyNMesZlfMGTxIhx8+bqYXGk7Xy0iVWUeiaaucCqc7
BPg9ecyuvOqJ4yp04LU3OVrA6KzL87ty6QibqGJkCNARGjQNB547FUaQlGOLTESj
5hPSk71qwfwKJVu8Q+p6Q3BZ2lGhyWyUoPVSxNnR8xs4RxGm7WP59mvEB2GHa1hT
sN5XGHhZa8G/xBlbNWb21Whw/Z12pU9/HNYVxstcSyPjy2E+HVg/CHlTVWCoWcZV
RhU8vpM9z6lZ6HaCEqe4J+WFandGe2QauRXhuyo2chKhM6qp7h5ulfIwpx3klq4A
FvSrCeaEo6a7f0fd0k4fwXD06laHE1LlcvdzxDGBkUw/L7goVCPLj0krMEw09UZ/
cfSAUPNC4t51evb+Sn97IVw8ia9iWRKSMRF2rqbZQrmsKdsASwR38903Ef6ULt09
I80FiWLPwtq0FYwsR8eURBZRvrH5SzkZlApxeRCkJg0L5r8xDZfgEydsQpQQVI2g
UApxOgGFwWtdsS4OGqvSOF8Lpgtl+WaaA0YHPVwfJWC+99l0c4AhGa+HOnuVJl51
aZ8P6oaKl6lkHIU/zxd+E38z/1aTfZ80YvnwfSXQoz6vOy1owQC8awFVxs6RYxPx
ddmYCU/Nt2/Zz+npkrAjCeI2WQinSjJ2JyswBDr0sPFrQe5jmJwQl4vcfbvS4Qe4
rm82prGNOnOCnIq28qqdePSWkUNTVAirUNF9UAA8yoqbpIowS2KgiYj7jCPPAFoX
/WUPkSUnYUCDUBVUJtp85Yc+qElYGs0efFa02IN6VJDcud2vM0IAQwy2gc3GOB3v
V0fdXhN+/axBaJdtdML4n6gftCfP5gzBvj7HnJssNSadPKL+hcqHvSlO9Vf54IJ3
vCnyTScKlNcHX5VQXhZQSn2XG/xvCFO4gVt0pSuv7ZUihuhGDVET+EhM0geSnEjy
WJ8jbEPevJpork9/9oH0nNeKHKr7fCILnoF2XyffHNGl6z/nwIqQM6nywJQlQC7P
176z3CMSRIWAnwW30lrS9pONaMjGYBTsOqHq0Eld398GBXcK5dwM/K+CgZPMaysY
Ho1/Rudoqye/rAdwmcnMMRow+/8JqI84y+tAbto15gnRVTMftUNucNiShLPhVg2r
Ubzofc35qZ/ECFrp84syoP/qWUrf+nZ4dXaDQC3P+YOiqQ6XAa7CmNy8mqSs18ll
jXCc0IFyibnfwoZy0O3gumbLtDTe9YucuHOtAwoRZmSAnV7iWcF/zxeOeoEAROs4
uhKAk/bl6pbEM8wOQ4I+7l8MdXxjSbnnAoOi5v4ayx5bONrwM5LH94D23By6/Oal
T0orzA5Daqh7MPv/XIdyEJScV3qJ3hM8bthJ0FTZLpAjuJOTiZuMDvcZvU5QKZuz
wYdbzAVpcEgGIT4+a22M253ub+aak3qArBnLjreDNFwRVl1BOKyrjnnGdE6ZOE2E
bAdBCkuRw92trkZZLZ9z+GEE3cMHjwKzllL3LrVqMLeLzg5dzuoSsDd5kbipVOSh
5Rr5mxDDzcyZijOW4Vxh3kfTgB9uSd8IDXY6yl5KLABiAZvQqo5tQsTIgcwNcyfE
xZ9k9jVsWbOia5K/dHaa1e2Hf5AP3mW+gjpsVVVJ8wdJ4eB8ZyYXBTc4UaRiOdiY
UFtaNU167Dd60omMKVftXkCo2/uNlXv6/zEi+1o+FWxoevGeQqKKJy468CmntQfv
6nyywP76pzIN/R0EG8ec8MBACDYlOaQd7JEznZ4JxYYebt65uoMIaLddWx7VqNiy
vARyMwPY/HfcqgvUVCdCniwttKizwnHjxDIHNB/apudtA+k00ipPWdq40Uv+AVSy
0y70Fu8dZ/qC8pSP93Xl4v9AgCFkeibGum9UsoXW86S5ocXClz87Ukdo2uT+nyRp
jx9ErHszSxXyC85eKrV9ub5Oe98TbB8gEEMENvn4ZS3cRhtDZ73sDR7n+mhDe8X4
A0OAcy6/QkkyOCyXbexxy3ra0R6DREliyjsPFaHPfqt9xzrnknNeQfj5YQ5R1fmk
gN5stPtJ2tytcFDCjqy851yM27WsKjLxE7YTomVs7yJXWf/+l9PtyLQ53zGfsbk8
h/f5wzFp6eWJrT3B4HNWfO+q2KOyzDrpY2QxNHL3HTN+kvcxnz5kqkj9vEZtXT9G
cAtYqowGvAtY6Z8V5P0LmFgKhFDa6UWl5sL6SNf2OkOEfyIeR5kYXzBHnXHtq30I
hCVQLqGJ/sdQbG65NRCcp2jV30aWZG7uxr6Gv2H2B5xrEJwz3UmiLiLHa1xnh/gd
WYZUktYJzbL6B68HvLkkJ2PfWGo0xF/V6BiBPIi3MKElpU2NPk0GqPYokyIDI4gN
ATEHcIaVj5QVXwNmGFsTzwbPPq1bqtIf+K9VxiLjkdEX3tg1OF5Q6tDziFtHEVGP
g3EDhviOI1qww4A8TvTyn80BUdL/l8ZT5dPte/MeVhmVSTObLFq8659QPljdy6I0
KSz4OV9xmz+YfzNeeZ5TdwtgH8BEs6/ZYNJ2imvG6v+31UXptlZhhwKPv1V/Wlu5
Pe8bCu3Y7r+GMVYZ43GjTUR8YQbJHG5vF5uBhrxXz0CZaO4nX0wntTh5oY+FazYH
QGut6PV/wLPXP1wysaPDtShkqJmVmbwcFT0oKmyNQyxO54isMf6EeFGYl9PX0tNF
bcL045f/tMQnrs1jjCpqKe/EsKko7W3Y/Q7IzDCqfWM5HmdkQmUf4cIbcYKnfNSv
TcfG7Et0K+wXppNCbTGfYfSDiXB/sEsfZTzlBwLvEs0meENn7ndX9rynqt2lVtAq
YH2pdodN3wXnN+oJ8Vk6JTdFsJQ/4Omr9LwN6cG8+AFpS9B7OPravwAaOdPfGiUr
dNjuMTt3HFIGy4fSiRXu3Y2raqa7qYkiXi6pPon0ugRw7ND+OlR10+lc8zZuFkyS
/IaRMDCOe7INVTK1WXSo+7uYxFMbrDKpoU3YVhF7NU5id/8DV5KjV2Xef/1DuoD7
lAeMPDt8UlIh4L5El9ZObghJXb4c2N8iBkRW0cL4ct0UBLObt8ry7Az/nFFGrLS0
/frZvH5iNf3FK1pWoSKl64qZWIF2+x1K/Qca/NbFgB33x5/lLegeXmO8ois7HV2f
Eu26qgRsEPSQqxLWb3w/4s529GDBe5KQrZuZk4Xb5/pS6OeU22z4aCLR+2DSiouB
jODTvNYFD1bd5qyBhYLSUtDkG3kgRor3KUxEnDAIbsndqe9p0kVht1NiNV5i+Tkv
ye/PxmuiCOjgWCjA5R8Wg7TwrEl90Qx4xRLiLOOvXGVzjkq4u8aK7RfUKE8Oo2bX
ZViGL5KO11l1sSazgMhn14+wAiv7krP43+LTMAkrcSJkFByOPvGg4QyhY2CmIOsO
CJ1B/sWzEC5n3e/RanG7RDLJaroeK0gR51+ECpRvohFPnXJ7Zr8NvfZuZ2R3G46u
XPkReXC29FiQ53X8HywsB2DyXQOCj2ELLVla4Tan2wwRlsZuZCbjmJTFwNA/3nJU
Wo6rAeY+dcklra4eWK5n4bifBLXCDjGUJnCIJUzXuxsPaiQmFSTlKRzcY4HrghH8
g20H6FB0bRyJijkoTh2Pg5HUeF/gKvj9bQizF1hT7F2yy8h8bb0IZtnguaIjVLP0
R00vsxiKSOF/LxA1Y9/OoAD70IXQ4s233aoReCIuI8YVtjt0ekHy98VueLGDc4ng
/VsEgWIAl8grRwDEV3xjEqYcDaJ0gM8OZZ3x6oSfIpr3dlaaqd6QG0d5WtJr5HNw
+G9vCmfTrp+S+TkhnlbANxkY/Le27nT7K0MYzqNJB6LwhaYXPtshgockctnNZPws
X35OKKdyOsBZUyx8WaHE/y3BRTcpZXYpdSJPwg9hOnL4Z/sm+ZJw3s1fHPeDqUFp
jjZRjswYb9/rGtuEOKirPaIsH++QyMIDgY9GMR+uQdnF+MinXY13nJcHJBDsqx+w
8m6ixoI1tseCZzi88o8y8K51ioZoODFrXgH9UYrF3OhkpJ4ejgB6eESui0ZFbDWm
vWgaLD/3fKmhsr7PUY2n7xuZA7GbNMqVWgHdhgxxa7j/I4p6WRZNoD2Tab9uS39W
fQJMobJU59fft+Sax06ueUv4YQqWnlL9E85XiOYEzWSIRMl4iMXjFUqnGfIVbyFY
gwzIJJ4Y8B97E4ToH8Qjb+dIleW6lC0l1m2Q3ywjjSXMLZFIVrdNajp5uYjag/WW
NkS07xfCCeqxOyy8bWLNfXYhMSVen5wi2TO5VzEx1Oc55opTuypoH5FaQIU8DOo1
rS9MMVyBipeFfCWDY2WqwPuKxybtXW6tvRZZeVWpf03kOa5/7I7KZMMET50x090D
cB6wqj4FbHEgWBjywlvsIxb4y4I23bDA1TI7Jp6s9d1nqiSojkPHoyoT6XucT5Wj
0p9MHqfb7npg76BwWHBap1xvOYUTNQzRbaInVY8Fp4oyeGNqWpAkM1lrqUG0N6/K
iO7zbZXEO7tAvS19W9MtB3AkoLkmcMoTWmbFKSsGUSt3LobicfsciV7YnfNlKTY/
oDP6Sn86LV1kglJ4FwrckFl3B6Ic2RTzQuphRum1qGAbPYPJGwChqPbRYiBTz49j
TYkTP5n+OjGZgbqx5Lsx8fT1J0y42VZf+bKUBOJ6diTUfkuA/O692vJVSrRv0Q+h
84KTb5jBztNqtg9tV+Emya43GCqssHehiOS5hvskdIXehQYuVGOBstovuwzZV8Ao
m3z/zMy+eYOlKs/axtVPUoAVNdIyLP0lkaOF4mbWOLAtn7Np2+HOZEf6qJc+e09k
VCW9upYfHqRn7679ZhTfbOsfcmFz7XO+763L/EqbqXuSN7bKT2uFrPGeDYN0v3mt
YJFG2T/mwvc9S6KHlpYHDwK5ZhpEgsY229+9oDo6BnLo1TTL1JojL/5OwJZxAKii
wsFxbE1Oy4HDydBrzcYCFQDXuNt+OLaD5L7M7C349lyf0nNqSEy5zy0BIwSrO6Az
emHkfOH9rWoaIwNn/wDek+XT+BIp2RJZtXJVVcev9Gcsb1rVr/OQoVktiJSK2pgR
XjYOUp2oRg8/sWdCkEA+QICjo4V+/QqSSE3Z7yiB1O8/ZkTPqHtfdtendjQVAIBe
2lwsorx7XmbIwiYwDffxGDQLxSJqEhv1aB6gKYSXEdwAHhbGTAd6zbTqO3pnZ8/Q
0bXSVyDmQtKZz1XnWvbek1iKZMCCJYlI4i5zx53T3bbaGFNoiCYBOIJRbYId5mDz
VvcRXLzEtXLRTK1wYAZ5xk0xJkoOcr13lGR+JOK/WGzuNLW2+5930lbps0OIw6Th
xXXFBz8O0w2uh84TXRzuEKvTFbETAFPilOeBfAQrllnJpjp/92mSqrPnct6l5+q0
x+vpVgpe9N8IDtWfZRrBauna+ybiW0yMMN36JPc8Bil/6ycBIcVUM1EI/kCQdx06
FYyPef+8uW92DbDQJO+8IYgHtzQkvfituxQABFBguhJC0gWS+A7ROTIb0Cn92Z+A
piSM6VaUMKhcZKOoDCchZtx9+L69iHrDMlS+hcA8HHwijLD2cWhgFBjDK82qy3SX
+5CD1DP2OB5ifVXfhxNe7oRlsamTC47HpNwKMPz20s0biwgFtHIBI/05EaFvX37C
pNmhlYzRJBkolQqDYVzYHFSXlhOgx2Hso1OgJLOuBIpRrWalnF1ubox8Xcc9Xf7M
Yg8NCG9gQIqHpKaILMlPbSGSQL6BivnmX3h9nEzJItoYZC/gXPGt84Hvc7uvamqs
qLboTFGjMSUHlhkAEtgQEApOcg8JVk/pZ/EhyYlzOLeAuA6jUCOzwwaNwO37xtQJ
JsHjLAZ9LZ0Y3ChGCiTPnNWO9ghemtxcmHAvCM5gfkKe5vOg++UvdrnF07F1eaIo
tyJL0ecOzTqBfqY301MGxGgFVJqJxcYSTBfECpXPOxMVHjzl1mEJOs+SkKZUVINI
txTEaycxkzbILs5Y7PeN/HmNJPbyOwww2pUai9WeHhGnPRaXd0hbaeDbxq9Y3uh6
Glic1Zx26PIj6n5VOvqBufwClH8xaeThy+cyXh4JjLcKafd/Y/4NzkmN30mby3lR
f5I+VEvLUsReDvPUupxLjbgnuJOOayg4hIaSVAGykRFpG+/HzsF77zttMWD32yEY
TB5g2ESS0qajUm6mTsH4HuNP7FGeTdQwFHcVmBQs8kV6uq8+B6xdcxFTjE0sXEOl
psY1kZb/ImhAwKr6OBIZKXeNrQEIjOgAAkIGqx57PdRGb0Fkhtlhgcl8vj0y1Ny3
A8c6+ODVtAo2hT/fydxgXkohB8cZQAYL7Pcb00IllPCpYUndv/sWMtNgGN1CWvCs
GY6ra3WAhazNg31TZpTcIeSmo7As2FHIqH84Pchk0+Z8AWxyImidmzPPceapuhCE
q91cw8PISywWpXZxDaO1OuMICtXJHBXkwvJGUZvYxasAMaOUy1s+xJHkdEOhjBjK
lHbIFES0wX1tcsA41+RubjWc7c2n91uz2NpjOp0hU/IA+LQalajKnJ0pOBSeEXt+
Son9a07TyzjzU8anadqdo87H6Q2Sg/utqBJNgDYtuqnsy9OgSKZD40QKDBD0EwZm
te8peW5V9S9nAWr7mk6N2//zCET85eatuFP7h0F0MHgQLmtis8nRk7WS29LWOKZS
/rSdoxHe533pjPxeQQlpM1N/PamJ8oX2i6Bz13DOLc/tlDFmyhSjdie3cVG563If
CYnEk1YjApRJ79N94XeR+qdaBzFIIwlQD2YPQw2oS2hqFHxBoP3cv3SJvDL0JfDc
gjJq1+VlJEPeC7eeiv7ItV7HdZMp2Oi3PMlBwSCK83BGo4re5cyb+Xo7e3jEuN5U
Mn4ZjSLgqI57w2MMpuH5UKCkVxnEmWXDagBuMQpVS2pqOML8d90oXa1kXw9tRP1A
vJgEHPxWWmYsVNw5smlpkkEIwiYceqft04/2LEniGdcUvtzL3IKOzLwdY593S51j
lVDpHyptOEbwWhTx7Zzrc3RflVLg2zC7EAA9X+OBD+1215ZJoh7bQhY3sF8rNvmE
qdnQ0beP0O7wok+iz1xqyn2Ex5CdXpkdzGS34W2A3hLdlQnbE1cnzum1TLtO9MK5
BOKhH0R1Ds2VGU42StiKFARSXrauNG4XUoCKLkYXCE/0YH4jF6z3TFqMwZWRhw6x
2zCKqQtxPK8rBu+FUtnwrcmSJ8kwnM++1SuhgQkviwxHyIxSQ87LzE02jtiTEFgm
gQ+XFNxkG215gCO+QILYS/Add0DpaS0AMSg++eaC0adZiL/YxzqBBrbbRzedBkOa
7aK4+e4YDekJ5Elf+Y2Blsl7LnC1CWXXxGhgRign5x4pW5g2IMLVtW7k2Yq4k4MI
HDY/mqIEioy7MQWCWxjRwiYelDWIGbuj6txPzd9pyM7WOyPZz1RkUdCs7Hu2VNcK
hzfOFEOhLmNNYUdBzFHbDsSxmAn9iygum3EWSzKB0JjcvHiiReC1ut9H7DPYw529
GEDbRDwfRfIrKtwjgKsB9ZDd3UJLdz/3a/FRaCLfM02KYp4wcGyefI+Ze5YbavTO
+jXC05Dkrou4iSRjuaLR6ykV+Nz77GQd+47XQJJAxHJr4cy4m3TiDOgP4jtT7xbC
wZ/QKm6h1+/Cujgae21qlH3kFhV1OTIQM+JtNhUJEo2nPrFUl2EkAxvdVgzFhU0t
pqh/slcdwyx74d35WLynTaAQt+aDAC91adqjhvSgP7GF3F3t+Lo9VkTWXYHUSlSM
xSR8jaIXJzfxfz7CgW3xECaWgRQibgaN2cN5/niS+xax3kWO39pXWonwbUV35v59
zh/fvl+wWFxsmdXmiYO7ZojD0jlw4ApRX7zw8xW+gFpemSGzZhlUVtox0YjJAl7G
/8j7Bm58vmVNwdTv/hIHlGIXobuqNEGpvYgE8mPBdOlZeAFL6MyaW5GB2pNj+Ak6
GbMoWwSRIqOp0Wop2WfdgC2cUsTo9jHqzTCNC6Qi//BjyifpCiWLzVGwmgpXyL7b
vTPXcO+i6yVSkFZ+WwQ5aKbI83ob9kErkgk26W/iQhExhcMoIkfR63hX71RJ+gq1
KoGqNvkA7y3d0bAgC03NanMZKh1M9+KXhJnErg4L+7CxKQ2cP2brrS3X7vagqQLD
Qsv+oHH/4JCyrvLPFoYMWV90X2y6No27ICOOVwIY8gYQCxv/cTtyfn4QL3Ug/40+
0+Qxb0LDeX+eGrIPyT6BZ2cY06RkgLhSqksc3SU4OmrVYKq/metpSsFDFLaLDsdS
YcEcCT8N/2Y7ajwc+4N9EoboqeNlPrwMLvxZBHYkfVlp4xjI0zZjCC/f1FpyPn/z
T/fCwE814628Xh1zyBun+jx6Gva+pvMVUHR1VLi4Cia4WhjRtECmWteaoRUjfkbM
IvfUP7vLuVEgnBhclCX9CjSjLS9qVr6bhWuAtSadkz66GnGn6KSVwfJf5sjIpRFs
PQKGPQqrIfc2cSJGVLupjc8/92aoULlcAo0N8U8gQGd3YvCbabi9C/idGqR7pfqz
haA63kquyhjpY33W5sJ17+lOUWcD4Li7JSr0p2djWGwZkd+eqdxhlB1RMjkInSJl
z4kpaAFTlZFnLJzaZ2wA9thSl3NCZzZ/ucn5fsMxQnefElgsDn3JOWbhP/hBoUrr
5Ru9SBDBch9UjDkxpxYAPS/M1E8tH+MGZrRytynn6cz4TfjZN+Ugk2cH2CJ5aoy4
Vy9gzHd1RbYEVplzGM+i6NEbx4R3QvSi3HoCUYiXTNplGU7whHKj8AuGZvtg/h00
x4GypkUWHUR6QVJKqfwZfc4OPGFu5xaxVaJaffcaWSbkadp+04NwOT/ncJm8drA3
uAd4flmIfULiY0REe9zj8tVf3kAtwgADHafjW52he6NKVTmfILZmKzenti5MwGfF
tTcgSNhMvHq0O7119023pGJQP4wUaE/XfWXf97WU+jr+JEMuUJN2WZpgtzDOD624
nJWahxMTFHKxr3IC1Ga0mE2gmpxpURL+CwaLr0Wzqm7l4NvkmvvggItg9nPhCs2s
fhEoDKcMijfm6/0GZ2N35tUxdoiy9dP/23B1BByvhwzK6y2uXmvn6oGYOFOGMyt2
Ft0LI+3LVkTp52DY/oi4NA8PGmm/Q4R58SqbZZN8BE4gIZBEegxwZPWfcHs04nnK
pnDGxI5wXW3NYHW+8CIis7j+6SxKc1T31QJtBfagjLkq4yEu/jbFxGIEFt23iYCS
G6O23fK6/st2rPjTVop7t2Ff78iNOUzHZSg216L5Fj1z311JfG7f3JPhap5NKEfj
hd3dvCpyuvD8LRbA7gl5AD8YimlfulBtt4Fo4LF+O4fBcoCb4L0qP5EqX49MTSqo
CYuS7ODFFvAJEZZRDZ6l7vXsA9CzgmQdE5dteppa5jyU+xHo/AJAGv66px6USuOG
edoPsEofmIQzPq2NUFQj59/TApPid0ELkCuJVqrkh9Wyy2v236ogkCmh1lgBqvNK
fl0EwA8zYFlwVgpJhFoCAaZkrS812CAs7BqVoJaRw2biwZwXPMgdzdy+8Hfs8tp7
XnXaY+6D9cPSK70SMcy3FEA2N32QxmaQJkIxemciQEem5MS44Lv480FNbAojbWcp
PUEGR127rKpJwpC5Gk2wbGDbcBKBhnjoxsSOB3LeibZcs+WVrEMdiSrZTHTSLZc/
DY/uIt5asySJbxWRNPoK3OV77Js4ILt9YmcqM2ED5OTJZ8TO73cIRVeRU1x8Op42
DEShAh4mvdIu+bUL533bt9yQ9k3cD7/rJGXSg5oBLGj/IpFY0tZTWOROaDItUT7v
OEcbgE9/2hlBG40qw46O0+ZNguEqkLNLNmy5KXfjE1A2CKVVTIXPGCacqbPGDH5n
MagnNi74XwDAT8B3EYGCy6dEhdCFJrgX5ImlF9dPyfU8HSLRMca+QNW7PKRlQOFR
ePFLO8P9FI79DOadxEa7ANIIgBGT8n0zJTZ9c9c10sVKjE3QROahKaxVzJOpeOQu
EEm5zp5QWFTgeS+zcHbmhmUEev2mSeBmuroc8JqVU2UTQwKG159JBN40RLhzYMKw
4i6IXEWFYg+D8IQ4u9fpz84Chz9RYVXJ+AwSOQHa8A2CWe6GmwKkRSJbPrB/p+DP
4TWaBjD6wST4vSq0gbYcdrq4EuX9EX6t6rwSyBdXWcaMo5OKkEvrMtoZZhOtV5k1
kWnJ3Js1iElkQz3I/GrtT3j98E4p9huGaHmIpE6lM2TXDihKb9brnBBpaS9remZO
h3b42TRQtXBavNYeLBLbROT1Xapn/zF0SA1yeo1PHjpU3tGG9Yh2olNY/4vnIGV5
0JSV0cJ7tIkPqAv+R4ylFVZTLETd8SGPNCnGuYZorYtB919GM5QS6qzFw4XHgjBj
ZVUPkrzkDo9749oUAs+qBx1tI0T3CwS26gtaSk18P6DSSQM6Byjeivh7ZHnDkR0v
sVHk3QQSc/Pdj7v7ajDbXRyA+rRbBznc5IQ2r3QFGTbOldlVHys2hWMhjoLeaEJn
avp1fbu8qlwr7TEydc8dGun4yx2g/IlkiukTwVzfXJQ8wusdwHp6Us9SUmwTtlqs
NyPKbTxWe+jbBVIqlntWO073pXSG00zVrroWBlKnfYbZQdj9/mOwYeJKFOtgjkCn
tLeZ012OrtENvTh2fhC2ge9p7IT3Q/brZfWYCQaLIbUPvS9BeDr0NKkmrsd2aciq
KMYSnaaQW3LygfrQ/kkDemKSQ2M5CdsnR/XfsMZ0Q2xpI7L6B9KkZphWCiVcdnnv
1R+d1DdzSNi6o22jOwEeGa0W8WANZyytJGgmPPeRg7ylv/lJHk9IxoQNR6D/VUoc
lEaFoVi0g3WhIaS84YZasx7XsOEepz6NH/NbrFBLNEnanVcYySgxJcVpMNA0qwNB
Jt996WnV6HbbDwEj3L/b7T1+SOSm2Z0mNbgoNUaLmUBHfLqUiOMNtZyYWcy2LLE+
crvrja5kfIh3dvLvwlbkjQDzqFaixLha/Y/JNlQZfcwIjBSvWzulugP6dvTRWz1V
HCig1ue9/1Xp40kMkffmwasdENxdWrnnMipzuYaGqEQIRB3msZRFNJI5evBOvN5L
Jh6Y6/aCWKYQ05SihsZrQGwICU0gq17UW9MMFCT50YRyXCKJu/bHHaSP8cDEitRJ
/Kc2bkbafaetRiI3spAMLoJpuhdjvuSkcuonl/UV+3ptVPr4lmIIOoebEy69hf+y
IYGoYhTjnSiSr9/OpkW84vyztIe5yoo0OO4Cgq52aWM1alB9TXqObu7mhqAB0M6o
h9feu5espMZSd+GAXznFMDiMq0CC7WkAS9V8ABqBvQlmXO+nV+wOlM0SNHBH6J33
25V3oJJo/qQnhSJsw/vlKwAU4PNne19oSSCSyE1A+iIiWatQStxZenY0OEcDalBE
Th7TbnZ8JG9aJyTgxNEBd/y0bowOeypOkezE5Yw4N1fpLN9fEmRmXh2l/q3r/F9G
pzCi5Rj9dTmlEqf36lMYII7wDbV9w5CmT3Xn1Ii/v66mqw9GyGjOO/FTPPhCk8bD
Z7ZU4N867XaubIqZ9STqHfqYkOj/2NbviTb1H+L8NZUQNaBJssyCmH7YFteN8ugw
D4DKdCb0omCdnNEB6YKBGzaYyetq19Qb3XmQDB7Q4E4AeMIz0VIk9uPfvcqSH6y2
rErsqOo1ddWivJ6jT70VgQ6V5tHe+5yuihNCGuITjku77Ti2FAx9wGZCPhGPYDnc
X4X6YG1nfolGxHLze0/SQWLz65SVlEsUJWOyvjWeXg+LA/4xEIR6LNHeaDEENwZ2
qhj8aroGVEAVzFlDZh2yfLTW0I3WTF3fTjxGJx+OeSD7FlqRqKTeyid/McHyOUhB
f+0HQM5QQXCurxdsaX/7UjgW0IyOoHS2UAwISaTgzNMtkjJGRD9Lq29EKeydVb98
D55an2fALbxVMmxRwbLEZRit9gogdr5nTO5rvZ0FhCXIbmt6t/WQVVTZiqiP5rYi
Z3jNMD9jHutW/M0OqojQsyTUxiDZiJ6wFtGfRA0IAR+rSEQuzfKL76OO1AS0SB29
qRonPBmfnCXiRs/PCVQviv/6JswHQceSxAaDm4yErnRB5ituD0xiV93pmAauaQmW
YUXrUYWvwM+SMzrmG9A7sZ+17ail3tQmE+hstIixV5GLHPHMH8gFVkqoLQ87c3sk
ZxlHyG42c6xVQbpI4S2WVyDUDpYFm+0LiOPmex9OEASVEoPA+s2wRziM/EaVZrLv
kWvTVh1J/TPTPn8E5aR5Yo1tyKWl5VWHtKmnwR6onLnRFTxoDScJy/iWnH7pWstg
FSopZxTpG8O4Y3cL7ZOexwxAM73MFeiNKVmPFceaeNEO50d1iYK9miGpHw8mPWnF
Z+0bBTgLW2/7sKO55HfZS0I1EJrCNy4AROMm+0qkSUBgGhZU4hxXFgJKGiTTe+HR
v5bSN+uwVsDyFBvtea0xybVslPgZqRRv4/09672JFwVL2S0xk9QMU+R4HIVAlu3U
r0B2V8BEcfXgpnisRnrohmv3m+G+Jq4CV+m1AWmuMPba4QSEBN4anKp8P5Ol++mm
MzFbxpmIqce3C9qCl+H82N/KbxyFnkKcrZNgYXTceobMlJ9MtN535tNzbSLN+2Pz
YmrW8Z9gM2uGE7rRYmT1YCg7Y7BqXp9a7EPhgp2G6OMSmQwjzv9ji8aiwJxhhyMv
/hc6pfxqgJowteHhGHEIswD+q47dqXKpf0kybdKGaQPL6bMBBp6QRYmC2zysB7bB
3xEkdAePwh6VyNhEM9beuvZK/d+45Qk7NqFZkq14vDAMc4h+qnzRtcEhioA2jlCs
hD+0pFeMMjoe9gDGtAXeDsdBapkhZ0N06m1p6Iax0vqg5cgufhnEKireo9FpGheI
7jPjBgyt0tofQ4R9CRJx0u2X+Bm39jtki+z2Xuxmap+8IiRCrDj7EeRzuXMME2+0
OpxRQU7Tid7X/3CpyE6S1BYtBQu3zuxhkEm5GBmDJpF6Djg5HCllzdU/2kbVxDUw
RnEWm2SmBfPmZNTZ18gY9+2u0Xl7ErziiESNpo5XWZoP7euCxOjcNcNf4ToUSl/3
g6ExHvCcqDy1YIvHZssDUa2Y8jAIFZD7dLB5V1vM2szAVUyxY2KA02drccvW8Aeb
98Fm5tDMdTOq3vzmd6joAFQxZBcVUIRYKl+iNWx9VhVMIvjkTFqSZqMmHUQ82yBy
QuI6fT4C0idDcm8A0CFozAI+xLEgcTU9qCcy8m+LpGPHOpVzTedqNx6za+binGIO
6j53CrTHQMqolAZHBZsQE5X9+YfqEmWGhgRZR1IVhL0CbgLr1d/XuPGH6PNLXr07
txXRHD1a8MBwt/02lXvhKUuixm3FLtbOAHWzpX9oTCYTCY31bWOXIb0u0E6Ysbvz
DmFGdIbeOD6H8UbLrPeGULuUUTEKxwM7us8KVxL4uvkOkkpLvTZUFGvyA3fM0naO
iT5TanYEamL/NkcULWMuiIN2vhpflaCdyY7GaXsKb1eqK56VYi0BQTgUcMvAq2wU
ZioZNsGzhjda+xkXtJRXgRoeAiH+E2nNeIVPgq4JRqoaYL01IG+mq1w1R3d1e7ha
93L6Jk0iWCc5e+2BwIpt0n0xxX40fzV2eKImmq21abZIqmLnosrXWVJXiMSqeryP
C53l434fyuKFxF8psky8+AxegS2f0Kf7EtXV2sSKOKruN1tJ1Cv5JmgA6PL7X5cK
4koZ8UeayHUjfjfhl0Za9IjhuxRH5KSujJpjYuNK0jVsszMF2m6cQoka7pE4Ny0M
nvBfLbbPYxDwkBHhvPrKUZbOyVpal6z/SciP02n8x4h4EUR7DjpyecAYURpcEU6E
jy4nM1JOrhPAgBApo4I5GSoS9UPuptG4yuJbfcFtwB/bhxvoPixF5oXo3d9cFO3l
2BMNGKfQptGvRtgDQdRxiKLa+utmfegqpQQIcLgZdt891ZjqGTCfmIg6PEUlHdhx
vO69FRu10jRi9FAx8CKemV+1HDDr13jcNKHo2InNH66hri0ItcmXdsC3Qo5a/+JG
sqb2tnd0BFEJxQX6W067SIiHlQqifHE8Ell1QJXSwRc0hhG7c2hiZlb3erefciIP
Fgqi7TavEEkJtXbwJuBBLKZdqgdR2GVRZwPGsMZRftv8dPLa6IamR+3D/lMxw4zz
SIfL61vIiFQppNgUVqth0xpwurIHHZ8j3rgTGJWytjww3mshXSYhlMwCIpZqITxY
qhdoiD+QSVS7h8/x9sU0/6Ka1T1ISEzJNhqyfQfq+gSFKObjdWsnWuq9sipCZ1C8
PqE3vCwRyodomre/Oo99pz7ueap13tDTAEz/3ArVJW3zB/e0MyURTuDW/Ggbe+NT
z23Ag8DOvb9zhGUjMT9Xejd8no1y2Fsf4EyZLVDcicAlOKLUWpXzr5CBeZxOxBhH
IjRLr9arRXAvO07CbgS4Gq1IZ7Q+InLrNsO5+P6ymWFiKpxviIJqUEK2MsBkM7I9
x/qwoDlI9mChDyqx1YbAlXa59dAcLtPwBfP0BSDZ8uVuH2HfacyR9iYew0Xhcpd2
NGWNWfiCg9yBr/KR6YxjOJn59SnWL8vame6twEGJVelRDjKo9Ia7MHvc/90AGLDN
fIz4z0vaMwAkSnAokKeNEuOYFUfXk9Mw2x3TYj0B3+LmcK5cATOBzWiFnJ8HteHN
KxIY6NVUefle9uFfu01dD+V4+kK4m/qJk6cIOGnwdDGDfyN13SROOHZd9Ztq72bW
hf6U9Suq31JMwYlYSBq56sXn6hYz+t2SFEbq6ATP2sPJC3U8duPXHDKlqM67EY6K
MHbvD/4aApILgJP26fzj6fxT/8vj5GGQxoVUpSyBrL6i+8QpP6ZoyHcv9vSw/xXR
7KSTBcYhKb2BjgVhDTfXmkhlbulSLF3izjjHlVBH359uv1Jhdtb2ZW95cbwIX/pq
F0dvWX81p9kp9yPdsPaPUQtMtsPehgSU+x+OcGwMPla98lhOEzDHUMb3iE9vp1E1
aPNky88MJxGMo38Eu9BKeahrrsGUoacUX+5wEQa4qsFZH4kbIZreeokABpw0zGhF
IonxraiZOWjg8YdlMPs87ZRGc9IRwkBAvy685Sb0+HJWtuTC2QeOyQndxcs0u9WV
wMCroxW1c076dzsknX3ScTIuVDfZAQhH6POdRjjS1JZt5RL026aN0ekCc8jR/w5t
AgVVCL0DxJM4C3tBgV9VQgkzkI0dSOcpdy+Rqm9gsTYKh/o5Qlq6ctXkBcgOQ/Sk
19R2TpkckKOwEx4uXlOEuoSluV8bMFbA6/0hIa8T1U76O2EHFQYggFHzTRopDIi5
X4F9JmbzSLMZ0a9gfCHMmcBTEmCBwL/n4ECddogx970y9BPjelFZ9uNlNQcrnBZU
ziJVwkS/eDnSc/GaUUWFHsu/lPfuGGweyajGa7u5sTxcPEO7m2Uf6T2SqJMf+SWa
lAP5NN3qsiEyHsglhuDx1t3gZ174BIUWwwUiAF41H0BLlWe5J2tHUU4KDOY3gCg+
D0g2kXPWCHmvTQ4KCZOQOY17txb+hDbY0cWqeA5F2EKDbjhxZtoMnc0KsV5llvEr
lQQLiN51NS4ZBNhIQgNZeJvJ2qJRHQi1Tlb4GNoKvewPPPz0Yppc8uJ7TesalKs8
g0Gzt2vsyDEthFJpKLPmwgG8jlUYhKoRHaDKY3LymvjokvdFbD2EL3oyewURCY1Z
i+CfsxdwlCirj6RIbPBKeiPKj7tChjxFaZoOiURpi70wmYOBGPYsS5jDaYzN4d4Y
eBky+qNfZyEG2Hj+BxGB+8UxHFXFuKe6A5ZH7blnu1NWhwExHJyp9B2mbbFuIggR
Jb1TNwxFLfoUqy8hxekHtOjur9cESP2WBPAtcCcbBUYFMLxL/RW0T7FA0jP9yGMB
YAg70rzQuZRXchU9z9YqyAQAan/PZRf/FodqzJqrxXqOuM5OqCwR/l2pm7WHDH5s
oSreGQ51kRnlsgYjhn8f9l4c6+u3DTj7Q2krxmKgopEo8QKoygaKjaeW+85Llbqm
O8nzHf0p5Jv98QvZp621459oBjgqerEI7T6JYLsQN4QWutPXzgfi3w3j2WNCI2Sx
dFdI6MHYJV3xfKF5Vw3Kdv2WWdgVzt1d391qrA9iaq7NJBMEHaHL6POxYd/cXzRE
+EBHL3V8OcuiRwxmgHmGT+bWS7jrFBf7RnHbaaueut6cps7o+AsvEwwf1kRg6Ttg
vh7yS1HKOx5ANYOduWCgEKL8S/3Pi0o/nrvMTvDINBvh6HvHmLXtzmIIH+0UUwqg
NCIfGA5D/mv+/TwwEm/SFDGPT7ZdLBfqdRfN6zb/VLGb8/v6gqpj4T2oGUn2oLbL
iGhbEyYpwxkzJ5FpJN8T1sMFW/Z3aOr9NcCm1Obv/RT2+xJu+Io/jcNy2pzTydbt
t+SuonVH77s8prBa/1PvPBlvA0SIBrnbdqREzMYosrQSVS/1LV2pvjBGClP5nOpu
J5Q8iPyok/pd3wqvcHNZcqPreRtPcvF5nsDcBWEH3PW/ORv2eygeFICfVdHHcmSf
h0tz+RKTFalAOF1fE6j9EWYbLWMzXMZrGfQXpl9b95BOnE3KrzJRIoTooYwvupgs
GtaGsJIHrmZKIqIF4Fa5LJyz0KPJ6K49Z4FXP90iUUnn7p5fcIZp2HoxRe+45R36
cKGqBtMBanKVbhkzhFSwwHpr8/SqTdgUgl8xCi9V/bQ65UhhuCQ9IpxIII7NH1ie
ECHBe/wh8o4xPYBExl9qZLAUUDHqMYR2VqIL/YL4iXMQwFrFduF4aQVdK9qIY3dU
+uEyfRRTQMySbL1U+xl/BBdqob0c9bhX+6sbuxMP8tBVvUlONxxIT2QyrTCFxVaR
H9Hrpe7WCZz8qidGLq2LTJG/ra/s8KX7h7HtUfjK/fuRGaB4kPsfqkFyWyBkcSD6
pvfmdVN25ABrGINVaNqxXFf0ris/Tfz9V2vJcVoE2MDjbg7z4kgrK8N0fKz7vmKD
zpS+PDMpdeFBXtuGog+DjZAy4qOCVaPQeBwbqS6uDaXsDVDJmnFSjS/0lfdnvKzs
QG36N/whDVzouR2FKxnTaSl72SJiqQukJAKqFh4Qt7ufnxIvmKdxv0+nZA8TxzBU
rgeYcwYhBt6a1/1oqB0iatB6MslRMbI0AJoe3ME+xvl7ax+hSFSN+MDwoyrJ3MkC
vsj/hmfVTs9bQrVace6571wfqVtNxqfYYY4rLlRwlehG3dG+HBjPLhGrZvTfumGC
fQA0iGPgaZInqEDQMm3Me28JT7SUuVXXpYVfdMX3LzPBaVLL/92bAWNAdfp6MB3i
vhdthd/xPU9mrnyanrjHQ92+k0SCf9y8+nJ1v+9M3YfJfnIeiWXtaAhflp4sKHfE
W5kpY0kTt0YEeGktZUGLjiwCnUqBvfL1jVJORIype/3UPLod10UyCxOAs71H6uFE
p3Nudil9vHaMMdcDamIsnMu9gwnjWrkuRXGPZDy/7o0T69FYtXjsPISqPOs+ROZ4
taBW7SQmXcZzOMlqqKwsZsyiEWGSbePu79sx05B6FFpvZRHV/Z5SLufoenrHOjet
D06jbRBclXIjgw6WTU4x3ajZ3FTuYQjFJFQwzhYntfodFuT7uWrCxoEg6TfZQ6Dv
AT14WxsvCl/g+VvrYoOcUq4EVOGySNc2jeIp6W/7tqlZOpAv5/zudY5Bx8eNWOyL
UuDQOGoViy5ScbpAtCv43t/d+OoAeN8vuPYwc9ax0qsm2bhTp3QKcl/d3SToQu6N
22M1WymgcpZudVHs0lN40ohCisPpH0+ztpCnNjCjVJBf3c98OGzQF1Fv4re6cdpD
kiWRIU5DVXjOJ8u61b9uYUPGhXTrZdREJqUm0h/wmDCYJVrGODj4pAgR/lq6jYor
hIEPccN7C8LB2RHV+5DKXQ3hxCih1gmEnAzdUPxTMNMPdZgi9tj994LzNolH5cqN
gt758F2/LCQiR/nUjOfdAitA95D0s9JcfMTxtV0ubH+pTxm3C43w7DLxJOV8+Jt6
lTfUvebZavlsBfHBa9S/WhRwKfaI82g0iv9tJcxpR4HgaotmYpo6KKzIYlriMjVZ
/QBKhaD9Llus4JQ1UtQ4Em0o3jQUhCqim9+Kfoa2m4lOu8zG8J5Y2buX+1o5xO7K
58CK1p1rOi0jh3oZJy7hei430dncnY1gHNtqgsay3a71NZmp/8uKxKGGoV8yNaFU
00GSG1Nz/NomdSMBAlEOoynRwgdNdNTUd/zQ46GFlzq23hr5P3htOZ3CeDPIkdaU
tK422Dq7ZLis0MY1mwdSAABn0A/Eygriz2NWPUXS/cDvhZVyhgdVpkd7UISXQsbG
ejAO8p6a4xmyQqzk2Bn3FtC117zyDMnoRmr9BQqLQx/SHissETHE8IpI95GaMx5c
CG1PmCyPcszVOm+8S+UMvxxLTRfoKF8GIiapa+83RuXH2RK2QuWwrJGL3Av/ieS0
egr0DQEcF8uESG+WkWEFuilDIr7tvfdjYfbsMZvIHVYxZmhSCyX/coS+ICPIm0uG
DjBZzxCWsmNnJIppmQBo7OuilJ1WVtpmynMTY0LP1sv6KlgpU0HkhIC1bNLQTJvx
3AY5MeI4waRflo5GcqoKtCaBMAfRPh2AAomVP1KgQw6iJPbE6wrJlbSkwFAIjrXX
abz38N0S+a3edbGcmlaU4yGkMImzAZdKXaE9JkHGU6xIx4frZ2oa+S9RA2sCFLrA
DvW4s4oW5j4l5qTq/Efaf2LjbNBxm+8gp3TEHCrbM7yHl1+YDTvSqkSKXhyRuPf9
a2vzyiFHdfA+UiMnXRKCgezJLWsCdMNAJFAiuDWTyVdFvLC2BS/IEe/CnJo6+WjG
E6B5NvGx2vuZePRex1JIX4DOubT67ZVlclD6L56El+X9Yc3IbALJSXc89rFg41F7
XU9W76nbhJQSCDK7Kec1WxFrLr5mfu7zg69OMXMSo3D+4Eho91F7J/T9imczzpeA
k4P/TEX5mDF0170C/S1ll4TyLvnrR2vhsn+6oC+imqCVrCIRXO/wAqWdxz3oJgZ+
rnLYkKVxoHjxpnmTpH7a1fSMSH/YTpUML7AJBDNp5Aapxn5jAViMZK8jnmTP/dNV
AZEIc29wEwAn8FB7+VCskA+6CVgqBRN4on0dkY4P8E3Co6vxMy/3hyoGAxn4JLTR
zh7jTY/qs/QEEWPH4hN5Zuiufj2CLpiFGHlCeu2mUQNkN1jlu1j7IMbe+NYFpp67
3s/r9Rkf8JoBz6OqHbakcNq0UDTCzls0JzEMMeuUdDVmx3NCjCIRgSRUEebkNBOQ
aEuu9QPahuOh06KYP86ulkFzmChE882w+bNHQe1ePC6VO6tFq5TMjeaGz6ckDQ8g
nnYXthaTa1FTIjl/Yrip5Qx8WAlDJpCC18mrffaTnsFmehC5W1igq+xeTPRs4Bms
As4l0PelTv/QwUMU5LmQraMh78TEgra92OsjsC4KMRFGRkaLVfcNShoIH9e2YwVf
/47IypM2dJpDNd5ONkymcPLpD229yAquZJTzl0lWbYf9wZGLwvYuBr3OGNtgQB5R
Whs05RQFGqcN885DlZ5mX+FNrntAC8Ox5bDlH8Ve5/mpJHa+Cv8bV24oYyb/wcbe
VqOit2uwuPcokfmWTsGBfdTkv+040J6uLlDn1eO3B90DUIQb9VHU302px0K1B+1q
GPQiMaVyGzaK0yYhsrpuWPw1W/Ob6XTG9FaL4exErANAKd84WtW6hMSGsz5PS6Wt
30SZMXzHnTJ/Er24mQ7YanbtUuakkG36scSWUi6tTKPOHHUv6ejPC1agfX9KDezM
f1edqxQQqi3xtTdEh2+grqt89KY1CPUAjKl/JKh3QTevXX85i1sGcKGG8TotaVjZ
bgTK3LKhIYyw2JO1TbmVF/tepIGMFx4DGOy7JZd4f2IqLkIvZgey+8+irznDFuJ4
2c7rWxW9bKtm1qrr0ezJvyKeDKYIG9+eJCQUKh0PE28e8HhnokO9wJwlW2HHXfJE
O4nCQFZuknjFcsAvCFCkI8tJHFMBI5karXlJiFUc9CBLdoE9fJu3vW1NiXshMDwK
KYQ1ES4zNmWAnsVtHtt/plbv0L3fEf3SiffvbrcCJixgbn/GExim6ezjjWw0/QoU
IXNxCgukjTuOTYw9WoQaX4MgX2QxD0z/Zz+uKhCOv56BDbAoWmAd9OR85F40lznc
MF0+eZcHzwGiMc3xYOHUJOgZ95Aksnh1pPJXWUbxFlDzY7YPVfSHIwEdrmG62Z7j
K65VdIibSIjtic1+Ssfl8QX0dH4Wm78PxWpwW48GgV3chMIv1YIXDI6MA0M61/QN
7tcp11D2JP35nBhSnYELSOHn7tiOFqS69vRVADoQFLx3CaP2wkVm8/CoO5OTfbnk
iMTHf0f8q6BBeAVghxn8Bj6tQ8rmeVsmlNtCE034+7TuXLVH8b3ieKcx4PXRNuPv
4UzstVXmojpmQ/6k4yB81WRwCYnWc0A+Q8rNSTB8799kGOTxRLr4pTWsB6Q0QkpK
imFhPNI71HiNJCXWjz+yzOuHr4CVl+ymxXvMLH/ICOB6P6aE4PSpUtCP8Bh0s4aT
Pm/3DLlWdZK1BPnG170LB9dyS7LuNfUUjUbbgAaUNpAPSUDva2cwy+DH64g+pypn
EDB154X2/tN1HgKUPENOsoRfEpSMCAJxsFxahGYZM/mug6ZrNNSgdTrxkXiix2Pu
dPFbj7ltD04eCIgGMF6yX8DprsDAFbs2TL9QGxzVaQsjfoo1UTGeCOOvtrSKMqJO
gXmY5ytjKfPN10trfujbaDPBMkEMOSrcR+ynovXEsdJuinleh3pOQ9Rvjak7xGrS
Aq/kbe4W3lg7wfno8JNS1r0fwuJjpdUXDcCg/BmFeDS5+rAUmXDc6LulNHBHMS5G
VZ74S3TzFB3qZHMWPwrG6H7ru7ItZxMcEUcZrACXXBSq+lz2iDdWrVoaHO4ngJn8
WT1rxhoJuE8g3twsUUM9GCMDx9BOYn1XdZ+DqDSCAE1yjD5uwITJA4zrjYZckh7n
FpRiXoslk66C8BGoxF2dA1TLIswg7SucMqPAg6UR8agA71XnaJBS92v9q8qsUxOR
ldPrFck+hgtzZxgEX5N/WhQCPfYR8k0lBAROMRNIUCCVqeReon/xLEf4AIpxw4Bi
IwAJiiuFNgk1DkoHg44ghIwgI+fIt4zlrNmQYm9J+lZocVQ7RUpH6yawOWFY37mK
ljvMH6oJWbKH8dNtKxnCZOiaJhyrWoy3nQR//k3f5jUw4CLZ+xNIJELu6S6mWImm
pXThUCipEsk328Z4RYaa5sywCo0yAMYxb7yYyoxvYce0rSEhs19+b3c9btUwT6Af
EFXFSZlxu1vm+mjgWCZ8IbzSyb7tcl9H9d7zgFlH0/kPU3J5BbmgjwEW7bcYZ8m7
U38oTRp6rvEnTJv4U4YR2auZc49DX5hTRALPfRMXiMpn7dnVk4dKd72uqOtJwm8g
5UCKdOAEt1V0gpRAOWfbTsF2fGSQ2Z0MWWARJvcLbuWTK7deUEdwYYbkTJr5ej85
yK68HFpGQQ+O5kqjQPuZNjreKsJuekAy6Egz1CKZUyA0agyo34UmiQ8F2UrxkBXZ
kfPmGLdW9X5j7l2n++jNzq3C+UUYLN6PNBG0a7TWnSaH33iMxrvp+5wkBK6Uj5kk
oEV4MiBN8of+A2NOkqmmdoNoUJhXk+7uK/w8c8rEfkCx2TQvpdO3JqK07z+XyLVp
8gcto3db9dZa5xPPaSSYWN2/JbOHV6kPZlOJyEZ/wWL7nyEUMeQukc/sBOAMTqxj
MD7+aUTq7xhiuzO2fW1E/ZLWqX8+a7QWvMqjVVrZ+qeGP1LXOYidgtT1fdXPnkfE
UL/BPgT/xXNUcA4tT8bUcEeNH3N+56jgfhZVM46RV5oIZW3Ie4ExYCATQGkLT58P
4z683QzALuccnTjyFbBbmenndW3PBRZOqvKWqNi+M+Q1zvtHfeNAF5vAy+SsQXM1
/6Nou5bwkx5d98cjIUkdfWV7IFbZjexrPBFunmDM6yVCQhExwsRdJmWBu1V++hXE
FO+1RuZiqGc8B2c2jT+rk09tw8JeTimdprMsZUqnruO5+NB/Zrq28A33gPzOTqku
9nkc5aRzyLXezonD+bb7p9wgpA7fHeaaKBzuNMqUFqYxc09Qd/BZEO+7BW7nY31D
Q6lWXh90Wjp258j5XLiy6SxEB07h+15X0muRw8kqauwG7g29/gDFPIuMIAxgpH1c
vUoqOPUYiMRCpmFGTaEZT9vzpd2ryFK15JVpKdMErtOMnbVaPkcYtJA/Seg0jmKN
UAa+C+gCoBOMl37h+gLf7+fYMLNDQjrF557S637MSmzSipTfX1BvzYyaMmyq1Oop
8sjWIxfHRT/wm1Xn5F9KInNrYImVTyv8hSgRP5T0G4iyF3iW+rUZ1rQjIhK3H6L3
/2qPRpccGVkV9tIeFPVYsq+2mu6FnfNnBLz5DYq/UrAHkhRxPTOP5VEFrNX76w3w
LQvAOIPMpKimAbSVv1SFDnpfUWP0RuBj0QVFqJrmi83DnBCSkz9R8MJH6EeHeqMl
A9rOypyjbfWFnATDGv6wgJR0E0aRYfc80v9iOvlWkBu+ziSSZ1r6Gn5y+79ykTbH
aBibkazuWnmRiMrR6eRo4J3lvRWAQpTDrA1tc/is4k4Ujw45nwDzBajWGvGPBT5K
NyKXGtXzjf/9mzyXqnVifwo4w8dIJPO9it95DUl9uectBzcOz9NkSXojhNVZzn3s
EGHTmRK3ow3sfyRGLnRQcl0zj8LFpLccqRNL6CzVCoil0zZLPP5Qyug04ukoK0Mz
LJGQyQdIbYGZ9hg/TSe7ywykQn16NgtfQYuXIEMA5RuUqDq86mLusZZqPuJUq1VX
gCVUX7P1ydJj2mill0ejLhct6Tb+GjxKB0vOvo//wg8OimYOcv1tuhGs0puDk1Rk
y72f6JwO35Pm1fsDuV8s3Wz/rbPf1moMfJuOaWwP4Yf2y09Q3gmROePPEgKpqPEk
q0NL98NPRCwHW2ZNAj2fOKVQ/rI4ovIluX0Cl0vvg/xYgJmJLiDYaLoat+LAWQ1G
NR2oTAeBQmYDQ3/3FW6jFIxmEqahIIKAFBCvPaANqADNtNKC3j4o0oxS4c81Qx9Q
McFUWFkV5Qb5nHeFxJFSthpuPhwdCLE2qNpQu/GOcK1DnQ2dhb4biHiV17+7Zhyr
fU4H1JbOyg/daFqCLn6aEGqGeaLiuBDBohx/EEH6nCEg9Cb0+JU3RZiadm8Li8gJ
J+DL9k+XteWDDZwgyunz4L716AxdpVdGaXTOQn/jeFDvZzwfY3VDkfBEtaTQswMc
kDw/pNXCT2Sw5E58FkDJoXvxkjGIWt4LUecjl5r2IvgTBZOWud08qr69kpvMoV+R
5SttwP5utKK9DwW16snZcJ4vrGeqRBCd6l5Qe2uxgd3K16NtsldiHB98CCfaeXzW
ReiKonn+xzBy50qg8bGy4pykSlil7LuTm8wNlJ/vXrCXHwiwWHfqMbQp453CFLYN
rxZynLDg6hfDhfiBisWIcqVqVdEjStV6MLWZV/89WShE+i72lVPKdeKM16eDrCOX
DZGz3QL0/2wo+p1vozlKjXg8BasIMY3ObFDuSp6zvD0S2vMpE3X1IcuXXudpjFN1
6uTEvPx323pJ0YnpiI4uKWIw7IdCx3YZjGgVeWuJxeoAkrACoewuU0EuA6lFKajD
Ej5SHyvx0Wlprj3Do76NlD+sKJUjTrksLjLSfte0xoxJ2jQ1EKRn3kleJZS1T7RB
dj/C1kFzHBTUjhhEaCSkdI4VZGBwv+sKrmuuz5oghRiAry++/9QRDfdbVKxz5nAJ
xIsThzIIHX/8Qa8oKVc2Ms1BQk6USiRaNsgYM+iuf19pDE/oNhWGNmxea8GQA+EG
ColUlu2UraWrkaKYJPG89ocbTugP1RizxjeWQ3++rO7HZ4kFJoBieJEcgvq/DtPb
iQ/fLGpbpGl87kbJt5uoD+QFouh7U9KEy/8uMccNUpRn2JRVR/F3ItSivW9iswZK
DVP8lNKJyRXw2YriVovPaVUeZOoAAbkDP1Nf9FHk6ryN92vkHXZtSGN4XlHkHgUK
VPkBqBqpLadJB7eb8J1q3E2Cc+MAZQlcepaHAhCHhsagjRXXwbs+UhF3WiBI4Uts
ZT5vHwdJ9KTKhWLia0RsDJaBl4T7WgHABPjSvKgwPYiTA0QfgsIndtltpNF6ZjdP
wPrXZaFVla/yzURT/kWfHdYjIPmnew4wrtdUHtVrySAWJmdMtbOru/VOR8AijT4p
Vsh5Mk2Qw1sm9wJwsh3eWeffLoysZhom/mSG316i1knTEoorvWKVtg3JfsOc+tqO
+Lb+xroqetk+AH7o9Dj1ES836CCfgYZheumSAcxAPXSji98k6cT/uGxUtrjpm8yx
whIVaaj9AcQyxfPXOTOeyAoBWleBMOM/QYJ2gYFotqrekMk1E6GsEmVn71eN0573
IC0drIXjSoqONXQGYbsGcJ1f6xNs8zHDuXtFMPdqwSEs93W0WeialdyFNtiiStBe
oCzQWzYNWQSkPywmIQwK8SRXZg0OGG5D/GooOO0Ub5QT4IiMQ80ZlJGTZ8gzqOzo
ViSUJ6g6JBcHxFeOFvK9lnwq3mMazZlTpw7BN9JOtvn848X5KPVXpgVT5/K0A55B
85ukAYXVHmskt7Zn6AOZU/qZn/+k7rj/qzt1uIl9MyOz3KBTdxUZ1UMC7BaB6woK
XrKUBKc/n72/kgdWbgS7R+A0iblQvvbSs1C05lLCe2o22mjV2DzogfQkY3mcSsUa
1FihP3J5lvtQh5PlhkCeV9utctqgBZbOx1kUkOTisB3aeJFPLxHvc99EEPCkGf0E
QNHi3whpFLy+TzMU3nDFaLV5C9DlbROUzU8lq+hwQlTaCCE//CB8zCoHnoX2Jkvc
nLsscAKbIehHI4oSLmrzy90QYGMUzLog3SHLDNM6qq7IO+/J9bbMtxckzJy05cPK
h1d68BMNycP//bgD6FquAxHyukRZznPOV1YCIdcplezNOSkTL6UHd5WL6w75nTmw
hQ8cWDwDHqPWnWCw7ymEOsHyDXkgZCgNVI0nXrAW67TcoHz+F5RDcY5nb4K5kjQ2
gjRW0VDenCVMxMBXcL1XoUtrN+eleBKVKF34Sb0GFPT0e3f1UmkOWF0WC8ISN21/
taTQVTbcKMwu57TA/szOUnysPW0JokOfZUgpUwI1DniB9sK3hznYg+zKIxYlbCW+
OzH6KwAanRnH0IKSPwFgeYgeMeCDO3cf0N0U9hToZLBNl1qTtwfOGstjw9eBCDIy
QiUHAZCni1z5XqlhtdNVHSRk33cXLBKJKO6Tpr6Y9lSFyZhxEwKL0SxEzW0nyAw+
Bjkryj4LAEd72ZM7Frq7WJ2HTmfS8wut/OvkAQlNGudDmCsvMBXEkSJLDe8PA9Gk
uAWUiCWQJPi3Nuvn3XFFDr8Y7A755RHbCmQbOLO1PGf4rBh6OfPBXN8WsKHMbuGU
T3BKiDy+Ls88nsBUOSB6TBJefqQiXVHGfRiIWWgeTAgx7qmRUL9xgCV7f0aUR2/z
m6tQcB4H82yNqgGWJHEzWRFfWjuxKqKX7921GB2Z/urDG465kS5/NH4ZH8+Bu07O
VZJQRahqdkgetZqn3OvxePmMFNoFJPP1rRJCJphfgOqWBTapLRZ5+YwX/F4e82Tn
4cIBQw9K0AmeuzW+OTMIDo8eWckiQLELA8lix5BLxM7cu31OKeIFR8YpN9Iq+Bdw
uOMkAJdU4NqmBRJ7nmUL0urEyBC/8+cz3cWeufygwb+ks2icrbuoj8x2fCWVv0Xj
30VVrqcW7/P6Wrgpsr5Oj90CzqoUmD4cZKdmMLxdDS/EvDX/8AvJAjlzjFKbjZQU
cvuzVCJ3QBnjJc9BfQWW8Dq6qlLYXVOXSw3nmbX96tKwf+BFkfmMbi6JAtktrODP
OCLolxwbZX6frKCEHZ+pMtgVO9gSksjqqwhr1bkLSGBeN+6QFsdkKGrsT2jR5VFy
RlpvU4v59zwjxUtjJuQH9W0R5cQf0zKQQseZMDeep7wNwJJrqxOZ5oj5AU1zYWe4
Tsp9ovd40+wmvsAvLRURMldVh7YhaD5SLZdTfOKK1IS5RI6lXiN/sLXA4NLPWMWk
RfSKqqMt0COzXorvm4sVOCuULPX9J89fegwRt/pLFlmj1uqCA3hbGzjvfFDl35cZ
6//6ihZs7wz2xOLZZIhRAyqohkUzqCjKoILrKjS9bqYICza0By9f+QIgnYqXbfXm
8nxc/Fbk8BZFumu6OzMAUbsJVXcOtNYHUbzXcoCbb6NTPpVo+WxEzT4OPVIxK0E/
RTC0+aA4KtKAyHrrUekWBpezDDNANFvD9DmLebpnlNo1Mg0zOA2YoHIsfa5E1UoF
G1STEkl3Pyf9xCqkZvghizaDD6Jqq0wmv+1botJk8McID/79Jph3OUPaacpWXdPU
vVZYd5jxZN9WjIz6LoF4pn7q+GYg0psVkuZrefEtHpvmYayhAV70vcHw8jSYe47v
vajvD1QpmTQEjwXJsiST2+xmLxLF+ktsFHkiqpXblPyzBD7J51SgoFRriyWb3dlJ
8BgjaAKXnApJhiCO/99kNnejlmvj0hi089uVRI35wl3dOU8BgHcjqqsTLb41bjuy
gh6YIDzEH7fsvId4+ACP+CtmA+MTqg4FB8FKUtLiYIn0PWFx21ZPxODfD6xb8tku
ewMo/90Fgzc9SiHkPy/ALNRgNzj2pgor45Mp3abx/tIJm+RHh80KEjNfVVjNlqKT
a8IPLOWlZq+8v36KnGzVuEZvJAb2ciJToBXrrpZnRNltPUs8ptlRFYO/XY1jj0Y0
T9J/2jQn8eGMoZqQDzzZZV1kwjZdBokAgxKNYOXNFj0YE8cwkjAapo7HL3uH9bkW
dxesxYswUTPv4zsxgMsKePlrDkYAArEwcJcatwOBaYF1R3m8waAPQt9RrmePOl+D
r6MlFnFl0EPyXfkTLNjk78QC2voq0BjCGKC2yUfUEGwV8CLnn3hwtfYr5RvAx5wJ
5QX1NNjXFiYXWjdhTr6UyELRJIuU565Ubpv2ytEQjnLYbqTaXrI6dUICpMUV5AAA
YwrnE8scwJk8QilFyUAI6DP4NqUbxjfcn8f9rwl/4NWYcqQ2cxvgPVCXj9A0RVlm
bvgCP94CGge992iJiQW/NEac2zDqG1rrq8aDorOLWubcEHHLcwZbPsrJ+6YCJ/7D
QBeRlI+wlUq1uMyvUyUQp2E78Lgij7f3w+1T4DTNVf+8axatUyabx14IC18ifQ7H
/YTFoMIVqnzSKca97WTCLdDbL0Rffpfeo496j8T0DxGCb1LtTC/YXaoAwiwbK7mH
9+prMC/3J4W3GsTD66Lp0cjtt0m8N0CoN24iuytbs9D+6F3XnEzIAy4cYELDTCW4
chZUPwZijesXcSCaFl8lUaUjdn56RKN7M3GJItsIS3ZDmV5mqOwWlWSAcurr52Sb
EyxE57qN6CcGO4d6/wt570q/7s82KE1LijqZ8E/oZbx6ZjbY8g8yQJko+x+M/F3a
/fB7Trr/g1W4lz1tkOyUMke1mqfQaw2W7BoU3vcn3hnRmRe9zeTommDKa04d9/wA
SDkIkhLjYJ1kQ2+FUvsUCJGCsaPbCDMQ7KIzasRYWvnwzKSOxAc1vWFSVJHaL43L
HPkO1ORfgSSYllZIV2XkeCXp/7+KXLIP2jE6gNm8H9w4/4wCRRRmrOQ3E8G0q9y6
vAqb9IadLCATbMG22ZL2qqS9MSk0K2fx/DBKSlZWGNg++8350JZhNi3sEM7VgnqM
Hjw8okX6Nim5IuVNJ1LYy9UOAndyY/eu++KPIt0zTvh9YbALZeWs0QcA7H99NdwB
NlJpSSqWNXcCELfA9EKTzclutHE+V2EtGJuXBfAkHkAjETGvqE1zZpCo8JHHQdH/
5V9lHbaTRqi9ybcfnZAqFOjlQrMPK25rqrTruLPgISyrqNb5+3xW4JgJoQD0sVaI
ckQluqAIj+5KglKtpa8a7cW+/treRiewYsRiU1Y8j91odRdSmBiHu5V7YinJXbWX
1UKdoSwNC6WaQFucILrsLGgcZ0mCC1qmCjaNX/1Bjw6qsTfFsZNRyzItW14VZ3uU
+m2h69WBqD5VlZ4HiMJ8lhhtD3+/k5vGJHxonI9HO3Qkcadp8ai4tk1APlCvmeGM
ZLT/7GmkFnJaE/7wstUN8am+SIQhMZm2EA7048dgb7vwyBNwaPD60cnVTnuuJcsi
aXIRhkVwKrEPGMoBa7Lw5tit99rcEI8gVCauyQSaOUjgF7gMnQC3a/kMW6V2T6Xw
WgY9cTDYZI0As08BSob6npv8Atpie7QxOv1q0rvQLxnFD2qk0TMElXh/ZgkitrdG
swqoLqQhIbvfDwyhcZWYY+DU5CcT8SETkPMd181VPt6ItjjpLD/BdHrf6SHaI1i4
LG2Nogaa9/VQunjjrzzUgkZjDQQUtk0itrjOZHE9cv42Aqf9wzKBi5ZtTzftpQYh
FAFGYQwNjfxhh5PSkQ3dIF6xS6D9JBCLKDluzkDAbDatgO4r4CCgPJNOWCvIzmRP
p6omihe1E4pC8e8fCiWGBojJillXieANc6zjBufFeac5w8xej13/ulkcNW1AU8dV
LZQU7PhevtwIUhFkhl6iZLx8/1Ff57HqWaJaxvMDwnfUGcFrNs/BzWPZ3PlCbutv
A27VNfsUk0hjS4TzZTrUY+0sMQTu5+SY6XUBpV8ivqc4+oLiSmARcdt1aqmelDWj
q8vt8wej8OkrkDszg8Q+fBVvcdI5r8gkJ1JFbJvnFYUcyuibgG2JHoTfT14gM9tR
SfarksFkP3/LIVcTLIbKmXYEcK5zbqR8A2XeSyzXw23KcEgz55l9pGuxebUe7XUy
8k5rPkQUKT6LTcnTTG4hKvfvWeBmDiqlG1hnWxd+9tqrgb6UvM8pDITS8C0g/z47
zZ/mIZp4M0SYBMZyviM+vLXMzCj5JJVNiu6Y9+gUccLzzLxag1TxwgdVJqI11I0k
IJrUC/y0onlJYkEJYd68QrxVLcfcAQfRrAwVLMyRJUMuhxsInhtFN2Q9CuZWSGqs
6HrrZYjMN3TJdizMeRFTDsDqdOYdZI2NGText0jLTztBgiDfmAZXY+5Fyr3Bvruk
2eRppw8CcGNpvNz95yYWgbyMUdh+nzwrrGor/8EjHHQprb4xkCzzTOd1JNBiMLjO
1TGvMNCHYqYprmWtPvWxWKzz7XgCTnfb8YQqhYxx+lP1m+buE6HYAEHoVJytLC/6
q0gfWlsyxjnoymJ2xK7HnHGCuCJoeiUzaOoBg8/L6pGNn/FuMIclGpNzRMpUwWYX
AvuIEgEcRbO7DHRwVrrPvatN2Cpr99IRZQ4dzaKclCP+jq/05vada0rCoaZLrA78
pktIHCAhzp8+l5089S7s6Ce/MpZAAA2lEAhcqm5HD4/NDvRqE1SCfsHrEg0wCojF
MwWrJ6kxFS/0ylgpeaYa55L4eP4AptObw9lOq7kYVIXcqzsicI4vkvNeElnJqMFo
rc1Ird4ffsOaOHvdvSP3G9f07paiqsT4r1VYb7TP/GlycTZJtExvJfZqnyZBLfSr
1f1eVzmtSw7tiO2XDZaKtFLES+onDip4aUfuIdQgnaB4ZxFcqH+RLadqXrcMmB80
HR5TFIgmNKkp5lZXI4uuMi2ZiVHuXkv2OBAVWfU/h89pNailK6wLfSSm1EZJ8iEr
47CTfY6f6XlRhZ2OcNziiYjnJbY9GY36PHa1+/XAGyCMoN4f86b2AwZwxGJM2Ha7
ZDQz28O8hbUSQEtmCzgbpYh26w5HlqsNfSnI/hcoPMKqhOh8KTtR+wLSq45oow8h
h/TQIxaIkbzc0oCeIuBaKerQPnFXPbZBTO7gn4VwxfHbzWHVyrLzURLIVnAsTP2P
CdOMqjhhEEVJacBb23KKhEF3R8qINJyTAKqfUf1iJHS/sKFhVGfgXrczvP1Ovt9/
nBhlXt5SC0xskEKkb2VnySjaLF9lPxOK16nkkc7cL2DBn8oQboBLvEqWBXQ7kJ+0
iyUhLmt6Oti6l31YDBBgTxl7ftcal6kGI8cvMLBeXO0mc6Y8xF3aSw60HzCby9qb
7ZHW5HY7GXu9p+NEg9eivyLh+bqjqHr71D0TTwOEvHZS+MZYBij1tylviwZb0eja
Wgzw1lbdpX/UAkr/ek7Gsw6gvEVhU6wAM8FfGGe5v7vQIf77PoYMROz1IP82Qsvr
/qMSxZGUfl5GxeiH9cWwPObMOgyJFhoD1YBDg6NxVxMSGeNRFB7dsvp+DTouMxPQ
6l9pJbz7/3XHOzt8IJcGOrtrXtTnfCgR8MHQqj9a6mmmkQlnhuWJw/zlAiMxAwFD
Me2G0x0i3KB/unitOk0/XqiObtNyyQFdNth1G8W4xl4xVuIjbN8jI/dYSJOW9nnr
FXsW39EoI5dVKblRbNc3sj1kvKyiePKxcEtkj8dUflXRsYS4ubnGqDaRMKLWp7le
6k/FxxcOq+Cht/PgHrgt/5iCAJ5coat6joCkoDTmgZzOHeoO1/X7HWbKT+Ge44Po
AJexgITmoF1YKv4Mw6wPNgYI5yAPL3LVpUyRcEmbFYgUUXe88CkwQGHqPrYDYPe0
qViLITSzgI3XUfgOQqawhfCcQJYBYYqMztf7c+GmCT67ESdkIK4+yWXktf3CwHzu
oP0226jyyedhjjgay86WXq/enIV+O7Xm4qdgzGMDZqLcJwxYajdpSikn+hAKynG0
/WdHqlUjEA3P4NfZlxhFegSFQfa5NjpFv7jI62a41KYnMqfoi/Hqngvk8iPX1zaU
mRtY+Q/3/1blTLNsrOFKyExkKbRz93yiURFrepu4auZ1CYPHua6j123hejp00+oG
7efAQs5Kt5gEHihcHKgdUH5NCheecxkeIjDZqmWNcBEsMRSthT6qmoZCHN3j4hBL
+3KMcjYPMG6HnjxseRf5JIt/lPAmdM1SMWS4KBIRfcMCH0gWt3hkw5lh6+34J7Ir
kdNatuAkqpba2rDLf2JsSRWTqibEm4B4lSFZzuYoxddPmWqCNA6jo+rWOvJC67JV
mjCKZLVcRitFg60mJi4hIzHgbjoslp/jAeNo4+K8XABcWLoVg7AfAM5V+/xMBolO
bj8exdlMPCZpphf39CQ6UjD+2UVkD+4/VNKSu+1Ff/tELnmiLYtAWq7NMvAGyG1J
SB4gn7CVH9gh4XAInjPp1+a+JNEN6pRW4IPT0BoS+XgvZs5PeatT4lHp+tV0vJRH
pfmdg2i/EAgBZbBf47f8N8jqPU9mGCcY9k+SvErz+GaZlOQQu7q9+3JyGEG9Kuhj
cGq99f3TvW32zF1JFPM6Bz95EkLQTRAt8Ezo9b3VZiW2IVFuzVttnVF4i4AZQp4p
t6VxfbvCHsAfZP+CJ/YR4Fk/R/T/xO0+q5Ljnx5jDtp1D+IuNoSan456n+lwy14W
PgVapmFb7VYStQI5u7nPFYbLCtEX5kUwZD2ykHqUsNUe3uLUZTM/3RKow9NimOKm
F8oDYbkMuJPI19Kgj3a3vX93tw+qkGPMejbqcBmwUxbnJrBtii8XKhcgLdvmSoeL
acn8ITtQZCbVnP2j7gclls/JXEz4UFORLE14fSdS2G0cAySXSQV2KdfLe2X+saI9
YUh2rjUQ+q3dwut7IttKD8sHefZnwkFT4WZRtjBE74019cSuUesjvHyADaHoq/Fq
5/MLhE3dksMhylQIwbIEDG4po2M4fpqaQJo/zkcyJFCt4jeWCKdBRoqyLVPn5zaH
vCNa34hvUF24qTNERDjSSmtYpMBwjqb/WLVn6Y1V6u1KpZHrOuN2ia0BTP0UGyIT
11GglQOdbdaDp/CHyynsrpk7kl02pNOIt1p/ImNHOyhileg77VLsxy0ATnl/V1iy
GH+6z8Tqje0/NqUofOlrfds6Be9w55oquG5glt4UdzXmWLfFstezIsMZWiKn9nGZ
Ht/LrytZogHoCKGkDMQ3MrAo0+9sNASLxwb/0We4HYjALCNBISGKOaw4MlNqefUG
1+7t/yw92vHTMYtFC+bLZw/97ObIo7SvRiQOVkdncR2chXBDR7Z0AeLAPkAdd2xC
kux4+YtQqycbJikua++puQdy8JmO6g6aIfG8LzWQQDLLprIs5t02C42BTHKE3cbE
iFF4xmVpQJHsaIbgY1sbxj4f8Jk/JygIeQg/QY4/pM9Beunt+6gIQL8UgKpDg/0L
2WoNJQNo4H30eqrGeZq7GPNfJl2M3yhcx1NH3HOpj/j2jM2BRVUNxl2eto+mgNo8
hP2DjbVgbDoREULDEQ3oCi9+QQJNx0vHN42Q7qetn8yVQ/i35xbSq/cI+i9LkNxD
APxmjxynyz8mZEpYQ4yTaFtz7FflUxqQoNhE94Avnbg3eQo5FPWEkEgRfzwEV4wl
Kr49br9XMZN8AIDnYGVSlC1QLq0j9WBKbHeWpP10jsgD+L2ymkSzJlltxvcPEx4G
8K2pn856AJ26UkkvjRsA+mIOtjNo9HWdpd96Xe48T9b6gxbMpcJRYqLg8eeFV5F9
RJujQicJwFK7We2SDfxvunLPCGveq3vRgu37nXghtzy7j0YMAlwInns7nEtMHSMy
cAZZPfEFjMkKbSXhIfcPRTyRPij3wCdkOYq6MGYZkFMboKVu4JwZFpe0jdZFQq7X
plOGHt189wKJZOjwl8Hj8mDTPjMHo6ZhnqopdsfJ1CR38xC7B2gmTEDqZwOMrPUw
ZwBrYu0E0+5re9kvmu1HlL6oKvS5Iey+Vkp73DcD2LVahpr4Bd+wAvq+khZ54Awg
tPzxZVNRG0KrEyYZR79VcgUmlZtDO6NPVbYgDaeEGAHQ4KQMdKZoa7TyOOoMC+EU
vVFiAnKWFHtR5LwHbOtqcRXSwNTpT/zbRioyTmgZ0QkazwL5P7MxslLmZHoQADx7
i+BM9/LCGOfu8yhEiA+08NzLHPnaUcd0YKn7rbbHqKNBu1SLPc7OQJYvZuEzAobg
31PK4XaOmT3J4G/dI3IWzmznsT1BGeltOhbqa2HBMzlX8gmp9t30bXC2nX+Gy+8y
iy8HTtnU6msuK02iMTyHMZtAKUq1KL5OAzOJJA4J6KissMKWEtL0siiCRq9dslOf
Elf9cfqw5f9yAR/GTOnMEB5BpCwsMoeuljCIOav0vzaCB5eY2sQwOMiW6Wo1XCi0
hOZ4PP0K/pXiC6TP1Myx5NwCRIdb0V3guFR6SxHScvTG5JQ5aQBf8x73dQ+wF6Fq
DTevEii0npmdpA5DfaVIVBdNAZQkskZM/HnBZjiTeBcfG3EBf7tWxlijeR7IMwQJ
MvgLBehdb1+5Uadjz58ofPfzUccylh9C5jsAAaTYtMpNw9R8rgNDSTIvmlXeHQTF
QT0YglBxjcCITn9MBL/VO943nkE+SUr3wnYCwh94cZK//nqWEjkAN9yREF36vq6p
JRvtqZGUbfjQph5v6yN6kaW+EEExMS/xSqD+ybhAD18SobI4n4O6TLyXBB2gDScb
4xh7amtDPai96XvvhGvDGsd1fVbcA8ivUJnUVZf/Sdo4fcJOm7lm4W9wcohS9MDF
FFn3anCoGpsmF7WOPVoBYwbZLEXLUnGdyPDSNXkAVUitJQ/COj8zNfxvJPSRZcGm
r8uI6/kEm4ukavqO8yQlptzscvvN8aFtLXGCxAO5tE8PgjInx71i9dqWZH0ccQ4z
MMGOovoP+xnjwv8FN0HT59R/wZJ7qN7aqu7HuTjVRMkO2Msildlb3RpO3PJInX85
VtOC6gYwfTLetg7B6wD3h0km21Sm22YQ4vjAQrj7hBc0X0xkus4yAYdzwJd8Aq+J
yTJZ7yixNVFQTCD6WwQw9KCeKVXrrKc7A88FcIIutpA+wiRKPNXrxTnnX/A29EUd
UCO+5yDgphU/z1Bm1vX+WUOZ5Su6bM7ejxbKi1QjMyWx+3C+z5e9Pc7NN6vjfXNW
iT+YRv3CbQmeZCswW1o5ZJmfaeW1lIBHPlbFoD+p3zDs5Dzsx7Te57SWrNO62lGi
Vc+jFlCfI/tp/dMAXhUlvy08QsZg09Q5sd+hVzGrK/0gYnKOQ4dF6QzRQJEeXBK+
K9bqxpAfl9l6lI7k0fgYIqIQhFkG2aYgRyozY9ciFM5zkh4RPlWpFTjdmP0hW92J
gcZOsIvMsr11i81yyp+LBxY4Vxo39qVRUJZgQzg2E+bhH/FeEi4i9ykHE8LNlHdl
S30gbQxDtU4RlzjGBOPdGCEnHQQOEeTJdaG3hFdOuDWeakCdPV3vGxpL1shZCo22
NWDcCYZR8CKLm8yXcxsT2iACOdM0WwnJATADQbsuys1BJrOSWG4FBDkK0L/Li1RA
S9tbu7GvQDQfbMzZxPeAgzoHMWpVMo//9VqIZ7hVlqLYo/xUW8gcmy8xcIzy4rKR
+pMOZASglEYcQXuNQNgMX1eg5Lq1fQJIFhZRjm3UoiviD0vUb4tVI79ovRTuVRNE
jCq3faJh1Gpl1iKspJa7SJG8bIlgx+lp4RemqBkBFbTWUhzJx/9AuwXcLCbuo7mw
e9eN6YRUqk8Slc+NtDNaxOUpdIaTX3WO1zt1uIVSouHiZQ1mnPVrKaQKdmapJ58H
VVb/t0ylvaqlmS1xs/CWLxwsZkMGJxH1zg1BdADusieMeEDVmCtwrkK2iq+6cvGV
+vG70lS20+UHtYYUmXubBtnJUUYCP2VSm4TYpGjiE+WQOliVCVqMAOUTXzoR7/xX
mPim6cT4RSQOEMCTdx6H2veGv5Ct/KcY7+IbuNeHMd+tQ6JVdkoZSV9XoZeMXHTT
dBqSG26Otc5D/li1IHkVbMlwoGMMpYn47xsROgJxuuy0j3LR/BOnyK/aEiBWUT4n
7/IYF0HZOVwbpZHiPKXpJ3tVGj43F16Ms37k1GAy7Y+MFHyQKgtUqHyUt785Ypwu
JP9I3hKFTAEN7RzKmEuiPGzLB7zvegjNjZPJIwtGCxSYgdi4WocM59tSPRROMt4Q
dFkqAdo+0CDJeMKEeUrCXm+izPr5PDqk58uW6rJzrgukDpNwEn+UYDHU8L6AJ6h6
fzARFcU+wvylrXXfsMqQavJlhNtMmmvXp3w8RInP3z094UMcaSuCpF6sRMSWXpQX
CTzcVMtChQ+mCFAp61SwbZlkNp3dbQA1EBsndzM26lMte13E2IUn3nN6amlHSjDK
sjNQdaZSgeSW+EN8kQo+DY0l4hi4cc2iQ7tssXmHVNNdBCYniCH4EMXgtqEuxfIa
SihajrlRcA48RmfVajq9JuhCHYk7ueZyUuoxxsvsSlCCP0lO7fmbflpM3xUIA+qy
LKMwpnTeYepw1rTSRWCzcWYF4Ou+nNnPkhwcNIjaZRVmcapUKZYtdX1Y8ZbdNti7
BNV+4MIiBgR6iI2+WQ9sOmc4ozt+TnA58eM9nvjlDzGRbtoA/kDgmpkQWQ7Y7GUf
l71bcwg/sbDpRSZTBh1HHYrlCy3/bSD6UcViA2XtdkEaktTO10gT7mzYeZ3EUJjF
hhPX3jJBgaXw8jTWPTEw3ksuYSzBVmkTZvH4MJ03Ly7TqsIjrXlM3B0v8RJ1yeAK
53mKaaTF47XchXYuEy5QSNyRMeUwGZU5b+X2rnw1yxA328Z5oBQ+4oNDCfUERPbF
6xPB161GX97KvbpPQfOIjD6rwPqlWPbz1RGLUi+6B0mhagdrCuJp/LXVRe03V0o4
FIzYQIJqyIxYxHnJMYjX7MxPpLoySvcE7v35BuIPN+aF4aOw3kh0RB/lOCOnSS2w
hfWIz3r39ZEGy9p8C05XXAeWcGHo1yh1osKlvR9izn8v8VTz7npTtltlCxcbcXh3
0zkc1HybclZImj1exeA7SNjlvg9g9r8kTZEM0vRygKcoNt3TbxH4NTV+C60bH3rA
M/aTSw/QyDwWvcLklpl/cR5+Ii+q3TR4BZOH92QBLmTP91OmIEniyQGTGTr1HcZK
ykYC17CVUOSPRMDLxcqZRYox085mo/EcQ1Bivp1ncjFLoKdEm54RxuzzKSxDA3Sz
weruyO0EELImoxynVMb7SvMqYwPTfrVyleykqAle7wDiFeIUIbh9cdjQbB/fMIlz
Mi7CZdN08nJh9saY596Tziv4ya6NtQ+mjqBzi1iavyMM2n/u5r7zV6JkP3o0lVqN
2LG/y9McWHojkYyCv6EssZE5fRzIT3o0m5MIvFUUFLPo+eAmcZ92u9nvDi4dcOun
qaX/DNXrO4nKM3XYc9EY2lq8HePM5CPcvpXY3x/JfA5zrui3gRYyOlKgktzZrPs1
GAfR+ChCXEjFkAgMjHtRYuWUdNeBSyWFpVIKKmj3/WqPN8qrAn6wz1qctaLz6x31
0OG02kXktDd2+cX8ldHfzsBO//9St69Zk4XYUW4z1QKz16zQ9bHwoFHVcyl3PUjQ
hPn4QmwakZjYjbM8rPJ1m/FhCvll06dM4Wdx+jUtCADBP+p0vtMmjxD+s6zkzcNk
BzuoryEE+mmQQj1iTj1Bl2S06BvW6MYYqENupTEkOLWI/htxV9UdSTNFo/wooBTi
PyUMM+dhMivj6X1YMnSxcYAX7kHqzLzAxRG/X4RAvO++tlZUk/0HOmknOcJGVnDK
I7YjfipR04JeTwb5CkLUmXnSwl7Ht2zezV7QryHf5aFO+4N7Z71p1VEILrpl2lUw
0nkNUtoG2fCAv/XiacsNK7f/irXkrKewZUl3evkmUkEdZ7AbU+DM8ZNJckxhHmT9
w+uQLNa5JWiaRCDH8a2Wduu5jReTUSluoY7eUZ8+pM3DIvm+ydLJ7x1rMxXwruL4
dLA0cPcGSJEDE7+Q0WJypkoYjyooeWCJxA5ID+1SKuUaK6DFcuxjRhhHDVwWxb0Q
euSuldFAqWTy36zIY6pdGmFyQI92zIIK39zo2LW8a4yolb54xlgqH1MPo4EgR0X0
ixWkaIYodPRip9k6Tn35qDKa5/gXAhousNx59067l3w6tTYtoT4EYT5ztMGVldtg
JdgzJoaqWIoAbi3ryr/hSlKMku7rj7Jq2RelcEIi50Mk5j27E/v/4C/bP7Z7VW/P
86AWWYxxSRkohINDECV9s2rAH1KlbZU2+eVQOnWRIPsDncdQkEeaZnF1hSCwL4NH
xlEr9pX5T8qYSXZ0Hys3bL4b9y2vegFM9oU3AiNg/tGxkPtN0+82miomSbR8YfRG
CFtlRF9Q7y0ZIk85WPO9BTzkj5JxqbBk0qiUxPBeK49zQ6x0UZkAdlUB8lnMbVrl
20dCQki0Ujtq8ub29NUh1XG8mdm6PsypTl6mlCTPW0ob1+u/Jh52eLLVosbUMTyi
FQFN/dM24CWyFfYpFMxVi4KVPVof2s9n3FubsxjSP8Fj9SUa4NNmC0rU38gK1AEW
BOc7JUVJbDwEO8j9/Tjow8ELShZHFE3NhuozCof6/TTbeQHJo7HW+COpxfb3Onxm
wPxFwrsqExSAiu8KNIJhYpYoYMNka6bU4E+UDrEN/9QTqsnPagrCO9XMPxUlOima
tPQVz1wanRThpuH9GygXDuWYzzajWqzpSCXvrLlus1dIXWIvSvkKb5FgRw+CldkB
WLHYUS03i4uPmxK/6o2YbiNtpX6iyMVOAAGi595F94bv4zmGj6bmhEzOedlxEckN
PXJwboSdJmO7zts1xeCs0O91PRlrZl2UYSKQ2/ULv+eddIHv1GSATt/SBK/tcbQV
i4AlRg6mHmmaI373ZlxInfGDXAOl/rdUXl5JZ6C/+I31X3zzPzV2Q0Jq+USMkqph
r/Pyz00oAzoL26GwCm7EXSojeKsm3/8dqusx35PV89Ds3BTXJRuQMFFdZyQ5dP3N
evYYS1jCDQ4rMiTGTLomdfifuE6E5TyQX7r6KD/yoASgVgeOr8R7pD6vs6wNZI9O
jFWIRXgPepDh5sfxWiwJ7jOrJjePUNo5B7ixduXKOlZINtHbt/Aj/V3t31uO8WXx
Znmmm9TliYAGKwYNJvtVw+hlp1/wOsPC4fiUTCwBx5UFRZVbY4NzvM7uLDOdkjNV
CeHhz9AFmOXSF1+s6EvX3MrUOQtbt1TQQBpLc+Lil8nAAcLmaqARMz5yjzmG6+ir
nNGgRcQcHpE0Quw4tA1XWBVLZFxDNLx1xHgbNPU6rTNLgBm5AtgeVz594gBD6WdJ
IjnFrBpoAf7ywQY1811kp1ksie4gKFZhCDOB0VXiFplCwVzhhTObxyi0k4stKAdz
x4nIamU7u2qQIMtQ5luY8VD1KcuscyDr/ow536Fdr1JElsm8kEZSzji5fnQzJBw+
/XpdJ2vPbagcmA5U8To7XshkD9emLYmiSiR2UcAji5tWlvBqgQSnbePMtqLa9KEi
zj/j3zK+2hFWfDvArDqnT3kUm922IdURMSmFhu+K+rv0tO6XPbwZ45dnmLqGgWof
UahCxpREiSU/3wurT648RSVA6Yz4NXfZ/+oJe8AYIwPkagInsI0BcyKkFaMo5SmG
kwtQZdZdwaGp40v0L80zLsoKJLo+/iKEf/J5Kg9oUBrzh0a+OV+01cw9VuijlH/F
yACr/Gfwt9OdcU0U05uPAgYZwQetNkoCqwGMyG/P3Z+3otr3LX1ZO2h92CdGlfnI
7XTFD4Uj5uRyXsQgyiRkhxLZ6QULEYh1FoY+75wQbtnv3gSM6BU4cISU9CG4TWrK
60E8LIM7qFcpW3ksUuVqakpmWE6r2HG2LtX4k4xuz9TTlHabiO71tBBoXLQYOqfg
LE5SQztJF73CY0lgt7bqseGtIfFdX906Zbfu/yneLTyZqx4FzIcB5eK9Jq3mWyzs
5cvMgaqKZvEKXqNYTtlg4l1sq2UdGyDhBQZuclkZMqo5Dz4WrjYNZm/d5973JTKc
sqrs8XqyC9h7uAp0YU7Zv6ZVWvXWE6XZtjOiINfHSpAapHLi+4ymXdML2oRdn/W2
A1KrOE+2hC79jhWJNpI5THhgCU01wNopAGGfuxxbxAia3aAXem1VnCxz1CdOMCmW
ua6QhTrPzhsgivmQL3dofurgsvL1AI8SRE1T7qw80NV3InK1aLYV+xNkH6aWGUBA
E+h2yELvQaoxcXz9J94To+Qx+xCvXsG3LsTRoJB9hQ/Q/5IVBh5ipKJ+LxjGSk0Y
caSh+zw0I/sM08KRchXjGBVMxllSsQZrRHmG99UxwldM4VUnSajUlPxHra2bbX3n
Ru0gbcSOdyuKjAqM4LmuAVTPznluM5EuiQOpV1mBTc8C8kFPrdqyU2Vv6fDXTlC3
u0tIyCfYOfThmeXfNAc/Va7KPonAJRhVUTFpD227enw9i7JPHv3Glty8KnQ1BBkP
Qam+VVoxN5MX6oIZ+QHJhfRTFU13so4n9wLEsVKBQZr6UZXaLxaQtELvUXNvr/jU
DWzQ35Xd9GWVZoqOxo9MY4TikyamvmPeV3ciz9BlEJq7lghSIGB0e0ymEDtUNz4V
fxIwlkwTh2nBVZvIjBSK2LSHni6k7RF64AQPEKRnF3c/7/ex05wddLLBld3Ji61k
YA4o4K4O+IVUOpme4YoNYAtZPaqIpJd6uOMNPqSGQFhQYy1aRNPdVo2KVFE806vy
AZK/0y7SfiisFxlRSi3wMvJo4WyC6gPmwtPoiYza1D9JPuWePveQDLPbB2XsCXqA
UrriIWUids21kjoiHehPR47tH8UVfidKIu5B1+TVKT7jp7XB3n6Vz7Wxhqi/DMx5
kCQYN1AC7PWEq+8vcR/6dOlvUZ7z4rO+hxUaJSY+wHTGFGhSpHKHOewHzwaqrnpW
elsmOlYdSMAwIxU9IvIYBpiFQ+egxk9PzjPOwqS4rSVUS6wtb4GdU6Ij6un42CyO
3ivXd6Vl3T/5hdv6ICCynjnpdvNoxTBLThDDG/7GTHwhn1rvvR9871mjIncSKqTQ
s5UiQg0pxhHWZt8/wTl7tIbK96bNI4LB46x0HAigEWfV6BQfszUWfQMqycpUU5jk
O1MZq2wK0kZ+p7MUm5uLGUYPVTioKlTxJ3tV95zPYCfoe9jquFzrgoBxyN6bHP2E
GgYDR99K6YwYZ7orY4J8vUxrk/Rdq4csbgQ0uHgcH5Ow6UOmUHn7PKkREgVENYGG
+mv1DpJF/i7tGle3ke2X5rMh0YSoIOv+61x2a4EGut6bY4E4UzQ0/BQIwmc8LB1W
YNM81eKOEtpRlIWZ9lr/HHoddpjuHJ82nvc5SVu1kOdjqiejjPyHKhSk8HhQvCAJ
efMueT2lTXNWKg3mUQKNQw2fP/gSoT+6CKnAC8A8sPo58NdyZDh0HHfKATnvR9EP
knpdf7I/udtOslAx5aQXYnp5gkgcov8jNZyJRAf+UsnZd/uWzi8dM7e0UbonHQzw
94GIyoiWg0U0ccvIrHVEpUX/veT0wcKArvCAlhuyu/PyIDPFmo9Y5ms/+2ZdDED7
ooP0r8+ZU8gVRLPEJQefPmc7m6HgXD//md9TRk0fZktShwXgpJ/NA+jhqDgNQX1e
d064zT0OZvbOrT1Mo5WnoQAvljcrKX0UMy5525hef1ZZMG6ql4hBPMXgj3ZI0pSI
Weqndk+CHJPEDCsNUYbLrQyph2XBy9hwdQkV/0c+kBfbNNMlANjpVw3op/MGZSCc
FxmJIRGdPR/7kZzW8ooQOsK8TVsDyo6bDYNnEQQLuHoE1nnDoAao9iby/5EELxg3
A9ZUDGVFv4hI9L6mmupHMOnObSxacns+HNWOCHjbmAvTUOeTXZDFvfesPApfm638
N1gxjDm6pXynr19TsoL50JLNu9ZjJBG4cRy6GoWIPZVKoawRlpH7ERXaRX4t6HYg
ayBesxMCdYce6mQ013biTfrOmCyGpC1TBTJkPWP8VFUtLssLGu8pzTz5PvR3LqjG
0VQSnho48cXOgXX066GRook3puGyjZV1zr1ToUwjxBh92D3YE3pnScM9JIgN+aDG
6HX7CjMUh6Q+uhxxkqlANyt7r0zXiQGIeyb+4juFalR/x2lBLvrFRo9L7Xjm6Kjc
bre3kVtQKgIQPJxmAu0fMHXQJUqMJyPgXHzFKO4rdByr9hwhm4rAB+Xn5BkiKd99
MhNYExB5z8ZSvH4TSPehIZZKnOSaQ+t+gZOijPvkl8UYOoFtoaUOhFdNeTcjxjw3
1dWmrwi4mjY5e+kuKd0zfLf8ep3x8c99iPggNMrWJvWOo4q9fwuEbHhKKzAde1Sg
U0Qu2IaSZMOebJcoJmQM4lmPZa9tjZ+1iB9m+dlr6pfxpRPBDRUXi3Vg91sUbiRI
df5SfUb+OczzpREHPdUCmdqDnfF532L0zPTP1L2JsGJezphLFmFLdzFPbBmfmbrg
zu0k2SumNdn9F81qYVKyMJg6gyeGKR7L7EB0tgTYXESFnpZUDAn4DZasj+BAeTx6
5CMzxXs9h72SpYEVLroPjS4+CJPxu8bCZdd+LiS6C44hTmb8Q3i6su2Btz0ZCR8N
zD4crAjNhDk41lSOOQCdd1WKH+cubDlKS6mmIbab66HpEKhIdO4lWQ/dd2qKmfRB
xTuFZMOhSllfx4saz0CsIojBg4R3FtTYK8WlsM78o7NprEy7yieVv+Frmf2DtD9b
EYbABCNovmrDulknwRwRLCLqfJJiDW2Dszdljh/VyIBY/oap5q9vA+sppIiW/DTe
zZ1NXmr43xpZtVePXPkv0aByIphCMK6DCUcxFf6Y0lBRwxAuSlm8ATvj1OMbHbhf
rLH7vcsN4TrPiYEyneZLvP5QOo0YTY0h4uOe9p/qT82m9CK8lEnmvDs8uXl70qmr
QUAKZt6RkLCcHCf3DhCuY6SnVCa+BivWvQusdg+4+/F5SboCES8ravsqoeXvEwWh
UnsX6s7TLSLCjjqhY9XGM9mZLqFz8uEgb2gqbqoHU+j7FVi7v8oFcLRIB5BeUN8i
5rK1KypjTqTcSwMzWLsHOMth0CsatLIDfidRRk+IIUtGvKpSxZS0LIdd8+C8NbUW
Fwqo5Dn10SBsyN4rjaNG7QBtQX6IiIsq+v7OLW4dEqPhfsx5pJJdtdTEP8gqtXwZ
nywC7dGXzXE9QhHZZltm8We+I91OJBcIquDTEWT/kZymtp+57CTdptgACi0x1U4a
B7X7LTW9dlJOdzG9mVyEyTFLt7inGD3wuV4Ji6Y0COYLlvjI5wA1k84qBmDp0bPT
N/i+yfrrXVRpQ5E4ovHzv9FvnmPXabL4OCVAMNDoNGyUqV4qOTHFeopW/yJeOhSs
6TcnMS8WD3/JGO9nSniPqSNLUu/NI7nTRprdZ1A9lTABUqgiMt2qI5MTUEqbyI1v
EHGSDeCwUovSynkr1PFmxgamr2RCutynyY3Pv4sx1yRySt9FZJVe3fn+5oPZdEeH
q+1YAEwuZWSh0S5GBJXEHJ/wmRL/BzZZR6ZV83n8bNhUpbWJiBbGQdtFCtMQEGMb
n0CnsE5+0LXCTzLRI8qsBXCZAWNSdInjMLikOwIeXOdRGtBzw9Wf4rD3B2Xaw9AC
sjRIRpIuQY3BY3uv/WJBViFvEpLIymY2ghldJWfhTpJ7sj8vpD8uC0c7sqHkdiAD
4f1d79poSLjOQX702oT1nvJDoPluA2dW/pMcIP6as2O276yGJhHdgSaH3UXLRll9
rgA1nk7UjS9xgkej3hWLblVVGFMU10ywkqcT3E6EUkTnDE+3wDoNmWzRGdmC55v8
r40iuEfUIlXwlhRFI83Y4FDpDUFQT+GGbtXIRDvMO3xGmbouThZdz8xL7+dWqr6j
gysaj4kD0bUl81NHN8bGM+Rwktk5+byzVKYQ3qCsNwyuiAv4u+pHW7oa5u87mbyO
/WVGu+P+K/7wsVFzoH/vuomX6a366ryoJzs5/hdD9CTKMjiS+DaRYwm8DUVpsJ8M
yeIeyMappvODYJZIzfTCckLBsSrvY+x9MGL+ld1D/KLhknjRfllX80wsCwNk6uxx
K6w2U0Cr8FPmbsBoTDleOn/aQWC+G73UdwUWz80KiFAD8zrRXGc5TdQZ+AAjVVFe
T0vEcPIaCb07CVhWFqyERXXFSfHl5JGHjJeLh2kjPstcwfdk0QkjGrthguNb4Cj3
ka2ziM19pabuJ7plVQESFzIJPiZCn6K51wFOeKfNXCDmnK9YY6pjw6gu4ZKhulkJ
X632Gvfy5cJF38oDXzOvJRivgvnRP9/E7kgrVnPlInTpruAsucBg6QHrrBN1Sx2e
fdSEWiDA2TfBud+SPprSLcGrQ5EtklduKHOM/8qeKomd9oWe1U5wRFrh+FgSKirN
D00g11dMSioC976jxJw2W48o6HJiqcmadYecCPNyoWJUx1LtnJfSpsJFDigBz0wv
mE7M4buavDjHxCW3lJiPbPyd+bJGLzUaq7wmgrv1ea2ZXPOOS9WVR9wxziTxuoBh
OtwLct2mP8CuqLw+dg69thFIdgm2ZEfnL2ir83/mHhE3GX2mxc2H3cEwVu4Ow4ay
XidQ3Ev2R8EW9a3QCqYKEJNYDeBtpvkH5W/aQaF9uyfFCkjN9uYxEjXj4rLHvReH
N/y+cZkvi/NxLp2zDev+3qsiP2JtRL3nnYMbigISh/a081z+4yOXcn+gSNDF9M+Z
lfyW6tgtn5fveyQcGrvPtGnOl7gNYeAjo/CJ+8mQX5VAykVkCu6lc0kB8MTrfqhI
z6CmNXwtnDcfXYUGwCTnMuaLm/ZCGMwMZgijj8umJ3wggo6tVsmuTIb2krlIwrzH
HtjhIHz9okvOHrQogycj9MgUtMMBD+ooIo0c95PqVK/lLOBZRILSbRHZJCOPZYK1
SoXlcEiYiasHcJQP1WLcSH090TEiBwVrOKg7gx0hLoGSfokpcuGXMYpWz0QhLMqF
GfRVzRDV1ZUVQtp5nlmB7Fl/zsW+lzhxbbwSWQJZI3yCn3BjROC6QYc7MbstO6Xe
3Cxr30OkHz5Z+Hkwj6uTd0E13cRX+pF8pHX0sb226lll3yD8DMDpNbL2UHW8WECr
aOeUL59I749FCbF+826a/Yb1UPrXslvu4LrkFNV/M81GikfpS23B7HImuuGFkvCZ
6W9XOiDVadmtKyJ3QUNGeNkjpZL0svdKABpolp2GLXj/mKSUtpbpN5ol5oNLIj/L
UtF9uN/HAlo2HvdWhKRkpwdRRLeva/7OYPLmw8Uv9EbO75CWJTG8ZuXsT+Iz4Wzk
atYl1kbLDaEPTLjj/+vlLvACB88L87z0v6A0sJiWFcFJC/W+iT2eCV6RmUiibC53
LWd8CqhQGIytIjhFFvqQ5dmMzPlctdqI63sUdN0MvdZ5BzkhW5l5H+RhhC9yvUlt
1oksgsQhFJj0Cuqwg+f6sUi+f8X3vx0gs+CNKgBAcmz1VrLDN1KbVIn1Razy0/wk
tO1XIDRijO9NPmAGjB9zI7vGte2/d/YIMECLiqH8/aaFKZ6+BGJh6IqbFWOqgc4s
tOzJqjoQOf/QOkvbDt79Y2QaPI4TLGZJjMp2KiFf8WAervvTZrHQ8qASkJIFDFvj
mClmc2Fkw8RBLhnLWXsiOnyIMisJ8y7R/JExojsW3PFqab4I46RZY1UO9Qmj5h50
M3STreSmkQvB99zjYee17I8WGBKi+s9mn9t8zyBZ4FnL0bcdcEWMF/9n1pfRqr9/
KwJF1vefmeSnr5d3XNdAN0lS15BACh65kOw3Eg73VVmc31do6ex4g91980RLCb/j
R902Abv2V8Ujgmy3lGJ0BKHEjo6F+f0/an+W2hnu2XTHRqoaU88Mw3BP0adJpRPo
7tIumaDPMtEpz4Wc6YkV1g7ZBwdSthvtK5Lp0n9sjug9f/9ow4gLof2apPPBh4px
3MGwq0lcRogPOlQy9sO3VV41IcQhZJUJrfLTeHy8fNwHPOE/RXYWyRWrXr/9z0gk
7dBovO+OR9xhigkfztaYt2dHOPYt6T77sK2HIZAKCeoy5hAeaLjvfkD+Jh4kcvka
C6ckgJJ2wPEuRNlN0pIifUnjMCT+eJbfUZdagrxCfXc6AAASZyNk0L3dVt52JjkF
NkpMITqvhxnqVgcMKcJl1DzM6tjZnLyMNDDxCRZ7piL2JFHWf19C/vRYMB9dKIAT
TZQxpyMIXrwkjEHD+OryQ6ogacKhSjxdK1nK7p5sBDU/kNzTO/RfXhFyVXfzPvnB
Mc6UL//USUMiF5EX9T/hqEOWG06wDLDw5d9qQix8YCMN7ekl0618gd+tPFr4Hmw2
Q63P5D88xbbiizBz+SravXR+9v7eOi0KaSSMv7rwZEAIwjsmVwd4XEVflnREXsQa
D1fqPUFQ03//CfeyX/TsPwAZ1WPFAJit3UGl926FYG2t0cRvtrkwey5d5bnKbrgS
cxA7ktp8ZFlgi3Eb1WNatD+sxHV8YxmHTHGKaxC0EKr/4WyxJCBUvX/iH25SBKzx
LLDN5jg/rFo9sYP58fmV5Y52EvMLrd68KR3twDymE37Uq0aTB72Z1CIMhg+8xTeR
7NBqnSZyODSMU3nObJKRLX00IqjYtGQwx8R0dTtWcdbBwAAKtPm5itAF1eYh0Fq1
qOZI66Wqr8jMIphXnr4EmzlzDMmBoPqQfXW4IBIWbOre7dyuAeYtu1v9rPnwHV3V
QaGXVPkG1RDn3gfUH3A5twWimeNfzt9J7jsz49kRImNufbsxVGIkkMlZsRrGdrK+
7lrc31WF15k26pQS/eIPJgn/2LUWqR+18EqhobSVhKHknuZxcYbRIpROEbEciJXy
KfDs9ze/uoMQO/l41vLVEjqFIcwjZqF7y4EtggLVJD4CCHU8DZ4SSXfIvuT7jRDx
t5JBzovNSs5yxULgscEVo4GyQQ+d+cfpNYAT/N+lnamPJ3kx3dJ0foGOFF0i+r4R
gAqgynkkidBUJc0pELej3k6PYUWtnmq6o/eJS2Rgt9/NX5EbyWMEH65X5otBRXOo
FiWetCm6wqSFW4HZV9JuuU4vUbiH6Ot+uZSa9Vhivdf9uSYLEjplo0Ln3NCsdjk+
kOc5ugjRdBlO4A7s17qyd7UrjN9E09cUCIj/RSd+XN21sHN5uAxK970XhvjcOtma
fV6Sbbpg/TAsbAT+bfSk8QJ90F/ba7yQYK1edeAGCEbwYL0U80RbA14BCiiHr2Kr
XB6gj4i19fdE7aRDWpbJxrDMFxdf9ixc6x9MPmd/JRqb8QDdpJ4+s+RcytPyrk9p
ywQKuTPDsW8bSWqOiMghUf87Treg7jpt4j4OW7yw4U9/aJb91U8DFkuDz2DsuG7G
HbYGIP4U/yQpGFjlblUX4L9HsAP3G/YxNK2185/1b1SbEfcYktoBDX0NnV4OcaHl
IhjzKYCzHLqZqetPag3P0lsTDolGK1WX5nxNgWBBi9l0f2zTxJHqhXXVIEobmtaQ
3wNiPCR9oC6HCnQN4WSoYg1kp+1o54D1WChAzuzMnt0I02xmdKezuq4Ng9CcxXdE
HyPeWr3rTfLMv0O4KZty0xlzzsk1Z7GaQN1yQamMdh2DTNdXm81Mbn9aA2O/QSlL
L+8kmROz1wxnVjE6NtZd3LFAqWgFxkourOwz7+1Fg1eIoKf0BlpltudPe2wiBAiT
G3RyqLdJ9aDsNwZRKlTq9Krw1DKvbqQMSr5Jh+dJnUCPlURxftCq882vz3VZ4rcs
dbsVEXvBK0bmxGGvMBq4J8l7i5/unO3Bid4q/6MTfIkwitTeZjWi8jM3u7lknHkk
N8d4I7410AzUbTV2H4fTaNgcjEWGRH4pgCk7jbj+sahdMEY5IyZvAZ8BNo1fvXA2
MwJDJ2r85Hinjl0mG71l85PsO8M3C08wNETM2sARfI3vquxaez6qd0dRUzSSaZGm
lF5Q2tZrbXqJ1N9+lmZNx0CP7qKkql8Lz8VHg/sGkgN2+wMCDQCgRXcm2183sd1H
Zj0fNGRzZWCQfvRV+MNFDXoLRePjD1q6pM/ftnH9MKWUJoNxy8Fwr+n3yn/FdRQy
dtjAt+Wev+wo0RIZSxSzno6RHNGoJMyuNQtM/HVayc3tC6b1wwujwXvkF3ANaMSa
6woxbUfGo8d7pdhvMgHA+Nz2FphsIdIN6ho0FX7hM+fw2nxBcPz1V6yIXPTeYNmE
cmjp5Ax+c5SeDU/Fb2gdQuT0Wmi4xVOF2KhO8c3KkkifaBMY8gNTH2Nr6MWUZqkB
+W4e4FxdNIv8sY/kp6BJD3xqYNe1cXOs9LcVFDzCFKKYIVteCV5K8N8fzpPKrjyy
YtSDBPjNFsoyG9kX20W6NaSTvPbYVYHXfvEu51Qpu129NSJGRwS8FPFkIQU6K5yn
8DWhIgOX+MqO60cr3n993PAJHyQYiklr+C3/im1KLsmYsZ+Z8htcR17eGZZYC/XS
8kKrS2kFka8F6KGJGBjF+HCiEPfC7ZN1fJ5z3bIhE8JoTv+J85+9af3mxAsldLxG
F2/39IVbjlkjWcpDIhF1GHMrxmcODUEJgL9rBz4L1HexZhtnLeo1exKYzLHENyp1
FJsl3+vFxWbGdw7KYVjxrvUzP8+jUabuLlo3U7rdCb3yOMJrBeM81qRmBTUtIkoI
ykSHNvKeBpZBgOLv7A12g7YX1YbuY+2GmfRXk/Lw/esgFWNQn/nn9R99gxWI8Zia
JqQCn2UMiYREZ0u26JqAJl6GXmG0+Ngmxs0mOu/eYGzvhwQ9EzeJX0h70b1UwVZl
Fj2ofJird5svSiQCJy/NKfPTDbOJTw02R87eRqhpMxkclS00Iv9c9CMHPF5/bZVA
+ZQ1YQB4eo5hU82rRXhOviutk1D08zi2VAOH/JFxXfEUDTb+PttT8+F8K1ffQ482
GQ+Z2rMjg826yBGQzLAUQb340ivukvKPXI7MbBgbxk6QRTswMNbCyqReyFRXWdP3
P/Sx3/wCAx/x/mZrjvpAsF0bSLRawXUEtEHWKMzICIwCbpkhRw90CrnWEcGhr1S0
Wgy0oWZMBONIkz7Qh6hT9jjsWnKKc5H44CdLXhVATSnswjcOPnOjt84ALRFmzhzz
XierLf/LsiJmPqDeZ9VjdwFzWCMyfhKK73wC6XPrqkt6huPPr5rogo6oTgWjM5nG
/TBzsnMQel3StaZjE0M1N67LYVp//7Ig3ouSQbZvzG7eJfaSDSVJtzo9gjbh7g1r
VHq0JQBeXtYNKm1rpVNSs5EO5nSYyH3OZkzLZCA2lUdsA5oNrI3vdNPVdkmabQuT
Z4iWMwGAtMlH4sjQTxP8LzY/PYkdjZ1dVid5JJfd0ZAZbYm/vSGLDXXLpOV+XIP2
GfBl2Modrua3t1XF2WnZK+6oR+rD9unva0Nf34IHYFmPdeYAZTLjeBSWApCiCbO5
7kmrrol1/zh/z8ADoq75cDvr7Pg64TA0RJnjTTrV/u6MjqPKwIljyinQFTXEzFOa
1S1TK02FfU76hl02yBvoLKoBPU1ZVY2vmt3KA/prpOsXhaORoFjwwDTucDoCcdi7
kdp1+rhEFiglv6ndf6cLj9fE8fTwLRzxfG4y0691ncAj2iVxYKqk2cz9OeRJ8qh/
eSwchOHrz5WAhr1UyNEV7WAU7O7W9rWjlcXp+WknsS9RCWtkgJx93WltpGQ/5gvB
CI6UwzNp1aBOc9052nYpXuOzrs7WzhrigMbnOlTnsw8exmLeYLwlid8+84otz0Nt
UgywvA0XgxiMma4oTJZ9k8m7OO1ONedXncnzzW6Q0iBAAIvkQBrvi/6rpVuQUVaN
fh0fTRThbqkm0SRtkCcpNaHIfHZGnN0spjh/piRtXHx6yTrW8twimgPIVOGU+rDw
GWJEhmNagF6fV2W48wax4ggBvBw+XuizW9n6u6BGB3xCJx54uJk0+i8aUYXY8Cm7
DzAuk+d33wP7GcyAH0axl/r0+Luk2cX+0Q9s6pQuwAf9DVxuNBD3JR4shry3Wfgg
wsyYxl95oO0TIZrqPmANfMDrxqQdM8tMmkmBfnLvQV87uHWaCgTA9XiDztNNw4eR
AA+u2fM7CND+X2Qn/7wdgrA9VNTsETmYR3aaGDcK1m2oubwnLb01cW5+dfNqa1Fa
9f1RdAEmxB9HRmr/GM5S2pnyQ9Y3O8qXpsC4MYKgt+M1/XOFOWqyP4LLuq3PMWlC
hpd2AroJwRNk1EnqBUwKzrn0VFBwAaZkk6xAnRTKjJ3f50fVlluwUi4L8LndtKHn
XdJCMR2UXhCtRawdJaUQlVW8Q+Ehld0ow8lsjF+XQFFz2wwLcJN90lmVOSq4xgkP
ZiHw9H5krwCZa8TAp+nmk/wqSze6fahR7ZixiORJPdopj8AWNMXEB8OfxhTW0hSF
zbcHQCOWgrLRaXG1t9WwO0+odwnfhsOm5PowF5i2q1QzR/Y1o1T7kyf8xo6vTO25
XoJheFzVrxBxpj9xv3TqoU2Co6CuoqGAV4PxZyD1nueM3Zl0/SIYRoCmWL7xsOcz
UlnyrYKHVLaC2Tpc1jgGvn8FpKFi7XmB46zm/OVStAqV9KMgIazczN4kB3OIFQai
CFhanMcccw3T4KTLTQYIHXuJeRwxEKjPWjnM8fj3Kuy+jMdImq7X1XJkfXG3aasb
TKCmwTFANadm6hC8TVuPBWZFUWziL+WWGKBF1A3GxRd5JKpaFtwIlYn68X+SJUeu
CPIehqNc352qx3d+1y6kegsAdkW+s0PE9vB0M4vSvgykBnFd7dm1xogrzOJS+BWr
2VJ1D2kY1cMjJZezSekQU3UfavnpfJ06aRtbq3cONl25EyHy3sHhZURBzdrDdD+z
di9EvNeadEvTb2tmU/D8A1qTPnzLw6BiSDH5MpLzsKN0X6IAgil9GHhhswtJyISK
1bbzPM/pq87+LYJYTFrRcx0LD3SCXgxmpe0gLwVRjV4Wn3ioAmCS/ENFIYJXNntS
gCJi4cq4m5QJCct9sN2c67PI28S01pcOcBVHMXxbSqSuX7vRPF2MXhWqQnFEZ3dq
xWcUrqWptBn5uZawMb/CQ5q2YvmQY5IyVkQkrAXWNCfImfSJCR03uqtSnQBYcOSm
z5Kr41oGY2EKQbcquV/uDSOkqFj7ZJFJJHKaFA6FsLQW8bxqnojHKgPJ4o3+cQoc
g/8GEmN4clbi96uht4sm/UP2xwsyuV1fAL2gUsoVFAwcuoK5VByeZCWy73v2pl6I
0af36TmgVE0TaoayigauaV9KPXPgcTwz3Q0KKchwgR8h8yr9P+s7MMdM0rPOdl+z
gEloWJtUYA+/uap6TXtHmoRpYV/tXRUqKaAVi5ksCze87zh39TQA1s8ARIYrtJdf
miUKDNwQuUhBipT10S/3XOesE6XyZtBxISQddM59HfNkbikTslcQE09EubTgIpFT
JMsMx3p4/14SGvpUNXX7ZWd9p4h3/HoNvYd0/rV2ko/hekwsdJRJiEgpiMjL/eiC
/qhJKmDHcVQTIJw7eVP08zppoYiLWhBKUKJvmxEc2qCYj+qKxZrvDoUqHQFw9FDB
a8nnXG2yKJa4M873gxnlwrx47K002LHfUyd4iHYm+Hy5nxmihKoqpgAQIVtExUO/
JDHcLAvFQfuQBtGiwo+L1uPmQAzqpAr4P1Kz0c3MtkpFIZoGjT4gT/XUYnuArFZZ
Kk7Rs9asxP5KbO+gIU5kqp54WohBvJ/ppbuR+I21AIl8Bn3VG8BvsqUgpSVqqGKq
PF3OGis3avuahiZy8/saxAtbu+lruHmQxiQ20Fj4lNSbxqpUfFIby1RIU5fOdliG
fh76CStvhUJiDzYHuPGI3XCJvVusUt8FSwN/gmkfGnAHtsW+SoYyqBoGUj6CU/Iu
hd0L165x3ZP5kAs8Df2DS4EDSx7ScRUNTmqdNOz0B7RbUEbp0zuj5sDRBs4S1c/x
PAoDCQtAxtig8m+VLWiGalHucmT/sAPKNdMg69MHlITrUBPX2wZxQ83+03I/+/Ig
h8kAuu2Gc3dNEGYJXZO0Ngfr9hXJjbpwna+CPTyKY0WQlJt+upaVD4vXzAXG8YCO
5FYDr3AdPwuwvLngSys5jZlq5KyaZLV2VnZy0Ob3FsPvmms4eiYRve8MDoWJg1JC
1KodxrthHIStPY+6hDgeja9PPq+tLFU0RTNHh18rMATIVCr6OqrrmbXlx0dmfi56
6bIMOHK/FbEqKqDkkgtN84bwADT67mmlwKuSIEbdcnlXUEv0PRuOIiVcWwABSZm/
HBzA9JfxkqKyi1QOGQe0l6eXrGNEpAfdHpVfc1CKURNqvc6Hd9l7NeJSHnYXBJYe
iki4NIZue1xYqTi6ugYzq/zJ6v/G6ArfLySqbBQux5le03iS4cjCqNrYPzoOYufm
FWnzZmuxhXMjnF82MTFcv/0xBGOevOCiTLXo29/ZOq2fO6622EaPRo3MTIEUDOci
xRhx1ILuOD/ZFziAoKGLFI96dkGAR/6pugA2Yvj1QpPVL7LPPVaXB81c7kOZvZcG
DtpwKL5c8EAQtHVB93ukTLDHPYZ1sDYyMa0M54fiXXyYJnsONLv8sn94YD+iD33X
YXsHN3LbvnM0eQ8DW4/4Kcjvh9UFkUgbFhjr/yL4qlLxNT1vpMrz77QGHgdsxBtk
4pkoFk88GGwYriNLQEmorT4fcLH5rQpJb1jPwApuMGKZn6ZPjf2slRU4np5Mj/bU
OayAIjQCQemYkWJfeSe7hgIGg4DcGcHFvMT//LoISo8LiGNp64x/4uomqNxEvqlp
zoaQa3CNXNurArGoHz50e6+0TIhpnXjNDU902FNqopTw3RdRyHQE0Kxc2PDzBUY9
3fPxvTr7Ta71ut8GEtfN6gDaRl/SbCQu6rUDyX3h0Sl3koScLB1yEx2JGGGTMN4Z
YcvdzD7FWcIQDzTDrCo6CxgwHfra02Vj/hgaEoyAfdS5TMwzN3xtV0SQtiM5JYGo
zSWdblpuB07KnYatnNOlOxZcg55ufpau5ptWeuY1jFHcHUFTbYtE/2A2rRgU+yHY
i3W0PPr/f/ch9duhDiYzX642C16w8kkmJxvVHv65M0L8/inHjPt9x4NYZisgas1l
1ejbAyoajXjRP8SFv5aoTNQdf94fVcEdzTrkX2RY1xDgGKWKP9yVki1JG6Q9p2Nm
vS64rRcIupbHfbDVigOMYy9pZ3GOMgw8skqK5NhmcBLmIMTTXbCq1P06APzvKGSN
JvQyDg8+zflcmhJLzphnYW9QkQu7VIGiyGaD8p91tZd/tkdqp56JPdipRS9w1wIE
1CeuzhB3O9KE8r0xaY9LRb/i1b5JPMIqTT7Xjz74FmGuFQKrpzYoEMwid7E0BCMP
HgbOFzECRQCnsArSsxEI0EANqQvAtGHUrz84UVWLu0xL0SYqCZ+k26Ur4Si2NZqw
0xPhjG0MhqRRcpEW6k3750FA472HR3ERNy9j8pLsPh40MiLxPF+ww9FWVPZ/zu1W
/Qd3umkqhlESOtutwGWbIApUTgDoNm6B9ulbnnaHs4bl0mymStSF1+X+45jACv0s
V/7WvxrHW/e++EPxG9bqnmVCKGpQB5jzMxRySrFY9vHgVI9c05/rnzRThTk/vhez
NUjEru+8iORHXjal/j6kZefzlHySH3dFuZYouSym2b1q0VRmEO8uLDmxf9ixzCGp
79VFRNJH43hH0kR7ZfAB6hdjENQkhOStQnT1+ve8awQmBJlJz2ERZCwz451HxI6s
f1hd+0Ax2z9po4DqyRMSFJ9o13Ja00nlKDrSZEkljqo/OHLTViPCmoF4GxySfUaw
wi1aldkACaxc31cgBZSJNbqJTMDlojIdTcgQlDoy+QIq0AOkk2emZod47N9a1w6M
idhPSk35es+Zlp76AJtvnk5uLmPfkKXyQ+V9gw9lpKBAUMmRSMrpx4oKqS73p/9P
UVTE4a8ksBfJZIwLDae6MbyoX3zeTWaeMzRaNGnAn7hmLQr6JKnkSPfBsQMcTxxM
VoR5xqfpjdQODF2M2Cx85U75A6fmeAzEEOQx2b5RSdDfzG9IqWofDviEXfBwPTmn
h6sxy1gFpixyZz1Z0Ro8a9EemheGPoPz65qalkoxdGQdmTkMDuD8qijObD9INtb5
8g23GERGTNxlZ0kCxE8nrrXd401j81caA69vfnFtbYJXj61qFWOZQgoIR+cR6cVQ
imoBPRA3Q4pWSVmPAITjx+Y0nVSwb8Xy8E9epkgpvpMgoWUJ3en5mXVtLP2R7inC
vMc2aBeawWdsR+mvNNewqe4xoVLnzBSz9aswgtYc2COhbCG6pO+ug1yx+Ua1FrVp
O8Zix8MCPAYBrwJseeHY6bOeilDkwsUIYCkUaf9lGqEzVF6+cEXstq7X8cE1q/sH
iF2nj1d6OAsu7R9aoIKzSlg2w6DHRem5vCRzC4TX5JZun/5QR4Z31uePZfKnHqpw
mJ+7tkW5u7P0FtsXk/chVjwUqnS+jN8q1NCyauFL9t+NaqMLHHgdzA1WIFYKU7RG
1w80HRSuV+1iEI/Q1Y+T7r3tFtW5x7lz6VfFc3UO5ndAkJE5QVqVM+nYVh8KM9ep
Om716XNZmuF5oDwEd2ncOywNr1XXjPO+f9UbBqlwEZM6BsAg4FdgX9d718OXviGb
wwL46sDiybxDAddMlHCnnIfsd+hw//mKREzqll+Xp8XTy66gFQLMeRmJpq4mYcHD
X/WdfSCRiCu8sHWDJeCjftWNtXVQ5B/fRJv6tHD1jLlqHkly2m4gCcmXzCx6ZsOQ
y2LorGBPdfY6qzdPvs3SlBCswxBbIqv6ZWUF+SpLL0MQUcMR0K3bytW0vveM1X/T
ZxDPdV4AFOZ1sSMwgsKRagaH44agEJiC0sfg1pbZiCfEMe8TqZdT2HLNXvs6AEJQ
po5ae12+7w8uBoEuYcL5awhxR1MNmu/lX3yslV24jM/OtTSboQ3knrk/14COSVJG
80oW2op16O1i2WTWbntM+CirhpBJiLb2WbIJrR31bqTBYg7Ws+LZIMEkGBj/mc60
yP8xD9uEEE5OWNldXVzm1EW5hChZ8l3hc8BKxaW+IenypoNRKrloA3d7p89HGwjK
Zx8SkgymEp9JgIAmUL+YDnoTzwrZumPe6CR+pVs5ve0pfyMV0FRs51acEy3UP/H4
sGI6tcOKbKbScMjHhdpGk45biTzCFdGat8sK/mCNukhnaNnkCDx7pTN1QIgdo+WY
t1E/BVn50qawMr66ZeGI9GNai5E3QigMiOpnCQCPkxFr/Eh990uIlm5RhxURgUMB
YwyWGW229nZQSpKmbN2dTqQts/9pPatUZ2sXJLq4P1OqnP1lU4v4k/KtGSu6/riF
BydKNkq4kdIhOxS2ghRoJgMpoKlowSxd31yFd0M0S4pm/unNAbo+V1UFy0Fq1yPD
Zbq2w3ExZqptxw/LQSqVo0K8IFMjDxJt/b5nt9xbt9WscbpTtnuJ4xiu6O8umvYN
r/e3EIdJCN12uEnI53b5ivPiygP1DoRt/mjbMpaL+TWIJmzT6F/1Ct9pbecHq8Ni
KbkdsTWfe1X7qYvV1gZkFgcHFhUwAhVJ3sXKn8gBOUElRkk40+AIxhkSwn86BvaY
4H1kGf4kSipsZfxueV9rLADwE9JkWjOqGWpYYZPx4bh6ohhyBvi2jl12oR51vgO+
Gajc3RJgcupFh4zNy1dwkKv3ogNBAD8x37bP/wTj47h1B3UKkXlN5MTx9yjpRTTI
ekUV5w1SzvJQcu6DwF+VhigVsxzY4zM0ydCZwjgeMs/FicI36oResLKKZpVnhteI
PeuQjOohFntEPz8fQ8wJbRlZrORok1ViBwLON6c1qydUp+pbwmaxCpG08J/+bjr2
p40YDbvqlq7YLuh6uvhr4/TnH8beFCTjRK2zhOQqECz6VXhHYlnontE/fcF8B9ND
2/N87neG/igcJZxqSdZGKr3POWZmTR0wERhBpIN9TeU0dY41JYuY70nrUacrJQep
z/GU2xlGCTk+eNjoOy7Ph1kVNnoNV+NjWAnUrnt6CkVyUSFo747uAmSncvP9Cw+K
3dFXd5j0rN1jgCScEgAf8V5XT1hKy0h3dVPIi+WKfSeh0cbIfPAGE7QzQEM2VcUj
XsFcdcVmzgnplfCc2nrE5soFsrtEbkVyvrQQ7cI5Y/wz4LeELZ/tCdxsiK833tCs
pJtJ4Q2zlvXFr2mJM1kJpz4aWG7I4LUAZ1jiqbikR/pHlZaml9pOO4rB7eeJCCOR
IdUWqN9+z19r4vjkNvvp/LwKRBTJ/mLHCYMiCvNjhv1jX7crVnbGIiVdcANXKX5c
t8jf24VVkGrzfz60yjkiFCTwFRjgpcpL4keeVHT1V80irIQbBX+xWAxOf4h3mPba
SapmdUK+VO/TDSfm7jkM9nsZB3uA6fPhVxXs/92i4vxt2fjubicIr64D60lxf8l5
8Rr1Sk83CXgcWOMYthE0IKh3kA/mYhTxI0TaWBBa7mhxI5T+UgxPTkEJH9c4yQ35
QMy1MFRI4QDh/CSgtMPJ6gtE0wf7/cQpFt2RKgMNHh4t/LnnLAF0SkBfo+fCuIiN
dO2qv6532MiceB37Mh9U8FfaurjntzC9dpbChZ/tw8+agj8oaU9SEMdy//3mCfvL
qbALr+3oblsg7WGsjnu9mNunh19weKGAgex44iKlHfu5P1uqBx+jgzJjgxJZ18RQ
sELGaW40V5LzXzvft1AfflN53UrX01RoDvLBPrVfTkBXBNUX64nWQ7joDo5xwSHD
UNWhKH1ZrlOPhMgVbW4tqGRpTnrHhddq7TuJMHWmNL04MUQvO7nfPLFhLBC782w7
OA97RCF3iigSG4xoJlQBaKfvQGJYx5jwyVvAg3jX5Vz828YnIThdMPkXIC8U20x/
kZtXJQZYCb6d8EQrk/JYTjk8zg7kjEfsW6q5l9PKHve2sGZ8iouBPzjB6C96qwpd
1t6L2BiZiDskGU78y/QERn0/zFRcIK+kM+motGlgo4SP+yhDV0JkAMEWTbdsdWJf
ivvRekUmvn5nDSSs+dEIYQK7rNsR3xAMhf04GMTpypPV3Eu9Nhm/2mhNkNj7DY3P
GYG8arcMUh3ed+johqpU/IO5dUzgUw7YWbiD5XIZYUDIrDWZ9+56sC0tvyR5gzaA
SC9kHuUQGaenudMW3RMdy8Y7GWkbfx5D6mI6oNqAJtio14HG/fl7eBDQ5Cubqz4n
ZaEThtOHEYhaagAoFs3iO3echKDQmJwALI8hpIzcGXRzSO9KXtUcv3ItyKu58byI
oyrneFPc1BKDQKTCGK/kijvJ0ezxrSzZ7nyXwrKNJwx+1eKe9wYUL4B3Zz6QKS5y
OGj7KZQkE0FuF7IWfYTrEkqp/AYtn2DMFhbeJZXZlat6lnJ76RLBXiwWz9KVVKBJ
oh6KlT/wuFrJCOfgSExEEobUsi7wspN49Yr5xEgIM16ejwvFOwQfFuvPcUpRLZUU
havtuUGH9l+rbjRlcpq9ab5374dBtc9P5V1IHU2hpW2lkOPNzXnSak9vW5vfzXtB
Mw74pkU/IELK1zEyuau0V8o9vjeAAx1FBgwVupkh7ZQGc3XsQB0YKdDjRd8jgCFT
vUFSNW1gDp//ZlSBhuXUKBRtR3o4m/Oyw051xcd0BwWjwZjuD+3Hz2JGJBZ9awW/
uShQ1JeXbHj3ZXFRuux1i5oZC/G6ixGvoE34r2GghTV/coFPTGd2Lcpl4XmFPr3m
JNliE5hBLLYIV/ZWvvj0YhmsyEk9bmI2V5XQVlTviAOu82gDd5/y051DD9IAle+K
jFFSYJ2wKx4DFZt27149Nc2fbhny2s2L6pSmjO7lNuUf4SbVqubhQvYmUMPj0MXa
HRdDd2kGdoMmgNbDy0YGiuXFqmjoQwF3/MWLLsWJef3500kB9Kkl8OkrvXyvE+71
iDmiyL/2sI607Fs427plBHtvBY/6u8HdeffTAsMT5s9ZhhKeWFXuy9E46EFZQ8MU
QkPUNCI6+CCOioMHfL8Vkd9yb35D0KwaB48UPKSvkv63ljjOIKx/PHRQe22iyo1W
oL9/Yjc2rDHe87i1+SIPsBv7uw7iSvLi42hLeNmo933rubw7GMy19Oox/jY7OieE
iHJCysyokoQ1vYnqRosTH3S8vWXWnyItdsZ9hvNrH+kJRY627zTFlW8/h/4BhUCn
3PqB1AqZcMtwywTDkVICQLjJrYa13gQYyW+HtW0aEw+yX7GMcOX5B/r6D3g57veY
eA0lJjna/VBAYIaNeE8IBwfTl+3F0DRpVIpnRkR9UMz/gxwXywcPbp10YKCSd8t1
WwUgb0mp0ZJDMIyEkjgPk1MEMC0BgWmke/RJeSo44evJj4xzeIwG8PLOaBYPyD4E
Z5woviiJTuLZToUpSXSYGAZDpt5Sv1m738AJD3IDNa9hTekm0UyiS3IJABZZ3Mj/
BuNkTPsf2Tvb17ZfKWPJgimYHB2JePKcdV5f0Fa8qh/g+wySDflCHs8k9wW4S4uV
t6FBvV0k/+8FvqEqBkTgSzkXRlb1WgvmpXv9ogTmFyfg0si5h3Yjp9Usb+gK0sRx
tTlEchMD8UOGlabtjI5mTbherBRF4HBp5LO9T6v4NuUU8xsBtxJBTv06lKunbd7y
2kVZIHQEWknNkg+6OEva35++tZoMLraWxJObC7UVljTet8/su1SAT52HzfdjFhKr
9ESCv6ZbTBHmzFj46yj+eq9C2LBs4J46HFV2mGaRxdY9hsd2/2g6UlyN8758BIzS
aRrbgIGBihkIzeRXuL6ZuXG2rpxDKIwVTVwomtOuhPPY1p2i/YoH8Yr72rFV96xG
3jfPd8BebzBMfOW6Ny2m1pHL8jaTYO9wM0s4k0zenKriIao/EwlOvaNILwVtkMe2
gwcj41Bd2horfGOYWVi/M5qu7TI5k8XU7VfqcBxcpv14q0IW9tfPbddOLYGbKbCQ
669etEla5QoDPPSpZ77zNFxY6KYZgK7/htK2KT2DeV4kZBzfQM6UtvReFmpLual6
8VmTpcNIEVK7zW2PXk5aJmDKL83sgRGlMzMvtyIj0YeZbhx29gtjM/OG3oWNqiWX
bps2HFngSqRRPgZmdvQcwaHTWWm0aifq8RadiqE0abPY3gLv8tyvJ0I3xr9TOGkd
EIGWurR0ZNFcrHikK6YSQH1nkDak+4DuakId10pOUNDAKvDvTEkJRAHEMONWIGHC
uDN0DWCvQifL0dSIZQ1zwqOXfhjgwrUCY2zIDf0GkcEWF9dYAmTjVIaupm8UqnRW
bTFRpadWg2381+oMhCdF0Mch2s93HLehh9NVqW6NcGflw13YIGZBBvwRRz3N+8MY
U4pT3b55zWn6pE42z8hpm+iefklmJKrdaaGp0R4lK+CANs+GrRulA3BlGRZM8Ikl
u4J51n/8CTHFR2mZv0dqK6Wv0PWujj+Cgfw7b27H/GuY0QO/7kU97klzXP0DQiJk
7NG3aJ/YZNO9FKbfbt89MfXy/9YwRTS+DNDLyvKDrTRvbqJQeUlvoaN75tcQnskV
BKmD4qMFAKSmcgeDqmEt0ozIcMno5Nmw5dYq03m/MOw+K2jBX3pGkNktp66K4Ys+
O41reh7kuXRO9kOulv6gwMSu0b5hpMvYwZnJH/7aaLp7iyb7tkXCmIu9brkgQUH0
dP4+qWMejILrj0DhfPyZewnSJAIp6961EDvKdlDKXdirFf+9xbrcgLbWWbXwdUPT
QL9Sjb+4FYXDT6aT44UhQ82TEIyeY9rl2EQP0OP3ZdT+1RsIy8zVoJwpgxeeUFRT
p/TUJqHyI9FNAXzcgzb9ZugFJQjVU1Wdp4AGG/RDBEXoik67tNqMCUi0gtX1k6En
aHKqUPE0J2ovOaf+/dWCtyDvvOAoo8XznCbvCuCAgH6kHTN1v+/d4ZfxXOnZxyrl
hssQBpLhTlubyJZg1qRIk3mE8SjUl5jOpi6vuMSOkW8MK/8H6ejKFMSawo4sklbz
Ft/O/6m3a1sAAZ5ttF9G0DYqPyQVAH/GcsOT77SHlxdbm2YQx9Nbnm1z7Jy5DycZ
7QMHLDvaMny2jd/d7apX73KGjPP+aUE9knoMLJccDntUY9cIK6majdjPV/vFe7X+
vX1ujLgPDcc/rkXu35pnlfZwX8+ciRLWw2r+ETGgMytun30VgiLRE5/lFpto9G86
5Hi0Kh6EoBcVmAVyCUiAIZMYtK7/n0RCvxMt5lpXTNPkTkzzi0Xfghax3KiHK+wA
rTXJAoRDFbbxeysrEaz42MVTksRj607hAqPkbW/P+FwnJtBHWceLBmaBQO7EMuEf
uGrM8Yxe2rRxhH8wcirIZ0Ms/5j96nxFZbA+J27MojL/EsbmIdJ0fz54vIJXs+yf
otQeQx+SAoZ+/3KSW7j+Lwf0RvZCcmxIJ4d12sXplgbKD8dtCVtSQY3e4tB3/O9c
ZobGP3+xsPpIT2UDbSbxUZDPq3Xuxod71pR+ULF1vTIqlUNS3RQ7dxsvZ2WU+B/F
rJifw5w0k2QZkZPmzHu3KwHkhUUMMighBSS5V3KQsUjVlm64zn35UEro2lGADfKZ
YwlQ3vohRtkotRB3WDCCsPEM9vxue+1Nrdw8JBydqllR4TEgaz8K/B/Xp0wYybcq
000/p01MiLDs39JJ17w3Uz1CErevMLzYBuGMfSTsO3m/ksQnpVHSoTu44iMtc4CC
gLJJA5cZai/r3jRtBL/2CbysXigS+NZhHUAkebEvgbJh79CcQyayOWtzr5DhHPZF
/3Ye2l+RPkCXIaka4qjAb3YxVvnYrav4AsEpLz4Hg2GtX8iw0phcJ8WFfyiWMl1N
9gqUkOeIHF3c0cQwDxKKOgMGiFTYV2wgfq/pc9jDejU5gPjptXUr7t2tmNzXTN1v
f2P4wHuhGB9FSRkfOyonnEYApiyhHmYNEf0fPa1G/LkhtRc/zUvRnBUVxuul47dg
p2BF2GnavscO3hf4S/Rh3uwKu5u4pDbahfmRcJAqlj5HlIm2Q1BveUAVzToeGCNg
v7ydfsWPnbyOe6CuFhra2KJiIwSYBAWCFkuxrq5E+AqldDpCFYXK8vThdDJ1miCf
NY+4pqy6ZHV2gAYY3J9IES4mSX2VA1Sbe5tpRMKOuUrfF4dz2iCr+3QxTrRYDVOE
oKkevY+NzHlDheggMZhwmgdRMUBBgIP6D98oLhuyUzMd5dud1QGNRANgGfDWs8Gq
pfisdJUyNg1Y4qcuzve2qfjLrIykesl+DjBYHQCb8cMwe9NcRxVjPKPAdErT4f0b
G6j9pdYSvJXFLiz/AOXjsroRfjqv6+ugwFKXp1UK8Co5P+9FXbGVQZPaa2nV3lOG
0/pqOmohQT7cyCbxLJrFDE0wiZK7dElcmxDhl4YqLr8FTuAmRsf0KCGW949HiMm8
AY5Tm3b8884clw0rNTnuiUx6ppLDnx+Ly9XgbA7C8j2lzq0RB7wMAEvXcdxc1VlX
jXP0+1YPzLsdNAjIlyC2+tWoU0nK0GMnZB6PjpmTLBq/7pU9uNJd6HK0zZphjEsk
X3voYSCkDovXDYxOdwo52D3uRlJwhaqoXsqIup4WlIcgfrk87YHhcJu/ce5Q9zN2
0hVuHEe4a5FpBHjQWUPC9PzvLqRu5pTxQu70r3dwueJqqrj+8IBLroTN821s5u5o
Zwh69kG4oQFBlcTU+ONO1fT0uGyGS57Oh0GIhsZwDTPPJRPEKAZdmjDpcWbD2FFk
ZFtnp/Uy85bMp2RrxT1yiJzxCWqcoySGHNXtpuASD+rm+XQfuz3oyoJyL+AZyPJz
04WpEq6QExLjdZWwJQkUqw3PCyQt7wJKxlqaMnau/U7WGqRB/O563QIQGezkaGe4
4VEpNCsXl8K7y6kvyhFfVhbU8IcQEE7CSwZhmakYe+t1++Y+FXygbQg4L76TD/8o
l7RXBqxtEbs4MpzpwlUsYk012ZWBFBKOxWpSPJFNrY/HHUsI9oRGn9Dnu94qYUH/
wwFykERSj0sbp0FASBbmETwOSEuBW6pg3mHIbUrAuPHIuU8PvK8UVrmXSn0MiD1u
HV+b6xs7etD4uTWJplLJWi8LrmvdatDCLTclUig4yg770OMURT5s4M1sYsbyrgAY
dV3E6QdtSOBmEdd6LYFcxfG0Rzofk1bGfd87IYlPGhPivn1TRsIOWwHXkuclXhSd
5oUSe+8ypc/RZOTqRzCMyXuW0kyUQSW2tmuxwMv8cXwPpuK51Y1Uibdue8XSsfV9
vsJtPJ/Y/9GwUt8dLhoMqsi2tEpe4xrwA+wiCmiR6fED6ePWu+pUMqsvU9LjrcTX
8reFueeBtb4IDUgXeNSlnG1zY6AiBcfy9YkGPSIsTya2SwawDVaIz29Aut/kJcB0
QmwmRbuKZK6NGmrGsfhwqY9Ata6W+BrcMnEmRsMEY/D/pru+r1m21Su+RQ2JZmag
+KXazkboIo61MBNL2T79ZKzn0yVIai4UVNe/lUSZ0wGtibFo+MJY6tvwMKU9dzfO
kZU2Qn1kQXXtwJSVhIFMTf4YrugF7OPo7cgxWMt0DKMmDO8Ln+ZTNoZyKtHdKUAl
L2/vCsP+Puu5TjOK2OrURkjNqvVT667g37Wig1fibYtuslCLz457vmxHzjJgs1JB
/iwA5sx4ge8DH2z5+g2SIqbkOfX7nlH3FkH6DE1tgd9uQlODkrFPB3Oonky6C26r
QeXgjjf03eQaJl/nYQ2jgFsPCCBmm/HzUpDP3ohk+Gntai0ew45ZWD3K4J7phU4J
UjlroBU5qzAjAA17EqrKunZEJx2bshIdKPWzK8qr1CaeT0GknSjnXD20gTgFQnkj
dabACD1F30eLfrJZypADlIYnXjShk60tMPUHWFzUkGdKyd82StkPiDFxj6/B9Sde
Lh1SRiRSwOikDEgRT6dBsmq5DmNNUPzSvRefwIhUpCIaL6leB8kawHQkQyn1CQbI
+K9sed22S+U78w/Y614dhMOMTY9/KrdfChFEdOR+ts2s0u+4BEJ2/DrWasCqfPDP
M1B4NTTfMjnjOEuqgWIm4MKKTHMClvMc6Ia9a5ia1DoxuRvvAbknA6JD4omQ3xfz
G4BlV0WlCFK9/hSAgg62T+D78KYiaIRcv0pJNwj2njUYcDEKjcom8IyPXHr1E4X6
g//9VPZLdRSwr8GQTr7NZN6hDAacLi3m/GqscYY2GHvC5rgcHuLG1BTEYgf7JYPU
prOBoPNRnxSrFILZKic4M4YKsSK0oEblKIlEI6mK6LVP/ihTTQ6UvJ5sKiq6d1o7
2SwJwBzai1kjpREvaEWAE//q+PdG4LXBYDXdWk+epdP0HmjiQo6g3NmuQpCmDfB/
e5yGJAp3ENSeNlUTtVr2nuRdxYpp56LSbguuL/D8yrMaEktoZBFC6qHRWDDBj6Kr
ePIG8LvTVGXMeuFnASAHln7ExJ6rcvwr1MJgovOlxaBpVb8B3sCjo3nEvsKbIw0s
er2fIv2749A41vCUO+x9xAxjvZAAO9XnE+1jAYCy6QokJUub5LvWIAio0PoVwACE
TpUtKgXkU2Fqx9pNYUW3e5+GiiNt/DZFr/9Fa6RSwy27G8oUkwZfLRnMOLvqrstI
2RNcV6BCckHvxKQdk3wwIiJNimeuFb4ac/3I/gwidd92M27qasVshplKAQ9yLanv
RbJSCusBkYGhND5P2nD7/FMfB2HcQVLO5lEEev9OFwqH7EgmV1kKOD7MmjxP4VEE
RipY3QGmvYNbu5h8HUTHr3sF6qNFb6hkCur4wDBblY2AucZX7QdWpajem9OO5zIl
AyIJf2iULNYo0Ya5icjjA4Y8RyVH4Mlpi/hXyicgW8R07iMkEwUZhH5UUkz/Mp6H
0QQziJappmNlopB2uleT0Ub6j4rEUGcRMbwzD4/ww1LlTebKQJeYa8NI+XoOLLBt
IKM+tGcACttIPnPFIzIDJ0nMFkCkxxy9HOawrcAmQlafVEZmcnK0NFvHkYwAfakk
cSUlqRRjmbA2wOuX8SbWqLjXPRCDPwipmHr0K5ixrJXP5nSfWZUkzeryT+TPEhA+
A3eGAEDmPqEkjyYM8+Az03JU9JzD833SBDx9QwR4LVIFGdzHMR5OBulTtaP+haPa
Qvvxk9LSFY6BpcGYmga4KF4K8QIRwMU/jg+vak9NA6MdhJfhGB3s+TuOdkw8R67Q
op3qSuOkQDuLZkpKMNiwhtAq4NgRR6Qwh+KuemG0Vv+Ep7fT2ccX0HUjyw7Ta0ni
kQVICOXjA2IYJNqwFyIup8/8oTxR2inkewTVsXQYxYHnHHLvi3O1u48l2udvpG31
hGH/VN4qm8JW7x05aAylDRoqsECcIrOLh+XiJjrHdAZcLNuuP8a1svBFrDt2iVeh
fpAgH/lIDqbQLhbu0fQtvrqCA2Kd4Gq+FfWh1ElIlnxf8XH8f48YyvFLS+aLWB2E
FysFN9piIzrBRuTn/rnih8KpwWwQ+Up82tc6yolhLOyCyVjIvJI0pALMmqAsNJ5h
0P6lbeEWbPgEJb1yAAEYGKlDQqf5couzUkVUzGxkXjRkCy0o5qI93J+wb4RgQ/6b
1YSgBJcZ1vv99smJdPVgYUaPwH5iCTPlY4zj1Yohe2ZrJiMgCPbdmLLpyKqaVlv3
Lbm2GRHuLfydIAUX1qMIG6vY7P5/SCjldD12PvzapLgvRTnsaM9O12CBA1qeXWdY
w3g+0OTbdcY3tNZWMKTAzSEk2mDLEL3i5JKkgSNyIhdI7RvbemjmORTeMQ7+8kl4
b9B2hPOsuH9kni+9Xt4UOtN6Y/EEGa8giAGWQCzGw5aPPW6xkewOKYt0VaCAbmxw
1oYQDbVTBt/Ey+aRD3PIXGPsX1SSp3KBta80ehDLjBOrzXrBAO1p4ZkWRGfWmgZd
D88ZTqac6hBBbio0gmBPXzKuCQg7ckNGvhXWXSDdjqxm7/WAEjRzkffVHnfjVTVk
AV8fOCM/xymGQhyUovwytne/pc73i0tkIhpjBSdZaJpunhZlRSitT1nZeEGVrhjB
XuRFRZ6qmw0sAPrr7zfTzt+z0NGyWLZvALlKo2Uj3UyWs3KbHxHUJuJJ6ehOu1Sb
q8rfjEdobpjJqAguIq/pwpd8JevPoJ2DC14dmETHv5yBiY/GrU5vxchbb2QQ6eEf
SORneK1MbdCO1xPY7e65dfhutRcpvFLGrS7RQSa+Pdn9+PxXX5r9qr47/27fIPBL
YlRQ60LHt6ViBQMnwv9/fClIOvsYi1Db8dpacPEGMBkXHAbrEVwNw/frnz+QPVhp
Q1fXbkXOz6tzfVFK+SWH8EhrpI5qHTNYPOIVftcurZqQRUjq+u8VNkU4XlfzX6LR
14BWhJHOtbfUKk4Hdo7xEYJ1Cv/0McqrezKe+mbY2kN0NeB8sGFBK4aAR6zE/wkM
UfrwsFf+IoWI+QP9vgriAdS1QXQFJW2qulW7Byu9Gvlq5lT4k3A7WRWAo3h8Nq+I
r7//eSHiDGaf3RLaZUmT3KgyTyqrGa0DiygwIO+GaFZBIChfpMSc7dKwRO64+uMz
bBPTfcbIY4AGpLtisGMsUHOReWekCUvTtT2m05+rj6MBTRJOLORTajNDQUR2pI35
nEZ4EFDls0wz0rswQkbFe/+5sTWmK4qs9XwPh+IVJWKdu5SqrivsLyFt4DMug0ql
Lcqz7qVYZiWez9oXWOD8InhLnVnDKiA9ttjJ3aW0kiLM1Nm+By9hhjHdsv3bmur+
Wo/M5+AO6teRnuwQ8HZGKDFrSRaKNuVNRRwRl7dDlnP0DkLlRMxp6ZxsiO9n1itf
PKjQN7/VyC0jBY46ttT2TAb8HlkDTH0eKFbvKYvCliMdrQRgzsWnWBZ8tZ+faYu6
rKEfmNL/rco45MWNL+lZhZ4iPki3ZPqlXiux0YwYQaOS97WbOmr5WToP3eArB/C4
80K3k5B6tjrcUbbELSCXN4NM6n6WQgfRHqRRMP6rG31Jy1w1qVND3G6+zQSkAEod
xDB0OZtXJfvzCz2jAPJzzwKMqrZ45o8bTSyKW+0FVYw6Svi1PXXVy/CYWI0eQ0OG
ovgKU352Xqf8Voo8lI1kVgqV4K9DZrSVABwDvH5ZrP8/PZVFUqzI8uPXJlOHcLuM
SN1kH3kvOW87N9lnR9QJB57aFaRJ3FR8gI3Ot3ketnrSgmh56H75TLAOEqyz6db/
n1mlPjE7T31UBORWv2+zWQmlGrTwygVEU0h2Mhw9Qp9lxUxfJp+TD+ICbxr3G7RN
pH2hfJOQW1c1EiJUOndopkyQ9AJJ/xMbcrOlyQkRxO0z1zjFKRHzDEZer43JdJw9
/xH3FHUKmZDV2CdeQvB/PCPJQefwevYfgACElzH+besXQfAsntSHCiD/1spT9/hE
lwsZCQth9v7kxnjmmHWDkmgVAsEUsMjGIl/QIgsUfs+Glt0VCyn0IqCxaGMBN2Wn
4UpZcXJFLrcK3+m/QBrh/euZZ237avg/bN5mJGHLthPM2nzPMK88yETgcqJIwNAW
SUYgqqJAPQHzLdv8+jYyh4UYchmRNBXfanWB3bhcxBti38G6tjkjKAen4ojBWszJ
CGsh5BbVY9cdPDp7h6/fTJghqEVzuE48hjX9mgxsh4z0vF8I1KjtoRKmkcoEo/KM
yGUn1aFDfx2BSzUMLg1Ax7myFTLhB9hWmz1WaOZsKyQyZ843vdQDhGFOw8WJfHUH
menKuk94J28S2IEOdSnWTXbrCs15CZ3myFOb38iEfZr7PPpoj1wlEzda45dpcV+h
owM9yrcp1xgGDJtZMfTzsSg9fMaIAmq/dKed8wvBeoyCvG7B8SN6ddm3G5Xmdq3k
L4fDcC/lK5Yv1zP7LqfMMV9hpKBXGZPA/dW8FCCdYn6bRTjV51SBNEX4AIeOwRWQ
sWUIQO0823U4zJxitLnZrbBlIeifSmyF1lf2bAv+EfA/KCFs+WMHupxAG2mMZ674
qlPV0BRAimNYMf4MrJnnRGKq19GuKPBNB+yvxtNi33/YnO6c86aty48QLx3e3w7P
lY3YCeAEsABk+2RdN0DIhQPApsuG6Te2h7OrzyHH/1Ju/3/TJBPvkN1et+X2GJvV
OcMOCfONzyi01uXESCVZEaI9R2xmf6RLaXwUiYztoGmLmrrRH5uXEwcD5JnitLgj
txN5vYxzATxyq9m2NwHItue+Dj8i1Z+rKbiVht9uRio05tezmANJFEptPj+NeSAr
8cpi5AGAJjaturTzTp2LCQe+R2BRW3VCBWWNfqfZG/5VQ0fhkacmDn064mjkaAng
244hccAxF7oNcKUscX9ErRPRhanVEAzIFFfLMhKsFFXa5lcRq8KLStn9Qmf0Zc77
TQi12mu51eHoj99h9kbu9CwY7ewXzebi+NF0kpD0xOpr++RcE0E1CwTVj713JBYj
/NAjKi6LvhoK6/7NsoWrgGnqRp5cpjGjTj90Rc2dY5IE+ddOgpummhM4gJRyf9j3
ruzcRwNU66xEkAldsHNtYzHts62ILouCE/kg6h93VR1z1IdHsB1obB7TApCWZRFn
zf1z8raTO54WV5rk73mLhA583mVisK7aQ5F7r2qvrgdKDQytl/EdIaV7oLw6hMdy
QVzVn8VLzHq3IJsbZq7XMbXRfeyHiZJAo9Rn18OivR4+0uQGCd2H76kDvLiA5s3n
hpwyZohPUdn/MOlokFzQiyz5qcVpgNLb9v17oJXcPWGsTCpa+aYol5zsLD4aP3Dp
bQqBiev1D8k/uZTEEGXNDPxwTp5gxW1HSOzVFDrpfbqEI/PIj2BmjXV7ezjVlLYb
ywnS6crLx/NUrovNzeF+izrZjadmf6XTSAwjEZXjKDpbQAtEq3bPWIiIFjtRGfkx
wN91Y4cjhj0koHwL0agxOOuog1VFkB6FgbYFFuliX0hrjZYnqOkL2z7CFGAoVy8B
b0JbfVbcl3De8r0p6jNW1Lg5yTZH51q0eaArCUtXhuy5LbrAunAZeJYl4tJFWPK4
nbw20wp41FmSvFWE2YLJRi9RjQCQYKhfaCsklhoW6vzgqfeUGdDW4QERl2p1c1yV
Q6PdJVzXAg9J09N2O5WZnPlUt2le1jpVF6MuN6ZTo4m5mUFuiBSIEl8hPyt8tOIs
nOQOdBJSQ91EDI0Cr9NdA2EsnaY/icu61yDbCcfkivxTF3Sy0AsOVfz6ENZdmvks
PYwzzztaK9ESOzTEVkJo2+/XdwjkNRhq0+D/HXlSYDWDBP6r38tSWVj9M9He0qyQ
zw+jfSHFSD+7BI0DBW2yfqvg+sjs+MeSjLt6FsTysW1CkZ0l1Y2u0BDEJAQgvwKK
n/rz1ncsEQcAO2wYVDtC1aWKhvkSQJarlm/7sM2ZNDZlJPCj6vM5g7lkRw4vX0m2
b1LwAes/qbijxYAy4J8ZNKxXmtY/3MoQIKXciBqHwXMvHfmeO3EvHf4f3fJpyhcm
kdiRuO00VboJtGjSr8N4E680zg+KlISv/72pYR+0+lksecFRh9IpzTKZQMxxtENb
HLin26aRLer0hsPoF05s7ham3j3lfjh5i1jVGAwKWC+SeXrKDoydVfKuYWhPgl2R
2oR5iXN5JbXeDLCuaAeXv3NOQVrP0gwl10HfE0rerYRDWKVnZ6FneUIO9j7FJd4v
2mRAC+QCpSl+J6atp4sdiz1LdOtQJyunQEqyPKSoMPkktZnG+ih7Qn+rfkWULlcl
/ZRImDlIL6pqZr8bmwb4iQGvkeLmxxmbhR8+xc7s4rln3FaCHcEpXk7D94XYRHUe
go5xSOMQY+G6+0D+NK414kCRZBhset4+ReTtTWu+bwFW1V7y6Pbv6pXryrlGfOPh
1J/PHKid4BCuBHRRtmGtsMN5bqhkbHmFKeEvRaY/ajN4VLpW28nUxvqUv99gfuP3
jstYjXj9R9CwU8Nd6jp9dPY648ke/NjIkD6epsm/NaarJxd/XtIZdv1TzntSVpoC
76oFBtZmHF0RLR3tSrqR1imy082wj6VaJSWfBs5PHnaGO+birassEnbguF8chHzI
2uWk1VLYfXe3a9AMD3wSkjAsfs7GmIx8fKfsLMwZ6JrW8b8Kwu6ZFzb0XeX/miHM
fl/hWl9c2YfP5QCTGE2hFQCYqLlyBTSpBT5MQDdLSXYFPSPdvYUmpR5V8SvOaebq
rthGrWbUCGcyTGJ1VR5FGqKG4stKNqhvnc7PUIBkCMjNC4vHhHYFnZwtFwEO/cwz
zm0UGZ2NwH37lKE5FjPqRGynmd7ylXZLaGccrCWqJhMZO/a2clBzeJaJx4N1PMh+
ty8YaeBFsEMKyvL6NU7KFGKVNLWb8ZN6Fwk9SIaXO9tfG8xf/hz9C4P3PLdBrwvv
dQoeyewGUH9HIAfr+REkeagOw4cx7+57Xs0Fu+9SGP76d9mC0TjZT6PUwSkNv3Y8
YGkMYGhTHAdCjEG1H/XahF7j5rkPw/Ql51+Dk2fNalPh3l5BLAg1moumJdGdLFQF
LeGNMo98Zs4h7/Vfb402sdtTudfZsXFzeAg0F7XaKbHyquTByWhSCi6562+J//sp
YS6FfFb6wacCf0qZTWWBWwO5Wr55eAM4UWPOvONboB9FfEGooTPGHM5L9kMRR4FS
Dx3PxaXMQ7L5kS5ESbgNi6XTnuOGlSpc07h7hS6l7eO78kG9Y3LN+44V1MRCamLL
g9UchPpr5SSHydAxAfYhVYc3Zzx/OSMBK0YYQ/mNgOqpdWW6ihBsqIIL8JaZvAUF
9WIhR06nJAwhnKX3/UdS38K/miSRA4asaaNjqoknkx0QwuQsOnjCBl9nqyMSgSTU
dKka4Ht4Mg5WwReGjI+5tOtOoIri2IQEqa2NG7AwhKCUYLhwHbzUi+uveMT8Foxs
e049LlppWkCmoul3qI/RIPBYKV1KOWCdc/IGJ5MO4xd/9oJtLcPKQCAAPyMQPQv1
/uf+tL2fVwZP3u27pQ+WAyvc0qkF/CJVfYATsmmEAkbYX38Cv2iKAHGpNKbsNHuU
cion8d8O6ckY7lHFXHJcaMOZyFTt9IRH/3s/P6aDBpb2EHjo1o40+rIrNvjPgWl4
dtK3046BDw6h7Stqvy/lkevYqarLReimgSxYLF6veT/ZSWeOE/oP7uI4zDohJYvM
zQZYQuFzhZbK7Tlz4C1ZoU706oYC9QhNebrUgg1KUg3cuq7JP8npHra9zkrKCa5v
5FdADIbPyeR5BXdvVxkMgBwjM10hh4zaAMkmAVzU9yZOJY4UwPlANW9+3s+Pil+7
ylB5r0LsQuGK4LEtCkqYJt917ILbSB/iCaezZRMiYxzx0uJdj+TRKnKH92ecQxNk
1AeHKH3GQgUOC7ekZDKAwAUwNFZxdlmZbSpWIoq2+3GUzN87/1IdyR/Ap54UalWn
CpmFdUQeUOMSDQ0MzRwOdVlFdzcZ/8BazDZfoLevwMMtYbjxm4fJVx8ssv93k0CI
VdrRSOC2EqrFAUsPKkffQJftnra6mLy8SNSXEshMiqU8fXBJnEKCmZK+6XD9L28t
6gQP4IRm75Z2rq5vASMLX2pdpbFYbl7E3jwGVsXKTb80t/tHwLnYHCKkCwmUS5St
HSSxuObvQOR6rIcVGrMc80x3khEi/PbgQf+stQEvUTTwanuzqMEUebJsO9f4BV/F
yaEWmApz4mmRPR8NXs2yLBmGpZit71GlI7fc5CE3LjvG+9d9Tc5Jd9RcbP/KPIE0
yVsFvFVWhKgBtETI/2bgIkxdsPyNOf3L/+0RgapoL+fli8dVytRkPCHlENLDklHl
QOtlq2I+1U1uQ5nyI6OdSpsgnjqYaI/8EUwmGd0CiN/8hb7g6LPtoHaDDm4DhSKp
q5kVxL0ZkrHPCEyilLxxvQrj/ME89sdPrUrm7QIqiIW23Py2NQmaKr57I7LOqMtB
WMPFU052Fqy+gRGnN1GhdI0a+EfE6W0rrLrisx0wkzg0lHvIS++dpGlPj04cb9OE
cz2KZSUa1p7FjKYmTVcF9QiluFcvmIlat0hiCWIaLmCoG0YkpCUvdCfWqNfH+2+c
5tgPpStGmDlb2ow/3ZCGDMSZJnBB2cc0S0Tx0Sybwxk00v6Inm9iUsfB1QrHkqfU
BtuPQwRl8xqJKYV/HvTMhEW0V6ZQGhUUl+wH1l8cun6V13dFtV7vRPKLqYm4QR92
T32LwCkbncLYm/WDpgCXGVcEBJqidYfT6FNKre11/6NrFopm/ar5q3hnOxdN8UXV
NU6HpOngGnEH5NORjJBITYokl6VP1tIGdVNYeY23NlwVpR0RTJfOGFEEN4SSlG8n
nXT6bTiCDBT7+VoXgFxfr0kS6bItTHyB6aF9imR3pafyIIJogmoJ0VR9lJ4adz7L
8zEhaBaJ2TIHWcEAHG49ZQLEenI+xt1YQZAgdpEqwmYryo4Pav8GKmN/fEGwqEe/
2LDzBE2AIpPDVaNEZ9vARvWgrGmK/i9k9j/yDvnESOjyhhUmfp9XnBe/AhxgT8K/
uSeuW47UXlDN45ifID6KfxIdtGMD07+0JXUkD/3Ad+17chVd+vp23U0ZRj7vK5Yi
KzMtpATPGnV+/gD1WyF56k/M1GDoUuYBfk3N8TTXEVEbR2xRYIAsSbetuqa/KlHU
V1qWCw5dsKNu0r3pSd25BnX+T13q1nOTWiZNcUGTx3MfF5Z10CAP6NIDMpvLewS5
8FOkvlaS2cjz1BQZHDx1BlqGM7b9LzztxYi/Uk/bCNO2VsELEYZFi1WyMQ6bmWZ1
r4iL5zh91oQUn6Af+XKYjy7ghYd5Y/fyZY2m26O4XJQcxqiUZSkpk6AEhyK3DjtY
21aQj/iWgH+CoueaAwx1KVt7dL1/55KKtODR1WeGXbyKKyxsm7mN2epDfMiPZnNx
dmw2pWUiY8Si+/16/3UuRU8xVdRBt626zs3rGnTJiaBPM922oZB9J7TxtMVrYMkK
DkTbG3zoIaueWlse0KS3EdiPeOLxCGvVi6riJAqenu6xc7O1DbMSM1A1HXixHhyL
gLAaAWotFAOFUdh9kuiidkbf9I9iAgl8K3O88xjBMZF8gabOLEmoB1KT+1Ffoy/g
etjrNPzjE//WSgpRz+PsTlt/DF5HM/wlFsMX5bnWtxcLmwqWcCtivg8PFZTT837H
2+a4fGKDBk7CyIkOix9AZE48/u+aawc9GMc3AnORDOLo9LVEvhZHSQWtAvJhl3gK
udC7gGEv0Zd+Aiv6/wwn2mUYWRY13eMxG+aXnKzifMZ8oiTveLwV03ExEmZmhtBg
T7HYrx7JGTrCmwkF8p8t2wiegXU/U7MF60Iryg7gU5DgeziVJpx6rGAhYsQYqcqN
USICqaqfbOc2DvGyxPSVV/c3R3/Qck/VRaipTAHQnr8O6VEpe7EiHTkyThsg8k8x
jKjaWcYwEpBEO9jMA0adxX9m+f6dIQNMKgdpkq5jd5/mzKEPkGfxig/u/ib0oM+J
mG+fqN6LEkExy/OrCCq5cWPlXucMVuoPOSR2W2qhAt7HBnykyLbtZuEwu+UBTyHN
eMXgXe9Lcx3t2ssAvrfDbbC5N7w425LslDu5tcpW+NvfO3VFSCfBOE8JROKNLiBi
LLHutijpprmmJZfsdrbc72wggnAR8dFeLwG2IEWJn1s2qhG8u6r2VyuV8i56Yf5M
w5/IjQHAHseSW1h5/CZcI+XdvhJf7T6QghBu2V+nJkorqsaxkaaozeRP3cQinOcI
TX2Udjf1n9nJ/seXOR3CJnltZNkzGylPRUqunyVYADBcyio6o0wViIcbBf3JHOlb
fJqjlfRoDRtB0+pT+NZ8Mq+Og1KrvHKaD28j4XPXXkJBiA6YElpKKzXAn1xNX0c/
jtM8qy+xKtoSir4kDVwFUoGCOyoIbZkq05c1/f0JllrC3gvOWNAOAzZgLQ+Jvi36
u/i8dh0uo2e+4PAiaDNWSFh6vU11aJE4B8lomdATNFudw+gLdlmoXgrLCYSKx6Y+
ap96neKvE9driQXn/SZImK5MA3RZQuwMHK35F80T1xls7LGsKMHluXBDLrB3sK3g
ArQjW+MUbqfkOGB13dlfIdC1gEk7s7tExhkkxdtHFPIyyARmGHIaCPPU8ahpAz3k
kG+6bgMGPwjwfFoMDdSLCr3c7k89o/3+GRgI+gVXJwSBaQCcdU0uB8H7UCjn2WUL
3NOzSzlawHdnwIXt6sGlUI0kedHlMWeTYX/kQz5H5Ri2x8zetrlvNYBs2Z0gVjdt
fBZarr4uHNyM3wv1wsqGWLtTl6obqgvZhKsEM8g1ZTT40hFl58dfXQNJLgXfU/DR
sYPUVM2yxc8tXX7mUnVQopTIphF6u0o8RBy7LGoWFvafcPMqeHbE1ccKw1/n22q2
G4wCEtOKQhQnrdMzQktZMADhufV7H+aCnj1vZIuCMZmvWARkX1W5hZ1Ert6un1VA
t8niBaVaft2/RLJOit+dIRJ0a+NlZcRPbKPtGj+ry6LPdRD7PJKGNrR2AQsVMvzo
8JmDnErcow0YR7meutjO6Ux0qmAXpujpd9jHqUXWGNRkBk5AzCyUmwMygM1/kH15
3xApI2rrMqPRzoTv+bolkRLPEnGdCxbkqpf8TCM4MHXUGR52FbwSkVK9LSszMQxH
FuInRhCsrK9L6z+H6aJUxXaM+QFtFwS12Dxg9Tr0ke4qMB6BhB2YofOBKsYYlcJR
0x53X7nAt3AVmBNEzC6MZ3j9+66pjABz6F1JYACH5SK4/BSkzDIpk5nZrCnyhR9E
EqpyC2tFUxa377VW1X+hfJ1kYswnjTTEanWV19/0yUM/m74gBcFC7+7qJSGDQieT
gGxi+Uk9kROEbJATcZm4ZIJqVnZQz1mSqYl+JvyIDXWaGfR4XEOSZzlPu9MLnlk6
RKdgPaUbkAM5Gc+GxNCxOEzz1sw+xC7rfIMMlat4sCO1oBVZG7IWs6xH6+q7+6cQ
/qiifxr93rjzMXwshZDEpg1dqymIPRBjaGKGq5UsFus9xKcm4jP3KI7Sxu1XO6yt
LkN9UgYcc4CE0QqBBSvqn15u4y277m9us5SKi74wg0Ie9eCbOdki6mTAoer8d/w7
RKL6NXbf/WcpRw2ZB06LVAK16uHhNwRGphWMVjdnIIft2Gz7DUv/odn/FlQ/4qk/
JSbI/xVh2JtBhujOIHtLJLBxXT+tWC07shXlth0AeYDLxAPZKWcIxO7YeVKNw5hL
PFQNBT/HCWkf0PtqoaRbg5L8hEAGmgWH5PyHoM8KhtBN1pOx7asC/Gelx/QPMttt
uAFyMkQkFXXF85EboOHYYZ2lMjbPJ47Za0xRpOSUA1A+c/WRE+eSZsn16MIHleLr
1Kyagol9e9RAPUrpdUaPi4dYPiPTa9U0mukv95ba0F8ppDrHqst/ZM0qtBSU7o+s
T3S9s7Nk1Bap53Sp34XydpxBZy1635a7hToPP2Nx+F2+RUyqKWe7gysj3cE/KVTH
SAL4eKK7mBpHHgy7SRgcAnFLAsfxX3nrNJ42G0fRQZnBKLwa6l/EWvC8r5BuxQOR
rDEg4EiQlsxfHHD9BzMTgxdKKEdMu0zovAC5aOzyphqIKqwGa+hkggAG7FcmpTbn
Z2STqtGwh1DPR4Ym6pYicAhVCNmBxt1p6fwkgAmIm8i/Lz+1zPfWRFHPA+IOqihI
8fVPeBURixdblRWOlivhBnz0kSHKEQK74arJ457Pb+9DVbPeqe6K6sXullAULY29
VhXmkWUPJ3qjYJpoXMwbtAOK3nHAzz0mAp66EySIG6P4vXV6UIIQtAl0shCDN7Hr
grGiqhkEKSrIW1/yMxujI1YpQIWN4mzjkurwHbAX0A6kcf010n/IqlEyO4OqPebX
n2WYfCRjnrzRGSJIHYVPJRtMnFGKyTqnF37a/z2EldZ6x+992OxEOjiw9G6jzglz
yPnWH1DU3/q+GSkXT4tn5VghToEXgNL5xV6DYdQ9EQk5hDk2MGIjLeJD+Nf/Atv7
lPk9yRICEAQKf+E+jryMOeQSTlcRom/4lCmIyqyed+S9NdCautkJj7OhT+pKgQ65
T/EL25P0frkztWleyUzyhm3gPvWWv79TdwQc1Iuhyic1TnwErbYsQsqKtcpskgUr
BKbFN2IDkPwq1ESuZFL33tzl/RuVBS84sgLxcL9w1J1kHaU6UxVmCZ4zC1CItdvi
8C6UDPeSyr2cJGuInTRzxpgeq7NLrVzras/tVxkJPlzrGVALsYp/D6LlphXI5eux
VB/N6ugTZ8rStFgrci3pz/mJ93kobaaxf8DHVKwH7KQikvDqXbNyJTk1cYjZ2KHQ
BJJSZJFbuCHxV6EDPkJvPNXcNe6aXRc694LUy2KAkP11GlqCOkSosVwOKbIc3pcU
Z/kQmt5/oBEBQlrc21Quy/z8978PgZyRSUdV1858wEZUN/WoPjCTP3gtkAZdX4qP
ESYnZq582LWiQHC8kgmZkHGFToz/gD4SWbnBrBNwqPGCj33X0LJ88ex0SKn53vpg
p6PivgT3+GnCu3ddsqAHxLJH1MHpt85oULIUfl+cF80qw6ykd+ukAxMUbouRhRPj
hmDyoCVW9EgOzGQwAaFE8RzNRFZxm7BkSpypC2ljgvKsZmBkRIs0BSV6i/NBItBw
WrT30lbDLC8TcVJkAvKzNDATbEzfmSUSn1NmAYvQkUAnb+qLuHqMA6RJYuWb1m7o
vb8UhMbBEjzP8go8iL4+KehI9Dp3Yc/ysGudPF/tvd7K6hMavgKBqe8QmveGGKvY
f+ZWCLFlF1nP8Vmu748WQreDaQkioNiPD2wtjJpAhhmJRxh2Sttlle9pr72SgWxm
Nw+sW7WvlOJGrIwcyAK9s6lq384v0N0DqBuF2O3cNvRdxQiOvv8uN+Mq8wUB4EwK
tW8V/NI37qjJYn6uROKUmvPPSzFZcsW+k9NC0e4Il7gKvlwrU7WFf8d4c8lMkMbF
VwO73Ul+vTHEZEJVuCU+uBdRKz14/ggvv6h/DU369CylRSMmsxG7JbJI6SAEN58K
5DcbbAeXsBpz/JhXqIDZhlmyGxwUmop9vTmFr//w34mkHkcvKzCNe15W7g07CVcs
FvMTBiKwDy7o8v3CywwKXf4Zmt7xUTQtH+MF8uiM5o6iBcGXUAxJ55VieeFhZ+B+
n8v4fBASYrfFzrixbgh/NVOpMNZLS9DniUUEy9h38ZzcdrrZ/aF5DZQ3DVx0DWdF
TSRBW045c73t+0fC24r/adTNwBdxmkihDtiHm/ImwgyLiCfydJWt4GDwYaApyVlS
0TaexRGaIlbLnExLpAavwq9VLYIckCp4z85+qy77dLTRhAp27AZLPaYWdwrEwW2P
VSCSrLTFOMOPIa6ylHo38cUXXE2F/6oCFOtaS76O3BMoF1qDQ/Z+tL32hZLDmR8o
n5WuQfi6Pgoh77Y4i/ramMc1wSDkc+6mYJNXjO7TYym7OIbb98uYYIlJcRZdEbAg
dJPGe7QaU+npQEcaQDqYVvbS/uV3i/1XzjOwC2Vxx2mxW3Lk6NnOX5fiD0JCyKFZ
xS7HaE1ShhGruSyMMBAkGwLv/+jGEHB0vaBQXCm24A1cN9nnqOmpjirJQFkwLkxH
ywhhKnA3KSvxfkinbFsQ2Usf8MGM91Ym9nySokLwFP9zngTnXJHJRZiURZZbSsd8
fHUQUfAGK1nyK+52xe1BsgyAXH+rr8GGXaS9yGfTFe/dbjwPKs8L2iwUYVNL4Mtc
EjirtTOtofAEwwztxSThM9gx68HZiyh1ZRifNupAAqU7ZSvuQj1JVfwBJflnPXAA
EPNeq68r8/FHKbJzimJ5CARkaleTV8RnDPwH3F1B4rfsMiFrk/bFJCRcTFG+/tfD
S8ckEFJA33y43DZBHWyi62TmlXmDhMV+9Pl6mcfzYaIuiIVwXXhZdV0lJo0CtONr
kgLHmTybCP9sLLVtBaUjy9RK/hubVHTsMZAlfFC9mCN8mrj02hcQaYI+j/9cgV2Y
V67OchKjCp6KODgu7glOFDg30WBUgzisCs0e6Aoo+eMTNLiuqxaF075vlQndIj2B
b3UwsiH5EmhXZVLPxJtZixfP5ORhfBQGRMgQCq67qdEgbkaWhVE/1hLVLzcX8sw4
6vpSB9tELH5iz1fEtxE7MDOITKuDs2vEzFqHjvj76vo38t4wpuf/EWa9ZgZxCPg5
AwJCWGAUOGcMMu8qEg3CS22rLx6vRMUTZCvrgjmvHTxJxtoN3iHnxbynKWet35q2
93CcnwPDapKMmu1w6Y1DNfTgeJDh+E0MI1UvtXjyXnevrkmQO+L114Rz+0NHsiwR
piKUmUZEkhDLMDpdOsZazMUl0QiFDeMplREX9WWE7MxD9uXOwbFIb33HWQwKiEdM
CYqUouIWW4W4SF4wmHBAl7Lp3FNjl9vGx3DnnJn8BcORMtSw1pcmCQAnhGAvURKD
sMUnyOyvMXGBHEDhgt1JbRglBNDfiOxfC4qYLiFeZRGacoiJsdxH81Ze7wgt/IGW
6PYljYozukjZEkHXd643Iq1oKLatqlkJyyrEXVwWjq3IPCnz5W/nXdkfGc1qZDvs
8xbbYhlaDxw1hedYCQuqNJ1iPr7+ROXgSkmsDGzvrBIOYG0/rhV0aIn1fbN17W77
pD6FVzc79L1D01GJfFQl0UXVxCHvVB0uhU2qLGmzgB0QMRun7Rn5WY+z9mqi3BLp
bymV6sij+EatHnZnOJuwZaepdG0E7AI1rwbzHQeIDP+NxWx/+S7d67zw8MDd4CYx
BnBNJHvP5RxsxKz7tey83GPe4TnSg7Fw1tzAuehXPk0/KwyoegNkGTn7hm9qR0/L
BRC2tJgDi5xJM1EFTM/UXAFl7a8aMs+qe1wvdOdMqwb5u6afXqWeE2TfCGW9pFjk
IUn9NLzh47T5gL/Ns9vFcyiMsLT1EtFymNf6GLhg/HgCzB+upVefOCimHyLKOnXe
Su5fpkd/G9oNCZU6wMgKD2FgjpPW0TBOvpi2L43FCrPG9N4weaxIj/jL7Fl1F/2G
hLHDQt96wI5d/2y2eONI/hooo9L5LXVOWkbz0h+TxP+Vg+e+hNGcifOwhMgNjv1p
khlkjz+PoDtrJCcvBEQUJWe+AZhNj3XhU2KPhHv8o3tVaen09BsQYYZQRk7JyLOj
TrzUrNzOmO0DtsgzCWmFCmL2wQY41rJds+B16MGB79jQP3x5fLQt8M+hi7wM5XfZ
t4Ow9SHrM1ys9yWaw+6aWXzUb+hSowLdiExMWP4XXYlh5VaH8sXnQerxxsNSAmU2
DMpXv6xAVsAL3jsDCBnh2RDXWgaJ+zngUwys1hEd6OTH5eU7CPgAHQyVQ62Nu2mg
oLQbMlfp/e5zWd/9UqJz9mkPIZ/8WAdFk53p3LQm/ClHKXK9CrpGZyStSOQUqWN7
gOv6B6vSLPADaQb4gdL5e3IJHJu1GEWmSoE7hlBmQKyzQBUXfpCydaW6xi1oapOy
OYhzSKlJQVp72Ir9uIaM/0q1J56HYSOttP4SkddYwRYRU6JMVS3pSC3YXkAlh2v4
ConYMin/lLuMfgsKO4PwKJXPvpg6HoF70zbkTIPLzt4P7E7TzXZTW2rKiEdbqR7J
1xhau2RE+GKmHYbN/ew9oOuTbRRX7lgQumoJPGona7cSrL5rdNpDOKIyHU25CUei
sjW/QCaOpKjrcQON1gAOibvOUoHoVmteehCVHK3x8kuean+OHPqACAGjFKZIf4pf
2x2oCv7ZXrd47uokKKLZNEBmmCro98apE8Rmia9DllBMAnvjlkHF2oNL87MW2E0Z
UaGrcgUt9813Cvp3dlrg4SWpx6+lLAgyWO8WHYz9BcObkVE4g4p4SItxDdSion7b
DBZVQVRWsiJBjsgbh42efMpGvp/QGosJ3VyBZtgVQqUrNLAqX8tXTHGkzAlxpYaV
HRcswSGlNq3ZvcxGosbjo0y5vIWOeVl1AK+97fbp2+DSL8plSI8tnFvGwIGssUFw
s7a1ad68bQ/h0tQ4YVen3c1+s5vOd1Pgnge7DlI4mk+G6qnVzLSjyY+1a8cYtxd7
xH0QiH26/ATpVqqP2eO0+hXktjTx6Gkx/uDe7C+w7UEC3JJ7bOc0T0y1EwtgyFPa
NDoLzNFH53Ut6KELBd94RPhUDz0BYI9XQZ33MnG5ubT+a/6NgFnvq304yAr/Mkga
lusn3iAnF4AVFd8b/9rP3IgIDsYy5K2r0/S36BmD2Lf+5+eD7oA+p8QHOTODzZYb
o1qw2tbnsdEf/MCotx1/JuSWmAtxbNQ56aIZOBXf6gN0pmKqzKCi3YpNxaDE60iW
AukfCemgtSwgfAQWDzCAX1WqORv7Y5yoAM7hdX6rHwaLzRe0tmrazwjuq99om+QM
SJ2Y5WCCQn60TsUY5W+6v8kkRaxR1Ir/E+nLUk2kEMpmvn2nEl6uFZXy0KlBvkaf
47UfXhuHjIGeql30a1laM3HjL84hzF8LkkWflFOsrHtdhSum4bjm2zfqRrVcGHi2
G/tdBbWcIKBZRI+Ltt0gHdoLpL4Xv9zy9xh7BejWu0p+4N2uAxlccP8yOgekXI2i
gyA9/OLSr8V+b5cCgU1qL4Mh42BfY5xnjKaxwaJLVHC/x5Zv5qb2vDhmV5IAgjks
xSl4EBGoWwc4q2z2OPLp38kYJCBZFkTkXGSa+T6GKWYV3qG908BF7Sn+r/S0fGMM
Ays1aYxCVDtD/7/vodzknbrXtM4gLxWqEydFBd+ZLQiGIje2QWcMeijnfy0WnwxD
pnAkt2DabXVDzF0uXQBkONn56ihoB7vsazbbws/T8/wZ0ZlVn1kuy/lWQ1eUXF7A
iPKHWHL4Poinacg2Vppeeo/HdFrAe0Q+uEzHSk1Sc1OIjOfMCw1JyLyA1Ydzpjd6
Bv6OXabNYJpu87+rZM/D/6a9CB8Mx5cCiggXADQD+ZeWbY/nChA5TsWipKtMZFMv
tNWuKoCIfWJFRR2EUs736Otb/gkfk+2BpfuUmdVaOFgSoHQC2aUqepL9yuQ/aOWU
HNeK7GRcBbNPR1hH4cmY6i+5WTBn/Me3isjmR7L7aRV6/wzJaPd5vknwp4AT2SHY
u9wIP14Is7ebVUnGfbZNBWLXkbzeAS4xm6KVYCyTEJT1TCUMcTx2V14AYckbJ9QP
Aq+ILin8S9/Sx+2/xVmapnLuIW6etlm2MQT4sZUYK+XBUgKg9tx7Xp1Ck3jDBNpp
V9vw5FgwpH3+hq/SLMTuhZ51GnhBKhdVGQMt6EInk0Bd3+0IdxAEO2QTfqo/z9pp
543Gw4a6n3VBMul6QXt6mjSaRP/AYzFRoF/eFE4McWXSo9dulcyr6rYE/kRVCAEv
ZcGDGa8jbjTReq+qVcoVRCkNxAI1ea6zbjmuhVyVPpgmAp0Hc3Ckwj2w+c9mZKeF
gf7YV7u9frMICpqS4o/QqTHiZFnMufrtraMAE+H+UUQhAjTziFF6N4vKXvKJv0J1
03UppSuY5rHZtXDfIQNGFW0XNYtBRxUbG2JwcQ1dNnK7FaYMxLNQthdGojKrreqN
4ZTIDKEeymiA1U8wVrtU8apggw/Omv9rSHcBCXyyBGRArKvjW0I2AhRmpTC/g/Vl
7JMO2PoJUAMSb1+2i62trgzxIgt9xoll8YvHXGAcmj4/nTNwlrHymasH/DHwm1Ps
v8MNKEocqvJdv09lhLSi+eIlZ8EGFIX/Wh69rbBUcSV6UCU3/WMvrklrSRdTKjF4
nRcpQ8qNrwrkEHtaPQrNKlsOarFLXb+pjlQe0ZgyDsduD1r5pwYAOtZnXdFpdkcp
FxtSHBdvbUBQ0nKSiyHDavN4wPsrrJrKlZy1sKZliTBKEzLvMx3GZw+DAK66UP8z
lkQSYyFc+2IER8aPFiutEKRNo4FGXk1cAtJzpHqiEeGG7oCkMRUc0SUOaKGChhtP
Ib3jWQLy+qVE6lmICKyunU5EHtuoXP75shjI3NuHq7T0hezAZxoAkDcGzsRbpwoC
ewkQneUFpP9EUcei2cZdsv9+/tcW3HONE3hLOCmbs3pY/LsrUFQQxJrykZ7y1wr8
bxV7tM4ht13B2zw1Hzo5E1e7iXcdBPdLAvw96CQqTzZB9mzEyWW7skghZ86qsTJS
zbgaOkKQUS8MLKERgpjmjzMkHFmbujaU2VQ1v7kDs/fVPvWAuJieSfDb7NjQErcz
sDlN5OqDHSbfTe2FSwRHcLXy2mGRR+q1h24CvP1F//+WZYWBRTLXnY/dep4Zu0fe
O6YvsjaSUbr8eZrebV39Rg2Bdu/Zg9mf0LYq/3UxU3bPjnQ1t/wn4mQaGzJIICg6
ENsi/LVW0weCiTv4UFbezzqAe3CqySI2EtKqLkdK4Us6MP/UWOxtvJ5j9j/z0dXM
mnb9ueDHymq5SZP1w72mCAmr9CgxAs7veFLkXBgtdErEjVbfU9zauDzPmgkr67P5
QhG9SOvh8+/RCiNH0FyDoctfKOjYyhkiPtL163giAiDuHUJOkEkxk/FhJgfpnMwi
UnzMpuWA2Rsh81fth9dhh7YNIV1OBhj/bSGRBNp7T520P3enHc5Uxf655w9jLUqa
M/dTySX4EDcL8fs4hUpAWDlPIjMOf84UNag/5MdbTFTV/q0IO5YR9+53OghjrsOz
yiUWXDUkackqiPFYRYwD41lOTZiDDxBOOJVh8gIOoj31I2TlC0vFH/v2xScJlnri
Wjq+BmqokCgCJ0pj4Rdi1IJqAtlsJz2Dt3UCWtPibZcqOCfIXRpZyU8Mf98tI6RJ
AycHO9qhnERO8IJcruUPeC3OWT2+UNh75ynpHIg9mSasFzX1MJ3sMfqEAg4rjDJH
JBqdzUhFlJOE4SnMHAl+TU3nzWFSS+J8u3HCW0jDqUSIDv4lncyejLYLD1NsMUxO
aXSSGmXK3jOEMBi+HFvyHzlSlQkWwUJxzHcu0wWEa9EpUPBV56o62cTCK08E1AD8
AVAbT1//BR5KDCvp2ADTe0W529lUXlV+VP8ib8G4z+Edpt2vfhRrOtiKBGKXaFvL
mzOmSCDiLCqRd1QxTzeJm4P8FXTJQhOIApny1arYZuhE+avyJLnnAKNCulkvH1n3
DE/dn2/dWb1LY8QsevXu2ZsAufgVET+ClBd3OkULA1y23Oer9stD0Abi440ZD/9K
oGBnRX+nY+Fi8N8D7z4uPdUKPzUWpQTFJg1UPK3B7t9rCVsG/PTqIdQxjHcqkKDu
QV3iS+fznOWGY70RzYiEyqiNvnlpUwvGtXLB6sWJ0Ft++2jYNCf+VVSo2wpgS3Aw
d53vbqpsS3hGfcKMVZlQXRE2jelOhJfiLBHV/M0EZL2P/4raIpl5DVA9q6iTIGvs
aU1pdEnmR10TLl39unXK3+kYwtlkRlLHnyNKZz4Udd6ed8bo1tEKltroMLcyLcK4
8/CvXGhuJe5Q3rms3r+7MKbbjzCHvK49FLl9Rp4S9U1NNmwIbt8TXSFi4Jsw62lK
KPLBA6VUCJJAVRAhiygdPqvqp1cqqH2zVj1VxsgILCjsIl3QKAvfRJbmLQPcBUi0
Ovr8XnRJZW2r254ukNmSVvYeVT3URXQb7Bd7xjH2RPV6O3QTn7Txdx7bcz0xC6fx
vQp+l/sj208QrHQ/Dficl6aoi+sBenZaUeQ3j1KwngWu0j+p8UXHJ28ghByrSKd3
3cePfY3OZF5nn/vNTOcNBAeLz/gRxq2pR3J5qQFH3H9x/pYC7J2HU/Ufkm98V4iw
N6HlleKuLRnuVPhXo38ofgtIfA4+5OJpPQzqNyGsWUzOteYucSE3lLazRLzcHv8K
2UQTmZubQGz0lFBY+Mi5+NAI9u9bUHRHKKZ9w8iZpLO0hmo9+FdRwVKGpy+ecBel
GCgR3dj45Zp733tQaLaALJTvOS47AZKlv292F01FfQCsYwJp+Lz3G1/bhAftw0dJ
D8PTelEoNpYC9LqE9eJ7O0jHEdmbADcSAW4ZQI+6DsNhgsEhRRUXyNc/D0PoAtsI
diDQH9eajQAgjSdOTi77UCjrV2JRjpIryAkg+MGAa1c0/RKzcAdbHe+H6coa5xJC
icxjKCF2e7ugSOXvFmgqWwR7PCvQPdIgulIyKpS0EOvlDGUB3rJGGXGUP9t6evfO
1saH7ZOZCDkzwDSMNhIb7kHyCaPH+KHUpcHtG95zOMEzliIib47K7YJwg98wR8+G
wOKM4i4b09X9YiTIgd/6MdjT3AQMNZDmhOUyrIzO7jUZTVFgYHrOr1PlfNGybnFy
Mwyb0FnV0KXHAcNqgZEDmLVIMKM8ipZj3wYAy0Tu50z8OEZOrLSEVZfnTjfmCvrv
Rwk7Vcv9KohyMgawfcB/r3KWGFz7SVinOfFSKouXBCJxJOWK11gTFWEylw/z3F2x
r1SUDaZp8lzLd3KILw+sKF4NZY1qZozdTHa78cBGB0CR+RUwP122X8lnK3nBjOqP
Ye9PKkxW7/nGKeI66AMv+9fT8OSTQn4zhAJYQL6/waxwgO+Lu6UgC9K2BFJHCR2c
rtgmpHWBmav9uYymQZ4GZwaNQF8hT8NoMOugyQTSqL94fYXKrL5rrFpLMwz0IzvA
t7N67i9Ie/OvxjRn71p98JzvLjx9smDFbiuaEsvIZpquKZQkOBuKLs9hqKr1FvUY
UVOlQwSXbVFWbCPOUyZ4Swez36b6oS6+/EHd5eEe2aOPxYuk98bagxUcd3POjY9O
Ot7xPja8eia80Kflmj74POl1hOUFlnV9blAd9LjsSU8R2WL8/yoGK7vI+N3KxwzB
hi3/Tjjq7fhr3nR5Uk3EHGbq660EKg7vcFG2l2sLPGP9vNNznVeXWfyD16ND6g/o
c4ijFkQSu47rlmMrlgasBOWYqm7spXgBXcuZmDo5MByWEZMOmYri5NfT8K4vRamC
2bCKoavdV71Z4VSkwYX5hYJeTLIKS6n0sbJgz+6oj9Yy1Lo4aLtNHrHDVV/AEdYE
pHyHyETBUcUEvZbTbiuhJPvz4TFCuv3hQRUCLfz27of9Nf+1cEAzPDEFuZtOZsCs
+lYO2sG2nR0UwdSNfeV+ZJkeuBqQzAJP9AJgKR1FKnj8T8XF2BioXIkwiV0SAKgU
xmREm7fqKjzzhGuJfxjQHpDixhvW2J4ygKVALc54fViCOs3NPawZBIv9Y7/SEwQX
lJwLp/w3ZLnA7Q+M1DxIGNmsvF21Hu1utlXbLW7nt1rBi8wGsoPOry+igEBz53Z1
CZcy3xOzwEmkN9T1jLGWaQTwWp0qgN7LfKRU5LvyQfU92mbzw6e8eRRGSw6blpdL
iX8MYuewgFzEpUZpJfu+qDgiGqbiebUQBPuiLgAs9JKqp6UDKJdt+7UISm1Idag7
aA5omVe7mRVwqUT2I7/zVYG99CeKakbX+Gc0EP9caPn+1SAdncxUua/Wf+Wdf7Zr
yoflseB1YnDzll9Vxl5ictlt+8TPYF2EyRnXl6uu3prRaBufD+eAxShcQhKgAD9X
FE5EILUdy29hrP3HK2E+aOcV93LEbQkFapKkwS2QHSncormO2gRtIEj85EpRrGmb
Z6T51hIt2JDLufGo00gy15oMI6A06ND3i7F+kPSq0QvD8Og7FJdXklk0ZrqAtyYY
sgn+3HX0t0e8MJae7ZZm/ckx1wDs5cI8WRofbXDk3Q5PYQGOvS9Rcbm0OIPqRfxV
/bcPYjkpQUfqOIeZF+Npe0Q+TWOMvlk5IPwF6Yz/JAA2xRP32xvKJ7/Ag7dbj5mY
C8p3Wxs54ejjo2uaVhg2MDFgo271f+pxyjR1khKvYksu9V/E4roo4Le8jSs0y7dh
emFDy1aTTyaNpGS09YulAOxZY7Rcxa6xB6RSE6HaQa+JvYagHbDhervWsKdskery
zRZEXq5KXs4pEJZiIQ3p4xbp1ix9WH2mDgtF7uqtncY+0+enhje6i3dETOA1zwo7
uP3xGv1uRRBC5zNFnk89I/0Zu70nhv1CCvTeyGbRN6WkRvZlChAiCgmiPDtvzR+A
WtcICT8fasTkFgk0+MDGpM+tUPdfOFEdEO0mY63blgrP4gBT0i9TtbL+Je1Cwb98
vvQok1rzwWYzbLnuD6S6Uks3ISOMYwKU0AQt7rozDKe280zRSLSkPTohRJvhHTQ6
TKXPlkvqSe84kzWjRoZChZ2sJxEn2i76cPHk2qBo90dR9Mc0IH0KQqZLZrkn0Gq3
5tJ40MIgeEYMXI8l4V+GYbhMTJcynxSGrzH5O1xUvDhjrUMldCCHjKDHEgXJEfyV
j1HDbP6B5gL6jXfgT83hlkE+8xzbwBFIEdboLRT3i/JNgYmlw6g9Uq9zI+RuSq8C
SjiHoe09hWAp+q1L2zm21WdrwhXrYM2R49nyDpluTKCFwN6busLbF6raEUoRBaRg
6LTbDjbhmA2dAMkW3RXR1dVPEjx+LGsjLZWQtEMt6E23whvh5mYXF3Y9isoN7tMq
XffJ5+VENSCUUE/rcSc/tt9Imz59zIzrcW7SwpbPCsf+2ucAiqI4lqqbVnAftRUE
LMa3i+WT//X4Bcgel4tMY/jBbWkTs6fyNYkO2MEKT94cbDwtbm3rJ5p+elHPzUSY
RCTM3kKaUU2Uyev6XnYQHrY3ZElYNf9eWvaoavpSFojW2xw6tuEd0IiS2hPh4GrW
PasxXUrXuIGoX3hql0ut/0BbtYIZ+M3iCQ6j0jfKCLNIPkJx+EHt6SEUcKy4LyeZ
xtTzwlkvsWwJz2zZ88lOMf5469+U2052zaBUwR7JK65YGjK+88hqqGNLvm2zS50D
i7FJTGwxhYzv4prMWPHGPGm2+6SHHrCMnt1Yb+S90MZyvr3dN20/AqXHGuJFMqJR
+9G6Rsgue7ue2DSPdF7SiSoAuvTHXcHVJKj0PqyYmiNbeofrm3/Q+EuwS8VNZV4V
zdfkI39iF8Qz9HErCZM5lavyAupvBD+g/stDm8WZXt5XXp0nmvskP6EDcDvbhnZM
NHQ5NmFGJp3zKQ6Tg+9RsfNkOiWYS/oTJNlJBl1J6Ld2YoaNciz1jfGFkFOBa7kd
Zxz0ZDv4rbnAYWMYPSCZThS+yXHz4z/HQQdSAn9apcDuyO88sM14wWL6kIfcdQuv
vNNcaNnsn1nb9O+er3/Gz+cP5DpeSVquBbwQlKPHym0RXl4PbD+MeRHeFCagqEFL
ZaO/AVYnNlsNB+ze8L5vRGA5o2tsZc2vg24O8Y6PjDBiLIAAxIFkTTROFGYxdCSr
zwc0JJNjYnryp8EfPpbqKR14lhgNqtK5ABggTgj3cbuttesRZv2A88yZMtupVNXq
mrHT4Ahptb7gYo4U3nAiTvM8gLiQ0g2xAlI5S3dKOY2yVoLutIsfb8ZlF/KvwsN5
j6e8wMZXU40LCYgi05IoZH+ozmzL0I42BjMiHFw+RnLCtgytjycohHe5McY2Ncox
JmthUWfM8RZzxBfpGU47HXz0o+qMnVDWI3A8AbkwEcH/mlAnOW5lmO1wrJgOatzQ
lcdyq0Vxpvj4SwMEPh9tS/VbL4dqs+PJvvCFXw2TtEenMTGIMB/bFOqYI6lnfJQa
MqtkFtOq/HLD3z/JZYDXB32H4SlglDmVquBc9ta2Wk9Vp7Yx0LtMTNLIHZLG0OWO
wIn1+lOmXMowy2Y//47PU2zLb7f4RVZ59kkwlpRzO47+5fFFKvZK8B9zjzRYNIbw
u0UANN6lLV0tIe+VU6Kte3Eeiq/ufjumdCH2jiq1zkpMRf5LcevDlNapcwL5K2HA
YROjmnwL0397NJiaBRtb53IqAJ4cCZXsNkuOSlb85M8J5w7EFs3Eq4RnNLg989c5
jJJ659rbxxgXRA3qEuMrZWW3n462E4TIXpk0SZsDAdM0NzITrkjO95GCeCt+Xqyr
cUJenk/+yr5L9aLk9u/EYo13XpCe6k4EynUkfVLMZMlkUCQiPW27wQYiQ/uvSxVT
C3QfmMRRiKpx3X4wJYjriQJO5h1mFsuST3Q2ZRBe6Twy4DmjjyppaXYCCY6XOcNG
7oQhFKARTLrbJ4sj681xWVZjx09Iji6XCXjPJ8IiD3JUo7f6z+9p7Zgt3PgOMlrg
HA7D0jaeQ2DZ4zC5IXLHXAlE3numv3/9YmPny5vwlvXlOAt+YgWwcTKQBzboJC1M
dzCNw/Z9rRUNPmmlTRgoUVpDUXtZP7GjfgHCEHEh65CWLqGcs1sZfSm4w0qePMHn
OsHui0hxM6VWFy7ylhY76Awg58sMmPoxXh0gJxN0voO5mcOsor5BoNDj11KG2yF5
bX8gaL6h5kk9Sw0S7i0zyr9VQQuU2Imz/2n2hdsL0MikYT993/U2uvR4q7JwzyUF
RF6x2nYcmyHrjXWFnkDANlGGtBF7KONBF9YX0t5bOwfKJLJ1AfbaWCmWxszXDEOo
boWFP6ZGttOVLSM5EA5rf3nOQiac06DbRolUZCbtVBD20OG/B8IjDtY4D+gfbWfA
CvHVN6QbE3yk26opdtvA4gXezCcjE35OLgvawgig+hNul8Eaz/apwqtNwOUqGkjN
yYv19tYUKqQu+RrN8U8j2JjlkfM9xHBeyGgu3DOX8EcJSBo0PIj+CD7ZX4LKeZ0p
FweHb/hKN3FR8fa7cbAUQCCxoto8tq8AMHGFpMwtw1+7iITssJ1JDi798i3hlnuU
8I3yUo4avl6aL+/r6xe4nmgM1MmM6TVSc2gELtY3jIQ1iFpQeRlsSm9RcZbA3Fez
XsdJEuJ4FQ7awnm3JO8GgUsgEQcmO3QVMptLH5sbd3YXxorB2ZgPdH9bbSDomkJK
BAlGQA6d5y57OYS8DFXgr3Ou5F/C6CtQLJIs2cLew6I3L7j4ojKValDjHTeinGb3
8wmQ2TW/pepc6SENUSkDZfQscw3lp46bLBwSuGiVe24Ax1Vg1gB9ik4PqKUALYEO
APjPXU7wKDJxvSsjTzd2wewwJYTFylB9G4d0HOs3WB415fqdjwbHPiFczTotxJi8
Vh9BSP0Rl7EGOZyit4pLqnCbLS7zrdHHrUkMUJJi1XcwF4fyDUbA56FeoRuttufl
bMIecYnD3Pt6tHbrTvGsNJslwBXDT5zTp3O4GlNWXeH2kJotvxyNGQs35Pja/wMm
QrxZCDcfXjOpjaHYH4F7EAEPhr3nsQVy1xufyJu/GtjyHmrNhnK5ie+JqJJ9VsAX
RL2yfAVfP89FsHQFy302EU+1xnC/ohr7FomqKs56ss+E+USewdcI/V+unfNO7LZT
KlB0rxk9rDoDeENNCA08xZ+s6BbGSkWvqkAwijlI2iH79APT3tJqfWySF44L3JVd
3wySQSZdr0XsKnLzBItE4s3u16bbw5aLoJJbA1+Dt8uLkLP51IYApcQkmiUwtVZP
EcFINqe6Jqy+X1tEXyORg6lr6WR4d8A6oK1L8wxKh7kdkaPQuoFEkOHBZw60ZCLG
CaJa6YhDXX5Co310z3xwzBhcKGZSx0oF/DtP7z2U0rhvspL70auvcF2ztPeyOMrx
MlLcMWGmxPQCpr9LwWgTUYWOiG6MM3KRLtAd3o8qUFHDZLPyAE6J8HINAK6/gPG/
N7V5c5v86Mz5cayVjIqggfzJgh+yIB9ZY8slDTF9jLtjgO6uzRdmMi4PRl3yceAZ
fTeAWEWWRehuRdLkqHDmCG6SCMQUUdzNk1xh8RirzeNJMyEgogaYTGAr0ysjxT0s
9tbKYpD4PrWTYPQGFHKHGCin2WFLMoxJalAMkv5H0Tc/tJs5RFlX/jeSYHJoi8JF
aZGrf0ZpG9BaDJH9gS4P82HOUn4teiy8XcZhqceOMS1T2c205I+QsZWK/4Aa1kAn
qMHD7GR4VfvRvLhKt2aQUBsmdg1lOYpfcEFb3BgQe0kpNKnkz0DS72z3g4MYuQeN
5vfglX/wO2Tm/Jn54/aHkITvjw0JW/Qmv201x0/B2Do1fMBYMwfYr9qRO0PcCgHt
ofZhFVEK6gFyfbNTEvynE5Q0gik4JG+J0PckEWvivA36H9u0y4sE1GkRZlu83IXy
mX7Yrgd3q94f2pl+Wl95Ex1CX+/0U4jDsJQKmGr523I+AuTi/TeuxyI2PiDQNNJE
RQRFExGoqKrzRCQOKUtBv77S4sa9rmAaHU7ZcY2uyBg+cq89ZI272nOv4f2UHNgI
GDKt+utFYcR6QQ3u+VxH3LnMqOYhVmwx3BXl9NPhAis9u1z4gD2+tOn7ilmUFIew
I9aKOMAIJd7/9PkHrCfa5zQWTs0EK04hN/MVDS9OZJn45gYRMQAApDbwqVsCinZg
8fESBiQohFBI1kf4egGCukpivu9ti9Wgh17rO+DzuL5D5ya1y7UPPHNJ3h85FyHw
9Ul+i7dA0jOjWwIjhysdb6PnCua+xbqbecbtbhXt+lLzbtiCllbapk4rfUonkdrh
DSrgs4f1eonYTSvxfaT5ZdGTjhMfDDb81/Yg4Su0e98/eq8t0ujn2iRS5Deh56sD
sV5HwPGuVY1Ei70NwZq/vEyUj7dmSXBR4IH33UXIh++OlS4HtFVgcLbUo+eYLExo
i+rMqO3ZAJC0CCFmr2d6Vi7A6HgkFu4ZcPXcqqo7TeTKb/nhPlQ15UJOkfxxASe5
FKByyHYCatClkS0W6m/hXlAIZCxdbrVaiVi9wV0XIigxbeo54wxEPgLsLthtFMxb
gCe6g4sX5cdPGBGA1VbwfhgeLx8nvbswkSwH40IIAgNgQoz4hyiOiM+mh3F3F+kr
7TJVH8VovruhWBrsPSTZVYHJ20m9iP21FU+jTRRzWjqkw2ghPVAnMFhUEXu498Cx
jcrEOqvw3prfVtVtAuy4T+Lfemt4t67tOPMvfDzXoh6BuyVAT0H11laFR7sTsHsf
mx5nQ/L9e0tYXftm9xV+VKo2z06awE1NlHygQQafurd7dW0tBhPHid9pky8Sv5kF
/xjydG3Qxd99y6ZzKfu5l4a39RKemX8e5RX183xSOOniVIZeFUBHfvuHvCxhuuMg
1PIGf4IrGY3peNAml1uY4azoCqBDUzCntMZRWKSfXZZBcsvdHCLSnZvIsB5amQmU
d+EJDNjqTkjdyp7mumdwnUK3L6/DhQ1xbrCtOm7ikaeVFlSWaHVpn4PcB1kiFxn0
TIE9rxx1kiY246VD1onbaEAJXprJ9NHQTQgKZsAs8i6QaLz2t1QBtuproUTbOSuc
AJT21Q+/Lg6xDzyYgzPTO7sKi1+d9lMplxyxvf9fBTeiCnbb6n7Cvuxf4Eyty1ua
5GLPRxT7NbLaLFudAp4fYTQs2GOR4rgiqyLdO/hZF6AFNs6mZkrZsrp6Y1K4bIf5
zysve37auLCfi9j40qcAF+DQv2/cpH+5OZaXFjF+OEzywb7mDNkS++azQlWxnutj
9MefVeuukBHwYf6jdxH2PJEfiuGTVN032v2qBtmQsEGIDfoGizSwtk4XsVDMQZJ6
0JuFKUd2P+QKhT+7BFYAdHbWMT3/NCUyQ6+qm7N//CNs6NxxfO1HJWzKVq5nGLMR
vpGh2QJE6H9kAgZPwFO5GAunw1lnP5DzvKWNGObklbdG39NkFA3kTO/PkhU1hmqT
UsnuDDlQy9UZLhBLVZkSrhHMhaB4Qrivd3xe7jzj+NZtU1Pn2aCIhbaIzS6By51/
XEb+7oiLi3DFWsrpQ1/L7PsraNSTqFPyMQREE2lE4BpXzxvcIZ8ORcMh36gUaNWV
WL0fEc+outYsPXCIvyysmn+dghva+lEI+5MgQI+hG2AMKq2oQU/pZwUC1eK9efDh
nRRNNe3yVHa+c6PCHM2z+z6JLxIcZvPV4wAUMlVbGjCv9lcDwS7B7TQxXpZOzbmQ
/cFTQ+KtIxIsDdblLEwcCXpLVSf1GeMW5v4+gwX26VUfWRF5gz9PZXEBqRwVHonp
baRIIvNZiVcJ30SeF35KWHkZDwjXkDN2OgdjvyjrUwu9VDotA7OmMcxhU433yXSs
P+t7nfYmo++rmUVBojnY4wpxny6Lzw1BzrMUI0Kdlbgshp1dE/iuzv7u/6uYEvf/
H1skKZt5GM76NLuC3qmmXZy1PKYfC1InL8mkL3P8QDdKuIKhkBt5EooT/DR1Ti5P
f3fUtXqr3fJ2i3Mi7rC38kJ7J0qwAnOlu7X7vjbFVTqQS2D6sy8LFEsdogCke6pp
pbZCajR3SsoeZre7lT8DFWvX+RhOFDI6upf6XeVDFNyIQOREzHfu1wnu2MnVd5/D
JUuuIwjFf4qn2WR2sAENLMMW1rlqMYnPgqWbMRepJBkcDXuRpa2N/MoNu2mwfFN6
+oA6vMARRzn+Nd8zZ7u0BMXmPeR8toiTJ6ASeMlETLN1pCLZ6jAmvJciqyPT717D
xaUaN6ZE65/rv8Jwtb+1od0hSgt8aBUah2UwIE8IOe7YgUghdOUbUyLTIoJltMG4
3Q9fE7fmtHvbc4FAzzBBdxdDyVMxWgy81YTKXTSQr+Rynk5jr1VAYQ9Hz0BQDEGM
R5sntBE7L/clTZtxcqrABzwDFiBSlAs25LDfy8OcZxI2EqxPRKGlwIitUKJHMQxn
/6Jx+DKzew/1ye45kU8XWlaABqHie76o+igW3DeJg9rOfvRr66RPNsLgmfPFlddI
9dqJK7nAaxZJw1sa3kYHBNy45Dw/Ioug34yxH4qWJ62TGydJ4vuvYi6hx2AEFfnz
85Q/ixVjywdS2j6WNR/f3Lgwh7dhn/eDBDUJDEQ17YsFmm9i47u6Go2cyEt+m9Jn
4DVXYcOLTfozcQHT3okRX/drzSI7C0yjuiUL2MiGO8j6/+NgnBSwjRp0nYXZFOdz
TmAAd0d+TUW0VDdhbwiSEdtK8Rrp1PINpy9hQCRNKbfUbhiSivJgC9ZglwR3QmCC
flZaY2ImTNJH6M586x9H4p5ZN4/U0BsEqELqGASG6Ny/Iu2G8u3dOTzuyAqAFE5o
iEMXt/D8VF+7FHqdVhAZ/1yO+jc9/NwvnTdsRDOHH/UPSW1LcWQ37V1g9Pb/aZZJ
oBPIwNBbmre7WijEU+SYtzCb7O10/14AY+yQbSV9TjLbJC9VVuDLOOLo+aEKYZd+
cAWdL+n3E30rsdgIcNxDLVF7hh/yfP8ssFPBrpel4EVCfoxJ6p7zUFTD9uQimjFy
5OM6wOWJL6zoVBoJNnwhjJ694Qjl+MyyjVzdE8Ojp8zVRlPTDFcqdz3Ysa0P6OdV
hhbsn/FvSNArejA5dJ/7swDkJGF44c80gFGCMrHEsGupgZQ1SsfEZa43MEfUwxUg
30t3kpdOQ1g/3VPmCECoI5BrnuAugQj4VhNKx5huwqEqKgsfktvztpmHtQfGo640
6u815HTWeysLubCtWUduiO74nEgA7Wn3Z+uNf+p/SagtJm+pfCbUcY4DNAGVX7r/
QpDUQNUaoliKnChN/WORMtR1QYTgm/Xn9N5pcWojlYlYHe5ejl8Q74sd0AIGP83m
k1usLjesUut0AI8a1uPli51qNuJPDzRehVOXpPRYrcfzYQv0F4RwHE2VOb7Uwkrl
11QgJPOtTDZqE6hpKoBKMpmL5b4T3B/oxCZLpYWD4QeGSMv1GsHGkmPsFHRFre2u
kYjVBV6VrU0LFenwnwet+38B7HgH6aIJs7HPUV84UJnVEczfzKKWhuDQQdmA7GYt
/sX0CJ84hmkciQ7skKdm8C96qLuRbWuE6Pjngnn0pmArHBQDBGzmMt/HNRWXOVt5
cL95FVI2Mu1W/4czhW9skNpRQLtY1Gkkv3nTyi5VFGa4jzN1Vx6MsJZFSQXJjG2o
UgtdsDtgLfhsi+aL1efxymijNZAZrno4jAPk7voX53KQ1jxchm9DXNs6j7mVUPPu
oiFEZpt9jrvaSGeS7ZSR9aIEqLxBTAM+1iqcBXv7vGaG/t1TfkaVXW1ErKRexM3S
GLe0v3vajy7oR+XYT15ql/PQfFi0izEUlgf9gJ/jGVbBJ447+B9/aoP8ttsCzBQC
zcB31Ba8CXBJHQJpPUssOXSD701zk22DCkazQPQyZRtO0rnK8QAKarNscffMpTEQ
4uabVwbpXt6WxoFooPVCXCdRST5GDIwxquZye+XHuO9p5pJpzKWJxCD/zBfeu3cM
Wup/m3ip7QBzhe013IVuV1pvDZLf3AUOdQ89JqTQAzspfyouosu7twiWKbmNWq32
tCfte/lYIZIJSOipaKYiVTHFpapV5GRO4BLMd+I6CNcdp/NiSYYmmYJ78ubNhIW2
Gxf9WfHMIiWzbNVfHnCpKBhPfIp+UaOr4pB1B9iocCmHGaYP8VJbFRCLWBVh5uuz
qOccpPyK3UMToV+HXqpls3T6RFAAqunox091NsBdk+VA6Mn9Ia1HatGkn08IZZ9S
oAyNATWCtDZqxsU3shQRryKZh+SGxwlkq2tm1Prp3nLMly77t8SMzcfV9Kz4yn7E
qbzSkhLlBdjgbvvLHxmS9D32m8m1FvLkXxA4IJ1t5xRcGL/QoasZHHT28Rw5H8lw
lcEjQDE30Lzp1DxA8STIEUvMHSH4Ne/62IimBYymUmgqOgdiZQkOI3hk2EGC6Sao
e0iXuAI+ZsEn2z3eDqEJCNED204EyH0toe6a8FARrrghlRyYnjHM8KFHHoMyW1dG
HNqryxvxgn6Lt76c4scdLAljqc/L9lgrIT6fnEuAy3LpgqHz3Po8OGdlA3eHhnj5
bdjKpj1vCoF4odQv5WJCFwMSB63TH+GJRTmRTTGoVLG/L3XOHobbnPnq3LHBdkjG
eXprzBil/33+2s39nXPZmv/KQtuZb+v6IEd7+bXGou/AUALpHKO6wp3VKXka4fGe
1drCaGLqfDiVHgm/T6Dy9ksZi8SFoN/cOgFw2xTUwv6ZiSXuPZDwfL8zvFRmsNOj
TQihhD9db2ZTQV+IqU3mw3ouvcr9v0t2Qx66o3oSms1/0qGan7vRVgpYMdW7kpaS
WZvA9WhlKMJauuf3ANnaWrn6ir/W3n/bwjUNmWxMkRGQHlz94ukc7w4UipEs3kJU
vwUUW2y4uiWeMATq8x8qsRkhzBzLEbZa86qaj2z7jVthy23Xmnf1WwM11c4tvdnC
+EarnuWqp+sLHSgp2cZp8bzx54lSunE9+EjFj03mZ3S2PTTgamcO1ZmasWUju86V
RjZIyb75ci5YuWXvGzYFWtJEMbBGUIZP5kGj0UEVcNKIM++NSOCZ0Fh68J2cQ7aD
iJ+sljjNHmEA1w5gW+g84T/dzSzXggZteMcp4SnJcNZNcQ8DKjs1Tz19y20k1p9b
Py8rr1l3KXWkUkij/D4QyH4nD0iVnY4/kfTqYNUZ18N+dx0OkrRyCoK70eTRVe+C
rekkgcHBetXwoErt5AS2w6Q/i+21Ed+JRCoT7vQl6iGRLw5juPiCV0j6qWAPvLPi
Eplzhaxhi3yCKTEwJKQWrLh/wf1UR2nBXATSUJN9gY67qp7yUiXs7SLh+0TFV2a2
/IatoBQhiADnWxwHupTdv3SkbGk0v40kY5iApxHrA+wLyMb/GQRAzDtwE+Vd9GPY
Nj9O3ZFAS6krZ3H8H7ef0sj43FUjChVZBCSexNDzGm3ZiyzTqPDkBvOBRB/d9MkO
Pkj3ajd1m6FZn4qD4/NI1635dRw2GTrpgdy7o05h8hLcSisf1kQRwvdq+2dGUKZP
E7RDG+iuG+WAVXgewaCvSFm8vN1douOV/ISFGaNUqD7+VfELa4H+H2v+injqLma9
0DBJ46lI+oLTsjZNaOoUscMjmAlf9oPoaTbvVsY3c9xzduKVnQGgblS+K9EHlSDT
9ZHjWwPSNh7zk4xmS4QfLr7lrZjroh8DM3ePWVKFedsoqDf3oBkypqwrShhCFVfz
Ld5CAjPORuMIbJ9Fl7jPg/5gCZTR6rl/2xfRZIpvwongKRzXamSlm2QIgKo68aai
WcxA8QzhZDevC8pg+VjhVyFaTix2a43LX8Q/kfew2lg4gSGNX7wP9xyUZjTakmfm
ps7uGo0D/sumB/t9AWdONdcz9m60/ihkS+pQSWRtbr30NQqmSHRIC4GnYVqXq+4R
yD4qBGfQMu9sscFDUj6+5DdDi1U2YeiCb4UtktYvvNyy/Nowsyk5DMswSjwdgDRR
7V5fEemBgiDBYVukKv9Q5IGiEQd4PXwroXO7Dxziim+hiUjWm/yH4g9nZDXPtX4B
EzRvprNXyh+4qUi81eZgZyH7iMP5BokUqhY2TKHNtEaMkire8r0hE87jmvPeVM1U
vnFyf731MFMfwDlbkjgQJDufiYmyrfwtd+8RJndKy9iE6acFaOfkAOryIgzMtBM9
jd43cPqiakfdbBGoFJAt4lgNta4GIpAE/4bi3bU6gtmJD8shGFtkscEKR8c7p1r5
fvk4fekLAUE/8qOIHo3BCUcUW1nASp1sV4Sx/7J+APikZmUgBOsp4BUAnhOxmGOP
5NXADXr432Py0U3ox7YVm1f6OhNCKtOGcaxyoZyy9/oMGFaCHn2g6h1epCn0CBVy
xpbsWoJpmYbtXJ3gLOGvGlxLXfUh90EIM5zlMwuG4BFPKfV20Ig6Y/gM6dBafDMh
RUKbmmqJJNbbBI/0ZdtwfrecgzrC9zUxXDJx6eTfNjcmFPylgeq5nkmWKk+AnRIg
k+t29dT6TaEllL4pGdBjYEagxQfOVN/Bm03j/MxN32q3QNK+IeuUYzoP1CiadT5H
ZDS5HwsjFRZsCgCX+09uz+eqj9kOlJ7deKepwDz+niIXGZ1bZ+WZe3r/iNzS+9eu
l7Wzt7hiblg5n/v8AN2X3yozS9nTyceei1fNqgelMdV7vPEJINGZoEoYbnH9I9hb
pZWWnzOohBrXB5KmBv51qWLfNDO2hDXU4C2i4o6/guM1n0Z6HEzKQqPqgW9KLnZE
5BM7c7VzsXNkg0ynSmhAltTPHHp8LNe7UqEAre0LGs/YAEyxFSNjk8OlSoVAJXBF
aPyFy8wPdwPpMK5mcMSjZTG7MnabgPgGD4rkM3jjbm1EHUqn/dKOrpaTgOfqdvt0
GVElE5EcCOpOvRH46R9yfkYCpzgtc7WplCN2VUXutzjR1fzzs5tS5NpOBiMJGI5T
a4Sjuy+N/gMUHATewZyTtU+IqcwA96Kx1iQQjrvVtwvT/X718suZl5lzTIy42lyI
J9n73VUvfM6oQRr0r19+uV2M6BtF9vcZqh/hEQlA7e2kIfFm98wBePJY9STyDngh
efAjmXtYy1Ki4dkdX6QgpV/WxbRD7k+VQq/zvDOhZUYE7FDOxmp/jVN7Vbp4GaZd
yQ3PmTtu5a0nUPZHwgYcOu/H6Qju9TF/DI3cUcvGgdtNs4zRdRvIuXK++ViAWb81
Zu5hmt1aFIjW23Zm1NuoQJl5Tmau/VHGzQgppZO3vIZ8tASp1/aRJtHs19HakvwI
TW5q6+QZs2qtau/YUjCnd49fhI4fwYQS6X/zPmwNCDJ2a22sQlfPqYliPfja4V83
7mGyKU+jl46k1Q3lgDq+Ac/y3QYyWuMJ5ifL8KQ994LgeyZwun72EMk/gAnmKirb
5U6BcvErqxDhIblfKBvfIMG8Ldhmki8Wg2PsbwgYIzbhNV0MZp3wJDNAmyMKkxTq
2GDa7eh6VeMbSWSaGmqwTAr6qtL2UrMh6mCgC+JEckLoLO2yYLd8k4DySsU42ytP
0ASUNjOdTlcHOJdfJFTbSjjCRCMJhmJF7DUuCcDlVnpxQtLxY5FC7zePeXo3C/9O
bwZMXGh2ZUkvecs6PuguluwtfdtJ3G/dcZTW/+J616Nkh3+yZre6i0pNbNXaNfsk
yHqZfToktpCnKSAaC1Y79GmiEsfZIjBNO4uXzrEI7FCjgSxoErXLtoHwcaoQxGXl
/wEgUr2QxLKAyBxph6VQLr7CeW9D9vkWH2VEilmt2Q+Qk/JRC7S8QFG0KgJ03kIj
iXTNYL8mkEKFmc4b0YsY8uZOnSLazPbirKchZrlLQRHNVtoqX9uw01881lOUpIoF
dFslyjhRifazueB5/QpAbyu7oo/ZMZgrB3Ay9+haARWGIj8VkJSnQNV98xHlkUSN
LhuvbRooHgHn2O5chL7R8UOBSYz/yl9sdBMME/adaRIQpIC9r6zgaD1Jli2PBwfe
BG6qRY8RJwo1QgNfkDTS3eNN9kTpT4sh2GRYz2ewBXnEfVmAFb3/E6ytPrirAbcG
tuG4nOwMQ7c/olF7X/DYlIHAnEJLGJPMAMu/UFYfabBN8RIN24ihl+hG5iyF4j90
0sYYaiXkVaIR0p1wU9QXzb9DUqYEYzS0Wu+tUejGlSro5SnDItn4dxiR1SuP7Pv0
HVphIsf13TRO4fTxodvjfSU/MYYU6HBs8+ra/V8yt2nJqT9LmXeEW/LZlNPFHOrB
WLDiyGNmadkaOTFlZDg8cwyuTFGnf0Sy9YesGZ1kWoQukhICQ8a9PyK4P0jWsKPL
3Jjaw5xX3p7FLs4UPt9tjmRfXWwwoh6MRtYykQlcrIZQ/kRwPOjyyL99NmAXdZhG
86+rSvq4pInCqNv3MfOE2UFb7RwWLFNINna1nMo3JN5xCGV9+k83j8c4x94mS87Z
wABXrDg/T8e7gI232F3gisBXNeaTY535the7IqQPgXT6Aw6cY/on6YS9l1cWvxXL
VRUpFtjZXy6ueq46FbGp5rsdow/WrRdbTaRPog88dBRr15XBsC2hWgcs9pWbJRvj
eY3iLvA+NYUnvIEPT1A3w7sr67HM5Cvru5/tFEO6K1m4BGc1ZMOA9T+WnRpohjaA
J2R+dVckJqfvI9Cwblw95ZXXYy4B6LO2QtJ1T4ohLDXX0L1VlKTVBoHlMPb3zst3
+fupQlRURjapupR+TBqK+aSkUgT7JpnOqOR7bU2KcyhS/2fiHgX1vF2pZiHjWbY6
lZYH6nccPuV1r8Zb0wHaoZG7gmDXC2Vms0LeB2GbjDBMAvYf5oqrmy8CD8aZUkm+
DxmU8J5gWP4GO05HSM3iq1zFBeLs1DhcWcNIj4p20IlhAhcD5k63ri13OcmEhaPC
d9ROwP3IdvbBP1VByUvQl1RLB02rF2dTPLEr1s05v8+x+ys0kHnCpXUWSL2cVYfv
K7iquUu7fDr364cAa6UexNtwo7AyVutbfTPU1ZFblU8DYXUmQaEhLd+FuQQ5J70G
pdY8uX1cvHbxj8Jbdc0KDjPlfjWhiFa5nS6A4o6gMgv1FD0KkxHihFaE+LDoao3Z
Z2k8kiKEeeNJvNB26naTnRG8p7nBoeeOxeRkGMRBp1/bHrWm80m6hS4tjjJAD3JZ
U2gbL5TWUgWnycI4jp7Opuwq+EERP8O+69isRFY74X9xvZLR6vn7sWQP+wGkBdfQ
5d05CM8lYRMgec+sqDeoYG459tLdyECrNTzWT2csBWQoO9CwXMstRYMwjDnhe8Bq
ahFNXmOLZ77vxTvIaumDSu+mzyQiQQuK5/6BITq5551cck4zUjeaRAxaVLxM7hnK
Z8s8iKlhBIVhAehOMrY7MmQbDNXrxxPuLMUsPP2bmnHrilUYWFJgbquTXNqiJKuy
+UTUWJiY1agGt8TjpxyK952/BDPU5gM6Rde2bvEeJshcUDFOf5in/Ba9sRuKc9hg
YZ1b7ihNQzMiMD7KaDPrSDyBXpdcMx1zeTvugO4439JrJ9+2b39SyeomNJrHwDmo
kYdxOMmhlM1un3jpjCZNFLbFKqgzQCbUD61DKJg5Z9dGuH4at++rQQ6b6ld8kaJT
/lo1ViT1y/g99ztIyw63dF7SVCuRhCzjFJQr9UDcKzutRumZk1X7JHaFSE/6Elu3
/lGx87YF6M/zTuzaXguJ0Fg+uxqLm1YpDy0X7qMLToiQuvXqrNnTwO4iy3qbsSP5
dbPNZ25yi4G7EFOtdX9FL64ZHj53zQJ1+VLPn70vbgqLi61SkrnljJTbpXD65zD/
7zkmJw1zWlx18aXOaa0RIWvNf3BB81BcxKrM/tTZ8XLD7TmaPUgXDRQ/ghrUnJ1+
EnKRmKtncIsqM1XuQl+QNNmjdRe+UJVwAjgBdkQtJdP6XBdfEon7u5HuoguhPGJP
d5oKd2TBHljDqBkSYtxqIbKGNHorWLBCqUEqjxM9WI9bK2UiBiCC1cOc5IOpTnLq
7jpkWq+wgTOzo60jrSbz72V3/wA9R7nVemL6jDNBiKcCqDuueW/79JRvSk3m+VDo
oL4OQLTYfAZ0r5JbHdGaKzZmEzFhbVE//4pqNMvmt/7ctT3rJ1szg5cphdNlx0Zz
yIJ6M7uuL7bXDLDVZAwzYVY2PY+iXT6ZCMtCI+6d1Wud3U3fPe3Qg+MF4h0TNIut
YtmkP+O2Yfo7c76JCgZPGwFCvOHy2X7ER1dQVwb4d7a8mHIvLebDH9ZuXPcDMHvf
UA+pyeaq/JqDBfOMnMcYh0EUm8vmUltAwQ69Sfp0Ce2gvxlUBTZ4AqOmueoy3jog
xaZVEpKlRNvagcRMYoKCZc8rBttVEQlllr8FBM/v8erHnfhsf8yihenPqes76ibU
kNitTn1EbqyGBQl0NYztL8xUbG6ps4Hx8JYAzkwCud8YV/BpOklwlPWqO2cd4yzm
CnXeB84UVwm3fNM0hTsd+sakskHzPPGjSkKGSIf7GO98GQzG4r6Fl3Rw+mT42aMD
rV1zYHoV2WJNvpwQKi4pfdjDJXVEimtELP5VFRE3Mxh4dtWkPwJwabIdiuoOoJ0o
C60LgXmw2cZCP10VOkfxoo4BbdqcgVxB9T8gvC1+hNN02JnFY2BH+9xx6vpX5biV
zgQjdU7xKmDjjxadR6kCXfezdk8RCRzZqFuUnpPTTqiAtQOFgzd7BAnxrj78kT73
zg0MsuFGxGBGPb7AX3wzJpTWhOn9OUhteHMqGg3Bt8FUxB5SqV9byKOBkxhLb21e
9q7Nx7wzMCIIt0Y+K7aAGL68zLcmBkwkpB2wbFUw6/PBypuwSYQutRnT77NBWNVm
N+4sd9Fa3DfL2jyrddlP2JFM/WxJRJ7FBiaaIVUAEU3zt7ktAtHtJrP+plAut2qE
pmS4owVZnDq1xfqt9/VGULFi1kWuaJvGNCn22dGK2wDj+MUtBAw5Fuj6EiaKYv2c
JC7plpPUoj9p49m/yPLpkx8e7ph7bXz3Q5tqQoMVvzW+4gFgi2GVA49LwRm8ldFM
jaSMarHPyWz/WabTxVqvrS2HHzZfu0ar08QXHMS7d5Tq2qa0fz7FuDbDKkjnEnmD
uyZbCAr1R6xc6InxuuX7bcE22R5HmcNghLQLGjTXOLMNIb8fbRrZlvp3bCuIWmJ9
SSLsZnsIJiV+cXuWTH/pM+SFae80ydbwvmKVTNXWR+ixaY1kghECHnEiu3gPGhGW
jaGdpVAFzc29f9frfBrk3Wl09Rmf9Zlv933rKKE7YJL6xqZdmLdtMkMWbATpNm+O
NqfCT22aUcFEdQVQ7NqGANswG+A7mT7biGUMhuffoB5Ofun3WWCOQAzDbeZSBtY2
zOQhbrXSbklxhNe2ozCDug//cylUAYaP+5iYznQRj6NMcq3PB6OsvtcQlVAWaAfd
8lh0/J0c8QWV8vvJi8mSzLvmtEuCo7YKAaPrb0x9PMKIRz6iYlZwvu+ftBUWFejZ
nPdxe3LIBK3FxUYyori1+pdF4IJxnAxHFc55yh/aDxDg+aPsKLE+DLi5pDPz2BQu
GyZcqAmxft4SXL5TO6pR9LfOmPhBaXi1cHjdKo5znw6pqy7CUfQeqyz5rYa6aV5S
d+UUIp2qmkZ77Y0NIGx/8ZxOS8T+ObEhEDLqOJZWMgRIRr0HofF/Cj0jFqQJUDBN
IXCOXzOqfCDOBHwz0BZlz/se8wg4humzEENVehU1VPUvgtwrB8TPYfZ4o3qwpVB9
xoqqedT/PtZjqe6enGLYomVeyLM92j0ohhtL6kz1twSMYdguxs2+uhMBBRQifa4N
0oIQhiXa3DoU5bN3XKtOmbGxQya0fAGw3h0IteK/gcDwaZQwxQhaNOcAk0BmiCgA
Z3iSN4nErpA93LgaWgVpo5s0udyaU00kwCWKiLWEjH5/0QOtBSJTW8LzoA3XnE5P
dJbVCQ/ZKsU+FKzNb0tf1Wvvs4+ne+Mfz6hsolt2FvG7R4C01weUYvWBOkBmsEWM
gks+OZU3uynAWZVFhjzH8xLWsEL+DhsECF0uEJWrVktT8QZcbTAWhcR+4mBDEWfe
kzV3vcCT2FmhMBdd1OUiXcTs1L6BrLlmf4zv202CERhBrOCgDQB0M+1rzqNHsfN/
tvYzUmtPckOuzKpsrPdAbESuHOxLIQBb3G7lv77HHrf9hSJitzE71w23zFCUo28w
B9WCAP1zzUH1KNqjP8wo3TSKwrK0mnK/7jl+03c/Kt4NXF+y8n1vrJ+6e/dcfJsX
GfU0ED38uv5WEIov7B4L+IHfCiTkm6R203iPPwmLnUBM6rPaJ5yq+p9fteGyN9IQ
DoaZTX1XsQ5e77mAwdKBDnkQ4hfSBsBAjEEIDeHhKN6RlYMeAPpleFFrLD4hG7JR
I9i94luqBH1WdY3uAA+c/wgwRCq56Oz2IhnANRtuyYsoD3SMtZWqJ5vtcQ6skKIq
nwX2QzmAz4zyHEz2BFTMBaxHNw/7yfmIRtGYWTXCYnd5m79qP2YQiqJBpp9bzUnD
oYn0nx48xHH1K9gJeRYlU8IFIRl1MNzWZslvPiiI8OMDW1byco3KwH9PsdiRcMpc
Qlj2ppr8tGBYEfo1kk7XNZzgYBXKvLS995fJpUo88DXJ0Ljpmoi+rV4MrOuSR1MD
EbsuFMpppYpn6y/m1yfbWUd/HirJDoFlv4fUF+HE1NPxEO4Ylb8fwhsL948Tc1k2
EyND41RjHc+C9Np0gNNfDGzTR7DJYbc9bkx/s+ptAS/ydrT9aV3R8dKC884LQY71
+SOWV/MdSUBeJB+yFQbaCMQlnr1pgDcU2HBKjdlb92nL0m7TvRvjXm2jzrzPiX+x
bDV8XVg1McLNF7VKw7fvYjW53W2fn1DAq0KDbiRrMY0HtPw/OlsLDrajjxbDsQ6V
zmgojA59x2N+eSbNcJFHsC7C8fAcZM/GuZ0+Y+pqPLkUeENmhAsdDqI1ZTzr+l5C
1cIrbHtYbx6tcfP4a5XXiD8MYJXtazO7pjuyAEiFvoDUClamowvjuhvSbaAUE7QL
mfn6juP4KTxA4EimPLAjHRfR6Eosgi+D4/gF/bf/o2mX9aJmQ0RPTANAfU8TS67h
yqi7RQbluBPNq4wFUfF87eL1ZhsGNflRQvbd8K/b8W6xMO3qZGQ4tF0JdqUU4crY
yJecBGKaZ20RYEO9l734cMJnaOvDBDr7KMHhi/r0G+/jCI6KNnz3fY4VgVrW6B50
XQiR3dUREIeS35t0EhtORyvPWE5T3lUwzpZ1DlhvNhbOwqpl2Bayn1FATVy/mbLt
w80OKKIOWEGk+dpwYaJDG4jqh1+/2deU14f0So9ShfBXn0PzM2/WnYsJn8nBSMx9
DDuUwTLPA9bYE4qOan8qjU4e9QdsCn91Fqph0JwLyZH2qMKndSnZv+8dzkTaIAyx
Na+pBjfMi1ufhHqSq/5ZHvxa3cy1jL3KWCZ+dqerRVJvj2iVrCA82TKzwDv434VS
BHu4OBhutLAHgir59VfMLncm+7Rx5MdVGS05VI48CbgusnANNwfXDRbomSYL3rWN
xlfiGMEA7vEAqij93pAZpMDlmzwikAVA009SaxuvI0P8cLZc9gDp3xU2qLlfBdi6
si6RB6ITYDkjAeETBRFMcgKrf5lyJL41NlW8ORAk9F9Q6YHEBa0K7uS5gfD+KvxH
ib5vWbZj+HQS5dKJeeRC/5Mr9wAzzbCT+2qZKWbiRnj14EBZlik3diaOnYcucO03
8dZWT2LqwO94rh5AL4TVvtl7sNZCNj/3LRuSmZO2HUFJTaWbD2RBWGInUQtZ+3NV
TsepB+gKJEWnXdWe6OiYjulWjINaMHKsI6/jILQEXna/d0T5AtTMwy12UNrG+hxh
YBbV1V2uy7T4LCYPzdwg/qhwt+2od9RMiQAmt0+nVHTipCreeTBKpLmwbwDYzqN/
645BJMKx4wBDC5qm0eiyRdl7TKTKGUjbh9v5QonlBQFHs2yhRnqBOvjgep1ULGq7
3huGd5T64f0qByAC9O6lr+g+tDUrR3MdqfN4xSapQwiVtKpnPzw+7h6Ughsnoqy/
Fy3hyZnJsDjw9k2+UAMhm4ESVk7NkFiYWVflSSfUUuGQTvrnmxNUojQssxXX/QvW
AOcbyp5xtD/eyuxGoTv4S+H/ST35WAy3lH/1TIH587Fpm603M8YeI9S5vYtCO5Nl
Ap/LQHl7oKlWpQ12i/Hq/22S9H/k+bTTwuIXsgaN80st23xb2WsB+JliN0BAdvjW
xYCKmFFlu1hkk5I8fiE8TltcVxjR8GQeLZhJGmJtQtB8bljmgsTRjr63mguJm6Tu
DmHEOo1bXcII6RfYmHB2awrwx2VydLrmTMX/kExJyqQTg0BIO5BLAs0h98aWsXhy
CIq9uo2IPYdX9Q6M3Y1bxw6+/8MIAyt0TYimVaHYe+WvjRNpkpnjrTn9UxCn+Wys
HGlpyLRstFiPuAmxbYNGh9/YMH8p5x1b7o1GRdMMysq+IcQMGQeMGhK9H6jBE9WI
IxWMkmyqB8iYpeopzEoURdSH5CAVUd0zUoWTElIIZzAvydAxKh4tMmCdJSQtp+Oa
M+zX/wghB5sdQ0bCB0XqItwNI/zTp9iWrHpHTEGtsvE644gksLErykKLXEwwRbYM
OKiEmgucQdWEBU2Z/6Q87Aqjv6txLnRHDma2zFgIDr6UJ2ax6orpt1HpPRWl/BTj
y5u7cyHOz6p50FJ6KxMyN6GWcOz+mEbu5odETNMt/tICmEDPLUg82LWJEzn0owPb
NgCN59l+e8P9bdQjx92f5lvh/bg196zWIFl2y48JG/I1Uf4iUzK0tvAI1FC1MU4U
JJ4YPB1wW+KyMVro3M7BPIs4Yx/O//lBv3xwUgcupArnN/oX+nvSUMpJMtJAUT3U
4uMt08J29/n7BxCnApfEHhwWH5G0ymaiZEPCg8jZUnstLAnyu5buw+bsIF2onuQl
kmTr9u74hOmUjm4dpXQgj/WA21FE3l8s2y/22UihBy4HzqD03IHRKJHBeV2HVOrT
o5KGC5iWG8NyRNV32zk3O9JhPOt9idR/JHSmw1SCkJpdbHb+2hxJ+SPCZOcfX1vx
8vjRV7CyBnmUBTHqpolX8wl8chu5Oo7N8YZ6e5LeMW+JGXTSktHt/1CvweuweVQW
5xGT7IVa919uCN3ck2l/ndzoWCX9hOnT1eAGPogNapFU4mthProcShoooOpSzsxF
Kuo4qAti6b1KLAsmvUpc4LFK2NYGPb7urz2/8oaMKFrKUt/5iT94QI/lft3EWsGW
fhblIiZONRdtHiGYDm584z2oq/z65LoUEo23xvASpDyvQPltcQglDLaYCAaeG7XL
sokFlghlvcsNtORtZXOA539Yzp83ByPgAez674ZjqC+S+A/JLvjNhqrRnNvqjb0R
klUnEJzRw+t4e82H4AH/LFpeOdjNzoYdLyhcVIQGV3iuJTqW4Vik/l75pth9VyuP
ADbIMnLE7I/7OTn2Qp3LgFFHmGrEBy2eDAC71L7RHdahlZNGxKx8gQKZZNy8IfdJ
WGGXe3WaJE3xZnGAMGfXwF5triwWVQfB9nPw+3aHfmvW+tHE61HLdx7+5ltsLIXW
XMPIm2TFzHGs4uzmexi6hwiY7l18odFqmO6Mxw6r985o0qrHwIFqFjTJp5SluxwN
7qfdv9c2jszYLNM0UI2qHtk8FotA6arPhsk7TLWdb8jwc3eN45RQ70ABQAU4S+er
jTOwD6S/AtDLbngKx0F5pfPe1inlrmDSVrXzSsANpExtBAAhYzrx26zjk05Brf6h
5VDateqso4abiRtMyckvEQM1PQprBqA6DiTRDB46Jp31BQPj+XG54P+LTe14Ac8r
CSH3KCpgXlusLtEj5CIbYEpwBquUDSKGPREZRJou09/TDypKdAVgiszqUXanb7GI
XrvWlTV1+JsMU0CJiy2OqVrDMP/1+047TuDh3u5KEtR6epmC909BMbm0wjOtN132
MJ3xBNc8gG6b39NchYaHlIJUcK+5rmWxRhDjNMfUUZpJ73gLhNo4cJNIdUIa6MOz
SKlnqu1Fxwspr98NWaMhsdKXJMYmH3zfA2bb7CEdzDyNtAKuoB/IohePnVbzT/+n
gFoYO7kTLEMpsOaKXaVN7Gb3liUc2lDy5dC4Dyl0CsEdmhe5CZLWLK9axJTsl/uB
IwotWk1mgcJCVh5+PRGDnRzlxfgpfitW/RNgO6yy1eUg0R5ze5fuNLsSn1OQ2yiH
2sXVjrmNWIkJlQ2jK9j8BL0+d1+eV73Mzem8w1QA+V2UPVyYUNTEl2DLT8eeoUMn
GXYA57JXkFW9Au2oNlnul3+7wJTsTE2jVwFicN8rHRnqqcKGXPDdVlWHMjUTmfSl
gb+VgII5WG2ItGGGzftQNuu5U2q04GKwPWVBAeEU1Qmf4t1P1/NcY2anik+ha4PC
NMF1wu9r4utA03fN/Uv3aBGN4zfzQM+VJd7Y+K970lBHNxQtUYtSHjzljqrGDpFw
NjduPEWnGj28YSXr9oziFu6rvtuJoobdTcVhAHkeZG6vyjUJa+1Y6Vunh7BvXk5O
SjBIO+OwGryUuMXNYg/XeFNGRpGnu5nO8psKAQorxz59LIJVoQ3g3E/KQBF6Bx+O
hPYDbE3TFVc5uJCxzzZECc7zyPT2L5NcK8DnI+eOxLmGvpfIa6oxn//IOme2j4Po
hb4kN6HsFsCGnGLERyg+aBIcJHyVkvyfkXmen8YAcxNsYhrTWM56cA/ACFvJCJCj
glC5AC2K/ZzCUYZwqXMmAJdoOdhZ9GTD8e8ayjzPi3uygjRhsooe6pN0cGgEjFGs
FMcFU3Srxr7QCsAhQndJG/gOrHWOrDtlKtQsuGLCuOVQuCep63layij2Oarczln+
pr3SLVLEgPBK+hQvFXGjnUwT/ynWx/q8SOwIGdfvA7sbjUnxaV45x1q+aS6lLKLn
QQU9wnqLr/y72ukur8DSyNzXGzxV9xrVBDdlIISfqa+cmHN+ebgduX+Hyy4OAv3u
y6jMVEkrOB5CvnSXDgZz218FzpP4x0NR6LluXoG2sCt5XM2aYI+9ZwBaMJw8y5jS
7MrHlgp9m1M6NKOEAVOjhARoWybK8Br7zWbsRlLEwPewTcmSG0AyMe5KSJYHlKMO
TYOAuGTEo/WAlq3ebqeD8MrL5NS7iq39QrVLNLN8MNbDCMHeJmLh16d+cWrENuP9
Gykrb/20jpQiaolJ315rvfhO7D67ZNvTcJpwMP+yDIiw3TSseAA1P67fGvhYjY+s
PEqKG/oi9O6y7ueojguDuXTAk85WQRhyL93X7eu5hE11czNh76lnGavgf7a13Xk2
GKbg5nl//jGsO+699SnWtFxu9e2s1YwzWEXZcLmQxFMXNkjFVIxzWU6UNTbSt49D
nA23diWKt/XAXgYEC5eDCefYpRVpRmKG0ufE1jgdjqwdYqKB69bzwMXxTCRoj7tq
vZppB3H0vz7IUIVtZQRZAwHXQQJ3mGNRmbirpY8NWCuBChqBPwl04We09/D+BYJx
LsQ912u/PS3VV9O6xffNXb1nb6kiWN7fWSHxIuvd49XU9vB5n43AQPuNzrcq08fr
exdXeTKiIIYasecxAMjbdEAExU3buXXm1NWipJYHoYJmT/eWVoTcFhoxfyqi8Qj1
aqAAFJJScoM4BizCh0ijRop3DTXHhy+02Sk7jCsWl54dEtnacoKCrIu15udfr/vd
VSvlDZeImby1O0jhh5s/TIU+j1JwlcoazwHW4F4f5yawdRRu1j8Pp9Rg6rz7VqwA
WjPAB9VKN/rPUrgQblzjUNiGT+YQn52pdTAgCFlWlqyKb6iXWGnrhMfWZOwyHXpm
7wS0xJW45bSJuCnmUM3RMz55R5eHy6dFNgx0J/k8qJ1ezGd2jAFdaNmDl26mrfuD
7JIYWJRE9sxP+Ltn/H85cO0X5Mi6HhdzLLp46thO01XlCTpGv2qR5jhTnB8vd1C3
fAXLMRwQjthuL3q20L4QXUlwGg3gTOpHG3B5jjFH245/tlOOfX2ZWzvz3Bl6AatM
bpAVBJubB4PYDw+yUaHV9PSwBU3ySjOC3Y77x+wN0rFR0S8s7Dp4e+Vfndqz+iyk
4RRF23PUaz+GIkvcfcPuHmrk/PHlp0qrA2RK+OptA44l9+MflAnVTSkTOWL2R8S2
hEKBSqyijojqN0yd5SLLDls6JAePpxLNcxdCzGBmTiYzxZjv+MdcNEoMdM5u/rdC
7Kt/in8PjAunV3yTn+ExyqJxXIMl59JDz0xcdQuohFttssFmkCoCxPbyuvS5X3Dt
y1NNbnDjFtjuPUpN52bWL68F/Uo1JgSE5VZ8AQBh/zykevQdnBG4JL2qEK7ol+/3
dAlUzlGBPPHvLHEq+zbqEMWZ8t9u59PXd2xm5vb3J/9yqIvxSt3rWA+IaXxoF18Q
VRkmhT5q5nVaUz9aDlqmeNI20LXIa32miNxHhXAeSCpLtdTfbDwpoXc6Cl8CdxAU
XgKkc3pt5USDmHo2QOcAwdWU4H9ZSSKPz4pkXk9O8mvXioBOWCTpriCzYpVu3USj
7Sn7WOuS5f98gURmSTpl7K9vjNSzweeCOUv9qS4sapE9eR2SbCR7Z0CPzVP/y5hl
7RuWmCpBQdIH+Xt2ZD0VMxxTP1BeVfjQzhdDkoQm0FEZuajGHTIuk980xWuD20MQ
1hhYzizw+TjjR9rnr3M4h+PIFKIswbpRM5gs3YmalLpPmX6vZ9OQLQFeB2T1YTX2
WPRj0gRuSMqUUgL7lGoccfqkakMGZLscq34DuEHCIpJYqzt2xlPkISneHW690JLq
NtsIcwPG7Vuqb5exeEUZ9AmhzK6DoPytwZjWceQaSJ4+bxLc5yk5icyKJVGjDjQf
kloyxlj8g/JCVgdrXDZ1dd3nP/QTwFFuLff2z8pMygKXEU3v62w5XZIsseFpT0A4
ZPPw+yqYhGJPlCJ41Bf/sc1pY3Sab68ZGepllT/wHmIAoNZRKoPk3aHhYW1J8aBN
og6iLNd+M0wPZOJSQTZ9XWAaNpLdE/FBzLYUbERsmCsC5esNEKOIHlTcI/LB0pOZ
qRNksU8kwCkT00+Y8RFxHvx1SEwiDK/3zd8ZhVe+6HHFmUDrl7/kJ9WwK1PvfiNB
Yg9uC72MXc3r26gHZKCJrz05spytZHpLzcYGp4h3oFzZ4KTko8IzfA7L6iju6++T
DhzRBaL/eT0ROsQYlglD+B9gmHVqed8IearlIpXFvp4O3FFukayuCBvRtFXUfduw
xhQpesgKbageF7HBUrkEQvOi6z3e/yBg3SMAB3as2pgUw9gt9UhBfAYMpL6RuqYx
SYI1gcn9tvpD4EuzfwycJStJfCUi7YVLCoxZbo63rhMnW1o+vyPKP9mMwBapmUUY
wkZeHflifcDAup67z7cd+muCYcigBTSHFkRRBL/RHkBgiJxh7WzbTVZUFmUxgNk2
N1WHn4K+VFP5sCSKd/MP5O6Z+TVVwMhDYtpdJPdseD5qNk2vFbYfu54txcHrTcTK
AdlFs8ty3opHZvGnZBeYAsvbjkMTu8xWPss+fCPiJbMoHvOQ8gGEZ5ZzApVB0gG7
uWPbpSd/k5B4oLMGYiJ4XduezdO6ft033KFmaXgDV88Oen29lqUCIaT9jA6BeECm
/Kbj7P0sihd/jlbn1pm5IeNtdlJQR+R961rVWs4+7ATLtkwSckSbM9lBIQkx/Tzk
YyRp9H9uksXnmqlBa1dhgNq+F4M5xVOPLj3oqOhv0oefX5YvsOl2cg8st96IGuH/
nAWu4WE+9a3WTni6WeHyENK+gpQcb6egNQCqlCTW5v3CqPbMcw4+ICmqVALRiLEa
EXr8OqngcoL/ITl3z49/N+l0mg/3Y+0SuZJ52JT767L3tkmqgBo3FBWMxAKpswwC
I2izW0yQBqXp5FCk3gfnneLbD9/pw3NQ9GL0kGIFKQ+dp047DXrihBnahFX15BAQ
mdeglgVY7+Zhyx/T/f99lrJZ7F59gQbDj1PpEe9fzUB6a1w2de9rBKMPNly9OrKj
zndwkI9flajexK7bTj7+mRUSkXexHyxl5vAfVFpHWepsA33uBLTGZMFLv2ICldJJ
7nrKYtcvpItLMRQoJd7wKJqwQnPnBp1R81fVBVMFyxCNqikYBGiBzC316pS/DTvm
+MSjVlAlqxyEyB0qckk6dkoFiIstYxDnRqbVFewWZMBGwoSBskfrmjO7LOoiNO6r
dRUe+ilMVO0vO5U87gzL+tV/SN5SmL3GdEX5X/DPH8dksOTcNGSq1A5n1b/yTQ5H
2YK2Xqw1DT+4utU+vaFAD1r6OT++kJGG5jw1gHbnOsxPGxLyeIQnotcVvdopn26r
cp8wqTBZOCcbdJyQg0WzcDw+UKRMxEKR3z5MqnFMrN1/2yKL4L0mNfMIrymPr2Vc
mBmBDMuz3cok2BJfDTBwJSk2WukYFfq5ROX7v5WXVr75rQ+HJFKp42WRI1aLqoXB
KLu9RVu05ytblW8pZ5wY0PtPQNclDUhflP1PqQExZ6t2m/IgLCEe7bHuOnNuQAXG
PsWjEm8Bs/FpuG7/kFJ47yYp8fvHdMxtka2hPIAjRxj/T3WCKsD0LuwXsljROpoC
Uwbn9e64Gfc3uCmfx0C231lNQrOLebljpVAHSy9HG2VCkSRe7cQdt8uahYZX1vse
oCOssB0mCe1pq68kIXq0vbyN5mWcxvylWsjiB0wTpSs97KtVf1g5OTG2fefy6X4u
JPK21qcyV7bwwf7j4wpThapdcS+eJpZa8jQGD2NEml+CXJrluPG1dB66v7yBfNVv
I1DDxuaJmG+dGTas6UzLU8gOhYOB7gtegETYHueYQivXnKHfZs+9Jq89Hs00hW37
ZzcZLAdxPfQWyVb7KqAw8hR1oKXykv8lkwf4CIdcmkqhz8M78RFKZGtY1j87Gg9p
VvuUbhHQURXaJb5FYONIELWhP+L+cMyjbzMb05GXBjf2JTS+WKs3NsWEdjNXaHUT
rfFZPeQG0cbqi9BLhpk4BX8twyN5PTrdsWjLxDE8qbqRDBmv8/sRC1KgEQa+oXYA
4g7XE0raSWVZXfY0wUTc5U2vSYjcy2/yjNBSjNIdlJJ1Sz/vnYTGe3zMcHs6QbZ4
Y4HIhMgree+Vq53eXCixjlIupJ1G/AE+o3Whl44K6rv6chid4YEg0Nn4PVFx0SWM
Ri1EtVhSOKxFZLr107lVkKz5O7jbZLFUnHiXys+xX8NYLVQJ9RScsTyylVFVVBFn
skVufRSnJ/7M5VBRjL+Fbi5XntHeRVB92ad7esO/hNCRgEDbMvK3Ex3EPUtoIdxL
znUB5Se3Gg0Oe1mrESyywl8lO4w0u5QKIfyxab/bFO7xdKHznEb7Abelems2d2G4
IMm9n13Kk+xTFioX305jGYkLC+3cJGIhicLXh0fG0K/hFvZgfdDaZVLzUes/3EAe
wj5UpIaD2TB5d3VDehphI9CxxXzlQWrD1/dUJZr2P+gdUf7PXwE2FtqcKu8fNGxZ
cXnBvfEkgdC8Wu2RdoMsEQqF8Tpty3dr3u8Q+MWkTSlPIVkVw3kedXvw76A32oSU
SNH2jhB1nOMU7NX0qWPdrs4+17ISrnC2NfqPKoiEkfGlDidzVlDz0oSGg86GYDKI
9Dga5P/NS+ZP6xgm8jFlx1AW2nMpGFD6chpsBbRRTb6YZfIxdLYvtGkMJV6rcw5m
Nfd1k4ZGLPBXyY3LIOM+Udemr5oEl7ys8ahMTLpvlpG4lYa5W1XBzcBKbP9jgWi5
wZFjHX5Cjlv432kB7i8tF+3mvpxAAkH/Q1jfH20x0D/yG3YfKC3S5Fh56V3yKeXX
5TuOTOlrfDLzwa6UG352VA0E51kXLOtr7AgEMDZ/QsRiD6a9e+Xkck6CMCyp/iDI
yiWwPLOnARvaMA6QP+vO++T5p0qwfXlu3aagJs7jRODSRsQKUIzwVxKu4kqXaU/R
WJY0D+W1bDSUIGHD/l7l2NzYG4vN1BvC05YZX5Try+dNvXYVkgRLd8LwlVVxzY8u
wyeGZnqDgIa+q1oIc7X6d34ABmjAeuxJsHbXtsnJIwtVZAE0zFamkEi8HB31jN4q
HL2adAMUvP8UszlmtLGLOQ/RRAtbW+d7MURlB53NxkZRyxjugr9jSpznHAOUOegI
s8/Dx9Z3ShjPRVHMcKfcAGjS/PW6V9a6ttsaVS+QTavzBqKccx+7sPMKhw6DV7SQ
Jf7AZgMYkNHVymhT9AVDNo5AAtuyRQIEH+v96vE8aur1EXaVQOlS5ktu0lHTRLRs
WSFIEH5xH1/n0Uzovuu6G4oPndohOQM/sEEd5wYlK8AHD84Zx9Nv59Pq8fGMCecO
p+PqEpAORa7n88moHmpCtKLXIMIUdOhQhNEgwzFmWtchmNlYDkd9fo0OsqCavBaA
UVBUzaBjXCO61/tvZ2wMss4N/FE9iZelIaAnbQevGNKT65WE4yJz8YJZODz5R53P
IgtNlLS1bpx7d7dqDuJ5JVrdHDy7TQTgyg+7byfQs/yUl5PqKUAsDF6QdTIx8+Pq
u4A057RSLvYPFyaAUFid3njrAzc68giV3OzWcs0tcBwMBQwE4iB/qlicdBAdJqZr
CI30xQLwj2B8NFJAu7BeTMHfHOsCLAddbiY4fnsVXfiZ0kYtIk9/CcwlIxTbDV7j
ashijJ4npdVtkZ9CVn1x0zHSqmSNi8ncJigxkotHgG1J0ETneDGXipGL0LeA7Rqo
ZiOXFO2bczxy/qKfrHqY5LqxI56CVLpP7Wnq40+codO8ToAJNnkJOrK2kS3Adfo4
owvPy+yPga6kJcGDkl+9FwD1BXXOcN2Nfnin2OdVGG1scDf7TPfzR11oGdjREfso
ax9beaYNF7v5VkA3OONbjtptlQfeVj4/lk8KORDHkx3UbNbi8qTS6AJU8opFeMrg
cIUoTXkdkNYvk3BFusCI51c851oTacbWJqYgK48csAgEbInxn+Gm/vZSlTUFoYUd
DPam3I05Tmi9BUxt6vG+Mw8XgHmL8r2xVS/AqsI+VAZNw2qk0HWwoFILhvToVkSq
zo61yOAgh6pwlQPHyZqcd9m0K8CJr7DSI78PguWwIsO3KeY+pGyl6jx4hce4tKUM
xL5nUJNWtuu/wbzaQXkn87SmsK6K5NyoBA1L2QxAZ0xi6tBBfHgdjdApA5uJlT0/
QiAaXh6KYvi4440qjQ5fSUWppLvxav80mYzhtnPBMWLtK0xUsklFNAV7BxEJfUjF
NxeerbcDxcmwlaSpPeUO4b79+JCG6XvhaZXJlnackOadABmE4IpF+eH9xnsajOs1
/F6L2dmxRSYpliZFH+yt8O2CcaqI29tCK5K3QHJYBEsJwkdO7chWDpUZh1/Tmj1c
mdfQ5gBiQzXqhN4MbshSV4Ofp8bFFbgRwFa03nDw+FDk0WOfmuslTka3j2I9LLus
lp9hcHAubMIpxoBKjjjLDnKhzippQMdtCFWQWsPmUX79mL3KhsfU5dYF3JHzYVNe
YK5U6G4CfDOAGJ8bjc1bMW8lihHqU1Hu22dbcMVaRxIrbOjoeN0wN9h6xiRVi1Gp
CkSs31sap/5Wi01tDq8c/75D196a9cgxZRYGmE+ixgfFvs1UjjK5jp8f8H2+RauN
k5zr34OSALILUw3nRTwaLl3dugFcz28l15bTZwF3taUns/PNHUHGGBuk7HrxdvnV
u66diBfbrRFJR6XY1Rz35/GmjrXDO0NJERuD6XArBcThHynjpO0NiGmnCyQDCUHz
ogrVW6XHelc11ujtbxuoexi/whvhqxbSEGs3wbhS/bPDAP7ZRI6J2wKl57dp4Q0B
U5szGwStXNxpe58r3f0a+XzNcWLk72pQLU8cEUH5s+BEjEVlHidYwvESdfSq6mVb
+39jgzF26KPMpOVZFP7z9nKaS+vemNggSKbSSuwgwbO28JVlwxtxCZJEMigcA/6L
YlRdYaSNaDz54Glt+go99KJQ96jmDkhmojo7VkM5dIbAtsrfBziUjmUjD6LtCVcV
76EZgX8gIiMliFTgWKeG4D/sQOCyUKYoRrY/l5Zy+j1U4pXzHOajQspElv1Dvqvk
iy38i2trIXtKzKxblgZ+SAkxLnGjWavt4Esgtq4wUUGmBkWiJS5+9K1DrsV8d8ip
2Ks83aO8JnTs1ThUGBVdAvI4lERpe3XPgZpeZfLRUwfBo5dwN3exTC1NZRYJPw/7
SthDTmL2Qhclwgq6L3btxuSZdpt9JJLkDv0/Y9P/i/RFvOMbVtx8beLo54mFOw31
PBTDJVwqtsCP7yiSaff2EZmtcggDbLYUiuktiy9NlARtHoCRcrMWqZv32WN2flx6
QThUSp7DjtjGmZXavJ3P60dk4osq/qRL0jDr4fTkUGT/4s0k6EF18GdXxH9sh+HA
peLsBokUpqywx/aHnWd6t79FjX/xMvPl3P4oD86nXHV3EZRj0amRU+BESk7Jakr6
XvEMUljqORXzdoPzEXkIlx5MpcOOKch5Zd6nY6X6Lwz/0/ZDvnCWxO+L248xw9+Z
UkaTnQbDfaFrOIg5nr1sGfqNJrNQ6IXXeGzOslOApjoP8rBkwIhJ3/4POeKZ/gCt
hqbZcUi3if4cMTwula0019IAdV6dVGe0oObAGa2cOV0mqMrww/gX9x2moqSzCgAh
Ia4kmxbeudbxxWJJnChRwsJyzueEA2SKbiu+9PDgJWIJzKw8mkoNUDN3TdTOCqDM
5+Z4gPQ43ARW/FbMj0jlMlBp+96Y8O3J7WSeUXK1pfvndFsWtlblNIiXqhDxkBmX
TB43efXWoPgj0WHoGbSf7fQUOc04DL87bWsQGVWw9ZRkvsnrN4XNhxu7/epsjBAM
WN5LbMTp45zSMqC7kD/y0uhU2F6k8zv9qVQEvjFzrjbSH/aDMdRbaoMEbsSmlW1J
1jBNogHeJ990dMRP84bL/WCWoWu6HB4RAOnyKux/qRPAK0vzKjpujnGLCXLdd0J5
Kiy0QpswIw/TxslkO8M1JgIzkE1tMbAqDmCU7wYdy0DpX3357v/0eM7xU52RLlsH
OIlqdAEo0t/REOYkEmftqQEPNW5QyMJ1oZDOxHuAi3+EM08XBBfN5xFT6X/Ob8b2
Lr1lQwtk189TqTTOj+WUVFyszIX/zcLfnH/ayCXGohyTLcyoCIf25122QFLGn50D
yTnc/bHKWTH7J/fg3ONlK8i9G6ubwXofb7heruxlmv5Tkbl5mTyVDbEhKAKdQcaV
bszjWAACgpIZE6F6al+lcNfD9vXfUI4vb/iW2YLWdEJfEcSesQ9fnV7Evrbl0lNR
3WWVdpXIdTeV+bRD7g6p0zrYMgxfQr7+11CZ3BcoNeFkEdOBG5TUQr0TDxEVPoYr
qP3xlubyRYVOoDjy4OX2o3bWq0d9dUuGDeQBckbOlYUzJI9Luty2CYzSOBNPKoRN
3lNvJ6M9es+FTSjYlMLUmM5Yz7sWuUlN9hzuHefmHgKAm2lOx3F2w45z6fjxsky+
INFrTVSzFcfBnQaxuFT6fxPMd+qHCEXGoJmUYd8z8fRkS8YxA+XIG5mOLMPDEuoL
NV7X6qJHjUH/4P8TnGeIXEiuUG8N417Kgvjm9fPm+/8jMFwslhYAkyFBzLga6c6e
jos4IhIROj/pbEKDSK4jdcgdGorac0hrc0EZ7J6PZk4X0vgk9ifwu+bECjTQmqbR
j+EqhCcJWHlNn7DiOG8duMamolAn6TGpJHpBstwHOfpqjonTRHW780pPNhOLg7sM
7oNQ7XUhgUJcqX2VvWwqJ0tiwQtnH4Jh4/PsttadAORz9OUKqb7MO4Tuw20zXIDZ
Z5tiMLw8TftBegh/f/z6BbJztcAyntsLdaSdcmPAx9wm4KQVwKE0yds5tF2UhD8+
DEXL0f7wL/NKFZW9v6lbd5PPMSvgjrb1vm+8wIglsNkMn4zafGk5vF0bT7RCg1/R
ejDr+2sB/67hp2WH1bNtVQHbytnNZlvasn7VFym3pNTISpC2vs49vcyprp+bLYNU
b58ag+oGzOsdYBGVR1cmrzoAwOV4AeIDfXAmtHYfVwuzBLsUXfOYymznbD0yRKKh
Jd3TussUG4ApiS0c9D9VOhI+9oI7gmYTiqtY6dzN6K8wi+HdUDWdQc1/uf+Sl0PZ
hHKtfg55+AC7Jjdhycp47edarMv8Yf0oTjJaaZ/UWH8SInkdMoHwobraA5kIUFR4
WDO5F2biVEjxXdyHM5AeO6aPfND4964r2gAGpOnZ0f8D35c9d4N2l6eLkbwc2Muq
IDhqldW6pWu4PDUv3+TT8FalQWu5hnfU/i31se2nrPmnJur5eatJOSPLvh0oUvO9
syBr7mdjVAagbZvvOmczhTT3oU4eC7fb31M1PYFSowRg3Q1HJbCDTYsdwmcOzBlq
bTzxVTMSOTtRWrqxcVPswzT8B8bn3bBp09w+lwuLRpa/J6lM0ErSPKpdKajhyto4
tJ+uySLHuXlUHGhQq+6Tj3UNrLwbH9CHzRuwsp0RwtmGwAZp9lA/tTY/Kh7ExIKL
FbLOCod5mDiqP6gWDU1nKxbm6/pCfgX9dkYe1R4ANs/t5cwQmpjIIvVV7nL/0mqD
v0LmRq4XK/5Jt7j3k2MCnffBgLAGHlpd3jQXuG86i8nhHHLbqTpOgLoqKnZIZZ8+
7YnaORUaFIayj7DA6ixgwL1OoP96FppnIzUlmjGpcVgGI9biPlc1JERKzHLPyIQE
tc27vVhNfafO69SvuSz18qLmgkemFLY+zL4fRdiyEaT1jcI8DEBcx1C1YEOPzNXn
xP+io2tgKjEi0USHHuLeaFxnOXhrle44+KqX6flZqvSKqfZAzJ4RfcL9R2O6i4ZU
GC6ClmOQnBvEL2bQlpCCZ3UnBJxoBiNASFeldmsFrsTVeAV6i87eZCagSr+jFCrr
WwJrny2jiEaH4bEXu+Yy6TSC/J610THxWd193xh5m/8Zvk8Z8baYvQYhnpP6o9Qa
dXQMTrd57jU84EP9dGd2s1Alc9D4YVi6c9WfCo5AuxhJ/2tkC9Kh0NNfn85bKadR
GrJWl0PwEZisfiTzLuNUdFqdf8UwdySUjbTwGLW4r4dBYEgoROgQQF+jOY9+gF5y
kb2SjclNRWYCjweN+/Dm9gEVpl5ieAbw3iS2uVwtcDULbADWGoocKsECXGvCn+mx
/X1dneqybNazmwWeHhB/ptTX7nl7N6FiuwyV181ggOuGscmZW5H5+rnenEZbZGtm
4mjW5ojE8MuTWR1U+V5Wblj15itj+ENYGCe73AAQc06KUtrhGkryrNwoJCLD0hV6
Rr566BCv8qWzkLFVi560OTHoBqm7/q1xfRY/4fIOqoqGpGFdxeX9WPZaFcro2k1e
2cAm850kGX1qohHDxwCJNZtGzZ6mgZBuhMRtUMXWS0ChT/QD16XvVPOStkliPxY4
nfGTM9/5YQgW7fwssUm64ZpM406B7pw3Qk+1WCNXPj/L1RiZ6KyAQ4u4k9FIC7qx
m6y8DdXXr/KvXaWOTAShaRKCgH8QegsJVeTRrv5Y3AdV2i4ubSsdNpc/Z1GRhEkW
MS3o63WzhFJTV/l1q8L66D78+6LxPqkOozxSwzup8xJjoamXBoJfkDSyH4KYqe0l
J1rzl6BjzjZQ9JGO8ASlMStFO+/77Ff2U3inVtW3A1GY3RkkB3LljkjGxjRA/iKe
IHHceHiTscJndnFFV++utULgfP+7DIGNB4OUapHhMD2QN/Y4tVAN/JIFSRb2p8oh
7AsdsHXaplI6G8SHFW/KjuhNGFnpgWZHHhXblWVMxap2xyge5lMo9NDU7W5TupKi
UM0XMvZnpK9RZfPdfdIgIMsGmRkvqofcOw2q3XEzRS9iJ1SNXx6CP8VGpuWqQ9w8
ZiOcJSQnPuJCGAvPeW3nSJDuvMd9PY8eG8dDSID8RotVtJhCpm6Mz9ZPOxSY81RS
URkyPHh1LADxQXjfj801972cgvKLC38jeDaZceJgp/7FvDQCVWxnZHkjRk3L2FJa
AbOX5+zdJvVgjBhMCfzjtfSoLKYX2BA+9FS8Or9oppv+PYDdmKZkPFeeBNrJNJgs
8dcYMavpNxR/TaPnulHa7Xxb6E9ywTzQBLg9g2FXLy2e32zPla14YSKVOCsBL85T
NN3oVDuyMyeSbEz2XX2d6FNjE/I1S/22TgqWDlv5TXpqdReCZV8RiTILfi9aN/lo
wSvT5oV1w0bd992sC6AfdAazUMTogFJ0TTxDTn463dEp+4lMsdbAtLJB8wWy/ZRd
Tt2toDyl1TInj0+mRQK10qEaEzOzpdydTZQOO9daiLzJslcDS2rtwEvW2DF9rbp9
Gu+lFbm0mW6ZeghVpE8ZDJQrcqgX7Sk//gkpcfGKl/+GzVO5SbyrZ3U3FCfTa2CJ
2OiqwwKqIxyAa30WGWM7BUKCnmcNK+QIZMwjVIAwnW6yBOxGlb7vGC9PiNs0+FwX
t6/KGmaruncDgOtn2caWVCKl/1zHlyIBapFx/qOrIwHdzGn/iH94kODwWiTozqM1
JdJKvrvqEg+WimX0EAs4R/p6t2jSqjz8Wd/pEO58AfIps2MV+Rwa1+0hktWemr9s
bsZmGvElEYMvGqynbINKzJar4h3B0Qcp50LHMdBww6b1yzizzySu5kOfR4BECNoI
MvuHCmN0DGw/vKnxPZNv/XO2uG56kcDbPBnMuLPNGU4eHUtAI60KR0ST9jMPetyg
EOXQsCc0P2TTGqTmtiyb19nKeZ2sAY+C0c+C8NE9wDRq5WbsztVruFYV4ciIEvM2
EAQs3u+H0w8XwmIiq6MkKbR9YDXPgqWpOhPoS77wKqnpR/0lg8fcK6RBWts23nYn
oLghf07F60egcbpEkmuXkkKO34dlcnA7IxXWZFg1SIcN7Hj2HERpDW/jOvUW1eA4
xgN7ZzoxSOxmsj5W0rFCsEVHcA1aITYSlUVIlh9QHkxN6UWplYvyIuUAYFoHFtCc
C72NoK3S9hNYIHtkifL4sU9jLDKE49fv6x7IXo0XNexMUuNFbIn7Hg3A2gsTxH8d
so2VlN/5ftxHB6b9fEcprl+NgS0mfW5kC/zkPnBZghVJfzR+tUOeca+eceEmI59t
R4BwyLKQBG/tjzO7+TupA768pFD0eP94wUHKD8X+OMvUJ6mmGE/Ouam9F1tRsO2z
0hvpCXt5KQCmEt+jxCz8adgUtWxDxPU1RYjccbcY/v2yiOL0oJoyqPGVFNxoR54O
tjMZWWvjL3G+A2uyZyuc0nmv9+ytr5EC1DM4nQtcTEaILBfpEifJt7Yy9WfjyXiJ
BrXwIh8aF4YO7RFhrpo+B72AvrM4JDENIw69PQ2m0EdFFJgRfH3Y684QD/2QvO/I
d2y4w0CNAG5jn5orBG6h9ZjoelD9/Cljt2vgto22KMzAD5rXswKu0lLq8goS3WZl
JI91XnhHUfcLTObevCAJ+vk0/o7B88AW0IQQzvB+GtH1aTLnbd361HoHuY1QeItS
l6c0w5d8nRiexVytPTaOkGvFMuyW6ryco+TsxsfJQ+mgCSj8/Dv/Z7L1SQOWm+6L
UZD2k0X2XrjQ4e8nh35Mm2DeokzxCsTYP2htyr0pVcWPFXsUwRsKM5M4VaI5LIc7
9WypN3+Tb6Rr/2ssQPVIXSwFnNSS9PCg4ewhBke83BTx0J+eK075I+f9CvRpho5V
GepInCt2J4WLdYi++SsmaTOOuCS8bWwJBzYwyYNO0HBO13hsNeKY4g1YK+s8Uxxn
Ksy8LvQYAHtgJsk/4YqV9LIZAHiYs9jcd8YItT44qZX8989P0oVlr2GRDBaQNN9/
mC/ev6+Cs9CWbot4RtdUTRFdhqjsGok4S4IjYXSp+mj/AiAz0t+q4UX2WBK/to8n
6Ms/A3c2pG1D7Zv4m5gIEnTz5bceOtXVLASoowaxpuz9VA3YOTzBSM8m3NBjES1e
fPiV4/pxhrJUtqQ0D+ghSIN4d4gE7K7OorFgD3DzFVXebFgClSWxLoIpjLCU1MJD
Qo0Y5hPRP+qJasWOb1ojYY+mRFQh488hIZ+CwrBilZFSMjLQU6tOfPQq8712z3/O
aNIhr9Z8b8FBdXhMDpBlnF/7WDHEuwmEOSxTJUeStCdQGDX/S5LMX8kC2RHTKETh
N6cDJYd748pGCP8KZ7LJsOlArTorgkjVorwf6Q7A42ofC8jJ+rb+zzJdpF41rCme
OnXSxi6bhrMTy1r/CbrYytagM5GN0VzmQuR4HNcIqNwJzA+dX72EyWs1AjPfVLwg
p8uScqs10GGvsENgsL281kAlrxBkoPECdOtUQq0VoX0mqXQ4td64O0BZ3DC8buBM
SV1z7VRRCbH8zqXlDuEf8dqu5eSP+ga2mgi1lRoLVOXgnpvJhxnZN+JFGqXC7B72
IUK0iuBxdU87yrUzk6hEzH0x9ehACZ5gzp6e4I9vchey74pt8rLpcq34v+ovezcP
trrUdZs5zPZqp9TIAF2rWBpIvRYoXZl8Gsf0EZFJOgr7XmymMWODhlFSdztp3HyC
TNrVhhVY0L8tN8CeihjClEK6ploNNm//Gzbd3pAaxKxccQiXZwKsYDKwhgS6gPwD
xSN7wzt2w/V8e8/7Rcpz6Oj2wN85gGIqkspQq6vzJzx7YYFP5uKHjsbzbGeU4pom
UeqHecekuqDSs0AlLr3naqXppPIJPlt9Q6OkmsimjyKGUyWtrHbUq9xQwmG1BTEB
zJ1xF1FZMI683b9HEZjOjAyAPPh4v05xVbW0Wz/LT9tAopCM0gyw6kiBPHERozLO
tXZyTxGtnn0zJHGf0nfvP/QLQZkwYrgN1d7cubpF0CkHOtxX0otolFgG6JCL2Iy2
S3TfaxOlxifcYxxdwh5CCHYvx2qLH0F/Nq3ywhGxkgeUMvbYVXk4iMuafoASZRcm
aXK3xw1r+6zqmXmeOlXjPQPyT+ncTwDPmHLaoMF3L4f31UiylFRNZqyDtHX9bLp6
+25db2soB8Rbn8go8HKPCkd21aZ+IhsoztBQI7n/MCXphrRIYcIJ4Au+YLUhA6oR
3iqeybSeZsZW+rNEJLgfbNlhNgWO3oirvKflzRS+ubJYRmQQPKLd0+7zJhYZk+e7
r2MT8GhK+EuOA4hSZGtnWkxF79P9Vwwl29kn9nYGyoOS2zti3cJZzJrZ3mWguKJT
QFn+7o/OoVNpNUpZgc+XZbuZ2UcACJbPE5C0P0359wEf/2NmeNW3J8Ri+iJgSmqa
hs1oAosMpYqpodJ9lTWvXHgjX2m/eI7CDQsVx9NodpMPebllBJOmGVg1jEBT+/gH
agCBMNChTRKxTvmFdLA3iMfXF2/QIJVWee2kb/p4xm7rS1HfPqtEP6/eJNTPemim
sC+EvVsn8ax8HOtr1dNvJxhtdAjcXCisGM6yDXDNlOzlqMBxqw7+h0vGF9FQgxjb
9TlSArdCsZdrxgDl1Od/6BHDaMp7j1keNHpygnhKppk41n5Ad6cI1ZgjRgtUIllV
r8dKueTQT8LD5yoJg7f2TuOkFlOd0xYfwAHPZJEiQ4zeY66pZ5NHYO3RUSYQNXPs
EVfVkgu/uoFipgwMcTEjhpexJtYLRp4X0+OCuMDBO5x935MiCT8Km1T1QwEmEQjc
ObdrPygwqXWmbtl/r5eoshVuyvPV+yFNcKDceY3gT07r5M2XsrayWkGgiiTP4ZSH
A4MGZ8QV+kAypqNSMYL22zGg+xzgCwYatWivsQ/HGG/3DpYCUm3WYDGu43tgfh/l
x02F2PtD/GGhR2jv9t4wrPnsT8gmhdg9bgShjME5sGTNF0S85Cv6tj4yMPKreAoh
yaNDEQGis5Oh8cK62y0DTRIB5zcIlHaEVh2/QEkqR2Sq/x+QAQK4EM8t8o36W6L/
LdYU4d5U2lZ6o7Ju8DPerf04X9y+S86HJ3ITulL4Dl1KlMNKNbGSux9mz3LbpA/j
cPMsaDNlJTa2sFJC9YUniEbT0jEowpNzTOHzK2tg4t0jxRE51+/UV24V2keram9t
MZ8K37lYDCnrgPRYGsefNItBO8I4TcwNzkKRCNy+hYPD9vutA/poHIuyPy6aU0jk
H87pTF/9WRYhKiCCzerm0e0appw1vqhaRxWU3sMjR5Q9KjbgpPFOec9uAqqLQ+T/
OVUX3jIc/4av7LwH8qwy0v8RQr9nSDaPHLDe6+rb2xAlMigc0alu4m8kH/InMY+s
5fFTQJ5F/FvmuFOZRpd4vlhBgjwmFis3GBYbaA0CNoTAzJUSvmDVHNrSOPrVLibt
0TzQHuMsZ/Te86J0b9v+bK/7dWwU6ExRvqA31f8Wi55ZAI/NQm6JjI8QE7brNERH
+NDwDqFtxpS6WqfNpzO+QcZAJTnhYkHwIXZofrQ37fjqdW5ncwroPTgqVRlDBm9u
WYfH4hxhgM6MmwmtE+IEq7aZHfeMh8c/v/n5TMhQnC2y6Xrsgx0HgJRR8zQDM11j
VbD7Yr3o8R8cI1B4j3z8s93gkwKs9AGaSvJp5EKZAsXZuEP7wVeHu0ZPGC8mbm1T
4pTyL6JXAfW7a5nCK5mRFm6OoDVmPjyHZFwvHe9FRZb4oxeX5sz6n768AoBEpNQE
QfDav+X491NOYsBBdeKkOx0x44k8lvzgjMpGVF8Tf0djijBjWFt90CcykGwCZMF6
EiODol/Pn/6Rwt99KRqKXmgiNtFRii8ZzzYnaDqZ6j5cpFqph4Ock8Wb3QLJobK8
3ZkXs50VakSx7P+J0KXJJ225sCe5qjGK6xHPElpFKNshRWW6nfddcpjHCFIQLsBk
MsxewutwSLiSkp4ZBRqgvZxNoZ53PaU3NlQiD3xhPgt4OrctuPNSP74RmTnkN+Mc
mI8UJu2sBWG9GBk6e0MvAqoZ/JeZ7X9EtTbBWaKC6C+DBqa68FMSfrAvp3pWHlMe
+zPmzdFfCVLQkpzPO9ButGMtAZYQ5p2n05ujGhR3zlndYAzXV8A0vdH8dmbGookh
fc8jdBLaK/JD+IYgH4996svne+ivAdBndEprPMOXAVpFGPzospcrtFwTFQgYgu1U
pstkOIQxMvCsUjKyi0T6lqDt5vMuY/X5k8phrUjZM5Vbmrny0qV3B2zNHSm8LMnb
EoTzThq1podZr9q/PPsM0MIBF2kvp3LDT9/T8W/DKLfzIdcHwoMCD+lcd/lx6bbV
7Cq+GPBZvnUJaTtrHhljON5v99DZBCnpMrDMAZIlgwGci5Rh0D/QmfZ9nfnM5OXh
ITywiIvUHgF2e8wRARuptxVFBUBSJfYLgfqcwuaib2X4ib5RguaUccUF6tYthXHf
bGwUOjN07YMSCzN2S/Ddtauwvy2H6R8BiHYGypdbi55Z5CzOuoGsYaYm9U5ALDAJ
Y7u79Su8LkwH/RL3PadM9OnbfDNpQWkjGxj3bJDDRW0FpFzRZ9enaQPS7XqrFI8l
sox3g7RjaoNWPoWhmgXhtF/2uIofZ2yB5Tvmf/iFOWIB/YWwJ6pMBcu6X7NuN601
Kk6Gr4a2obiAaOoG6xrqffzuy7xcr8idh3Eq6Ar1Y3/iRkONdnqvBRWMEpByAjsF
hlVDFL32bqY9yhr3PkIiZuBeuzJAOfGVhSRbAXV28RWEZ8p0nYtwSk+IE1REI+B/
cmGGatYUKd1QSJpXWaqvqD6lKjVN7f8oBgSUM3hTJabPk5H+MpXbKy9+aZgF4f/n
kdS7KEyWSu+hLG04i7C5xfKwZ1JD7V0G9jr5948czCapFTLyxOqSszJso1c5wnij
FKavgYMPwAGN/AS0Aqzujl5xApPp8LWYbzMJhwRzPhy6XcZ80enHt1g4u8bnD5fD
Y/EI7VLQvQHmE/VCBpzPDntcnF00iOBBXQmPGhQY0FfLQ01A2080zffaogWShUs9
5MUL+ELtvPomH3kpMcF+mkBd+Y72fxec8hbAZ3tQIBopH/grFR2spoEZuOHf81n5
kT8kGPIBI454JiABt0a0KgcISirsLKefl34WcM+MKfQeR35WmP6bVtG/1iudsYQC
SF63DQcDOpdtRq9pus7L63ZScodnBALrdN/yhhWAo3YLgEeHqhpsCdebVWVNywS2
2f64F6b3+JNi4AQk03Mz6HhCoGauunJOCcg0H28XKlK3j7+y4IYI+fvVIlgpfWTd
5KpcT4LR6S+ZCxi6JnnwitlAluXwsTLkc1GBjVKSGvDf8jNQa/b5gfg9DjpA0t6g
1gd4zxtjmFXbnTLiClfCuAxWQZgbbkRIkcnLlFp0FEU9i9jdbfQi2+iWHw/S1LmS
lmQ6LXoOrF9FZf1ExOl3SX0a4RaJCcF0QMUPJmTUs3J0gzF0tuCahhkX9qhPpMbq
+e7E1hJgXSw+Ryd+54Og6GYKxg47CQI9paaIZxXzty2zQXTc1fcXy8AJDrt6CIbx
CyFgbPNdZq4lvKMI9Grfled/QBv49GTfEN3+i18ScqRwiiOepXPfbOfc7LHKusG1
LQAERPEuy3Rwhq6SAiXi+x7xjLUhM+cAyYbMiYlM6A/5BP2jOKUDXLORl4x2Dg8j
aOZvGTFkTeolth/Ipd31zjq4XbnY0KsdMwezo9+1EH43QbEof1wve03LpaFehqfh
Doo4P/+9JPfd2ufRNf26HynGBapyQMZsxoYdsmCJeyOHqcjMRf39K5pxGmajDIpt
QbQDRKvrI5OMftNbq9Ir7Yh130aEnQz8Zfgydaxd2PpSvzP4fjBXvU+5EEfHLFJu
eky8NJzcfj6l8d+bxcpnN5tyv/hOBAo3O3Qz8vb9NMmhjR226ho8qgSJ804JuRxm
nwOAOTHzn/0RaJtp9jfffiV86UdM0o8d2b2ufEJTrwhmhVd2X52mcacClJ7CgpE0
7Pmox6T4jvxY3DzDihTbDdOAPLfRG4j56dP5AVFT8uAqhO1pzXY+6DskL1MxaMm6
xeocBFqqsjBrs5GCG/BqH/IDpdnlb/sAto/f+3FH0wz1U4hYZBMQJd7S450rzTUJ
tnXliWs11V8TDolVUDCIkSkD3DXYPMsc7LzZW0OqPEt4wjey1iYWRsf3npATPEmD
3ASRevNywSkKgXJ2UJ3wnFAzWLXATe9vYjCsb7ZcstDyDv2O54TQ8JC2iwPIwakf
m4sX9KgaZGcV2cxxdx0TOiO2nAbEY3bQ9OLpzXLAPo3o58AB2+L9MHP3KIo38UP/
u5cs626nzcYPMinJMHtWROAYWULvGVIC56ERiM/d+wbjGXDHEK2wL+5MRnSeWUyv
jX8gWccL5ONT2btvGZncheXqy5FY7UpZGDaqURf2xbyWINTQQqYfpO4P4PXZB63i
lSnvNCpMAqHH1iqB7RaL+U7baxuP/0TfdaUSU+ZJYzYmLFFpNMxhiSM/P83ka3dj
hL+CJXYknWBNfTsqzRmCF7ubth7Ugv5hDpJBN/Vvux90MOC6mpuz29O1CLXh3jax
vUBsm8jfWdJydq5+KBeDKh2VSW/OX2DN1MV+RAQDvvcA4PpzbVDlbtGRS7bra7VU
UpXvR70abvKYOqJ0970m28XG8pll6a/cQuavs94N2pNEKrEZYvD/ufhRUE4paSHD
UaAslf6LFKYvvND4bHVFKDAZEF3BEdHJ9L66E0fquSppQk4jbnHF4QcF03d1yJdC
XPLP0SbX6Z0VhXjjC4HnIPxjEpc4jzHozNsEn0nnG0rYU+jmhGf2JO3R3KkWAlxX
HfHn09WmOZoB+IeOTFd0YAoWx4F9Nr2uDI98EOSmwauqrzaSoCXI9RcElTELTAdo
fwNidrBK73qBOoGuwI87Hdx6FTRGcpQQEJNs+lzvUYd7k+awA+G++QHwFbTmeZqi
91gIMTahKR+kfwvr32w8How5CuQ3OEsA4aOTwH8RU/HGfD+bINr9KpKG0AO4pFau
CnFla9nxk2SUui1NpUXTIUxulVrF6Dd8wULwT7+iomTewv2sgG7iuBO//2c5vQiN
RD2Ng6B0FAes8wmM1cNstn62EV8IbiyQY5VHuCidotD/wIrLbPrsvLqbZeskzptK
odz3D826h0GVZShF3efJMrZd8Lw8pSA5dFcF8uHJOubwidvCYewiesd2tyGln1mL
QutHmYvkbbdC2src3qZAlHVuguvDj7P7F9navRvoiqNtr11xKeCK6UXXAl8lDhgx
g7ewKX3hux253lo/LMVkX2M8MymFMmHbsWkNDvlZdnjCl++eqwaY699Y4mirlea2
LuRaQUAKZj6E5Ge4I6QQozpvHeSQcFt5vDrGZirbvK1SszpS4so/grAo8pUsKOPn
gZZ9Sj2DOuKmbMzsBQWmdyHgF9Acrsj7AYVkKYa1st/XZTyU2DXGCmat1XansYod
V6xLkH71COcp6nS4QwU/LJ5KTAcmjp0sJjMNXkwK0TbuZ3VEr82JuzLiqrHHOKtN
pB+6rxEZsS8AMCAZz+q7z3Kzh5bC6y56q3VI6rN9nUmsBHDd7Xtf8WFQTEdLTxqk
5zC8ck5sokg0jSksYhxnMtkVivBqYV+bJo8Adr35MykQS4P2/CLAZqaV3CTstznj
0zkPobDqeJCv1vhSey2WC7orA6R3jZBCFL1vr2YXB2Qu5fRNUqd2xGlSMjEr7dm0
9wLbaBt46MW+tpXnVRMk/nEizS2ZrJb790QCynzsokiw2ze1j1GuPrf91kknJGlD
4V8NNMDKNmFWl5bxjazsZTkjCxtz+BFp64FX+B+5Mg7C7wtq1LSw8SS3rQpffUTp
2BduJPkT8xttRHQbKUX2qJkMAhJhkOY1Qy3o7Dx8GFzVvAfYWPEs0+QQcXyi4k9i
eYFhdYEkL3PVY6R7uRLw5+XluWYeWOzsrGIZwbsrW9kgOMJ3f3vw9xlImBqf2XCa
codC6QQ8mRek/WcrKr8oyffKJSZBd7SyUeRbKzrlZoIk7BD9NuHXFafFFA4vGy5P
4pJIgZqCnww5IzG8gmRV1g6l5OF1E0HcCiXv5j8wgJ8CcBMLouLDo1Lpnz5U03sv
1JzWrJPV0JjNIcByRrNDhSyYrUuWzEGPB2zAOheLAz812UShkWwqfUHUfIGdyjlO
IyekIKBzVwGQBZgn0NivuYNGqlFJrnF3uaYRs91vxitbekX7IonwcGTIfJIxvSij
MGg2GLCizftRxzGuOicQHcfBOagiTOOnOzBazf6Um6FnKRbofo9WFQ6Ij2iATIga
716ErVPJ92V0+ALWNsfoBzXgiW01T3nWt58xyMwB9drcSKjC8rD/ZPFFNUcEifFS
WCn/rtVIjnXFw0a2LEkmM+c96OS8TlJLXQT/DA5JEx7ZEMt1Flo6Jh5TJ2DApit3
1fXNh3/XhdTK264fG6w6Lo6OLgTKn211bTAJJ48iNMrDm3Tgg5yfu4ZS4K8TWOiC
vXOMVpeGAKKNjjV57560qIpP2CehPKwGT1ejzujyufMvaHlMbnoodTYmySuzvn1o
M8uqIwV+bJmmqJhaTRAhMDmEIq2dduXMzt3NMfueDuqiZIHfOBIXqkng49EakhPS
d1P2lNy93PJ+zSmcI3/0l3UURt97V18te7MQpqQ7nkldofcfEf/HZzxu7qG2s5g7
ozoBuR29S9G2nNLWMqAzdwC4OwVmmzEKfG+KQvdutBOSPQVDGrm34VnRrozcPgpN
BgpwwqL3tvS37ZqtzRg1BbuJnpA1yLhVPpXjzIZgKtCHtfokIED1g/syZb2GL5FB
TUShZOr1b1koLiY22U+g+xy1O7BZoIGwlo6zvbj14D6ZBm3H7x1F1VtIrsRgN6S8
ZNwE3D69IpcLdluoZsKJodmBsIfx6Mkjef3N/Dd7sV/skrDLHrUEYzUX479Aw0h0
5YysLzHP/zSPu8gOPw5kUr1YsXYOziR8QnVuWvQtIPwY6jo3teB6aihZxoQU1s2j
r3gq1xLZ1PKohB1GCaTQ08wQ2//1/g0W67fbaC1WMu1hLIvl+7wW0zlNXP+PQ9Jd
o2vlfFrOzZDXuOzBnEIOYihOqFf+Q3EbsZWp9xGZ/Jp3SxW8FbAWnum1dDIct6dL
AkD7nI+ih6aEQ5s7dz/lgWS75d834j8QXhMUTfOiAwrmKHFcXxBqh1KPpU0I+MPe
wUtDqkT74rMOtNHVpo0pP1l9YEhlU8jY74PuCirzOPT9oi+9r+InH4n0EHrVZkSl
JGZxF36DJpLP0L2tE7bQAtAYeSVg4YWHfhbr48YLyMnKMNXXh3F7WH8LkWpydSRj
FiJcZaPY6wCyX5KVUKFoacjoBVKW3W6fFge6Eunb3u4NDF31P6+7N8n4M8jcHAoE
2o4fMlmfukXkvM14Rskr6iZv/pBvCqI8eVYWWdjXFcl8Rwjrch1yBGY0yVkd6q2C
+zjdHyCEYw6xEFhFlt6n3Il5nL/6IN6dSU6TIn5z2miEHAcK6eRjoNDI6R+3nvDq
DhLUf86MSRDiYStCVZFBVAaDAP5WnzMriqqXkGmHBmpVycAq611f+NFYMZT3wNns
ad5sAN/5NRBApceqXONJjpguQy93bPXVWlWRIgsuMoNd1Arm+aqNIWtkNtiFoz4V
TdouGN42SVo4JzjibHfmVskeOa17XGC/WVCMK8DNMtthV+rPrderCPq3XDlWYezW
mIGxVjUGtwTDlDEzmsCdGIscvTwJmS6DeIZI9nSSPhXbHUWJfvwKImEiNnrujVs0
z44wxEw213U0DNnoisf829UHWx68Gxd3VXrTrV6nPocDpJkSOqqgh8byJNSdv5gV
uvzWgCR17LaJuM/YdkEJGKgrmSJnMT8uTFHRLGtrcxkUInl6BvpBJ2LGUKfXF+S5
frRorLZHecU04RyxMfSCfTEqksmpc4sCJL8ylkTvs5dabhSInk6/yvw8je0seKyo
vDuCDPcoxjdQpbd7OmK7uJTjV8uZxhIcrcgaddV3CNYTPwFWush4kUSfmGHT8Etr
DqmmgodSt1ZRBvCr+IuD4IxBp3HxWcq0x8JYZpXXEPBmjtnFyn+ij4aLRkV9zFnO
gOjY6u0fNHt6wth7bMk/DJEGq6W0kCjrNZ8ETkizS0x1WK9ywJmS+FQDGycWu9vr
Js8Vr87B20Fu0ba8X8WosIJXbT1HQyz0320m0M1kSH+z7wv2srbw/DCOPOzUAwW3
HTEmGkvOIrkFq+hT4uompSTOuFzrI/AEYcLW0FQJ0xTLGAS3vYCeWqX9VHotHjVD
318dITXRO0Sft6p10ZhMYQvA6un4q7ZXf0pv+9A2ESHj9y5ORyyCda3YRBuReyNe
NfRijgCXBgiGzfZufII6Xjf53NFG3f1jCVamfFAD0Ggci4XTXnQf0udDmF939s09
iuB67AsC2mE1Q5Zs5IwcLsX4w+KeJXrWsYVZ8QJzjWR36S5Wq/1U5Tkicqisat8O
GCMVTyMCYRtqlWibon8nFSxTm445sBpqFJWQo5+a2Wkwx7NnzGtnF7Guw+p6hMTH
R4w5xo7yGjBvB3oDlar7ulF/b9ntP3yMJ4E3KXJVT+nsF1NHIEILX+VbA8I/W8vQ
RTN694Z68BP3lDGB8s8WgHIBelQL7vwSV5g9F+5p69ZK+i/aCEsr5XOfbI6sKVCF
6emmpuRsy914aavNez4nvpV/no8mJGxr3FCHZ3zAg8jGex68xL7FbzoB6khockSM
ujKJcLNbSrAN1SrcBAOBVCprcGQ79PioQxxarzQYr40TrmfxGiNgQeMEYrlimTHs
vpLqsePZJkmfOHgWfQWvJvV9xoKJQhEeHr+YAOsgPisgtDKZ1S95h5xVn7cWgpyI
4y779ypRajvxFovEr9QjBLTUMr3lOnOi5EgH0zLIrFUGN2rJN4sZea14oN0u3ku9
Jmqt4irxeXSCAuysq/CL7GRucXQWLhga1FnD14KTJZhBPJmdG+6xV4vFb3jPeg7e
gZTzwytn6gi7BJ2ggxAE2RIgzFAMC0Iv1izvDcapnQmOp1VmWhFGSvUaG6LnJzdo
XdyIte9CTQ0sWsWbz5h1160ij8wTgeY2DYQtv8PiBzqpRUsrjsDHsJRDzSW258Yu
+CxM3GEEA7Dw+HuJs8+zWeynETokgGRBBCFA+C0vJKfakFH3rOwqJSCs0GwIIRjr
BjCFd61AQQu80ocn2XkkAHeqSuV3K8YcfCpp7uANKPsUkF0ydGyiJ47YSPjkNly5
wWmKl18+OwLaneCN43eMPTfMFd2psJ1VvkG8WYoSAc6Tc3aSqYdfx3DtVR/9DzLH
I4VGF0Xm1AGw7q+flHmsmzP52t60uAr7QhIP6ztELx+TOMxQ3OLScSz7oHBulnjL
S2ridxuP1DGLCyv9c0nT4sz5U5L/Q+1iD1AsbntpEMv8L6hyOIa1ESctukq+h8/b
AAlahWyDwnXNicjfKihT5UkaLEY9QeEkE1ie8PKoWa3/Nk0C51B5hL+OJ71YE2ZM
ACuQujO9NzHS4l7w0BupXi4IytkC7fnJKDr6zwR2nVHXxyI6mwBfh/UfCyaBmP1W
yj4W/XHCank182WxEBAWllXiff1q1zyP2MwJjRYt6ZgSoSDCW4549Mddjjp8SlCs
JFpAIK63Gi3CuyQ3giiJHCwxIHwcJEjreXZiskOpEDiTymu/l3MzLaE70BOqIdrd
XWS4t0DveHQdUQCyXIqzXndhBdU6Z4RyMk6XjT3XsjVKoLqrJLJiu8+wNTIGRMlr
LLVC214BOa3UBxZ888/qsw/Ff+DwFGuKYVbAAW2bEaQPBnFkqwHkgQ2vqf62ClJO
3TgGQ2fjQMmqBfiJvks3CjUQWxxISuSYB0IeV2jdtZqdJyhUEokbwnag9aoD+nf0
9KooZnlGKwNaaPZjwg3DsFuRnAZHZsM2MymClobS0xw4xh5jgBhQM41xO1anuBg7
KYaELDAnOUwWmkSm6j/nt7VEyWi2qtLPa1BM+/Czt4Gt2myybtuDE+wt4g4J8DmL
l+AqelVq7U/9SmKdxI14DYP6C73gTloKlB90MHCBdn3VyyiCowLvYqxBVf82Jnrv
Z7qjMNn7xGEYiayF5E/xVWXMdJP/TtyNAgMLTFdrdPF5yulsuULyWvqNei4h2WJj
SW7B6ieSGETYqnSYL5VLj6iOcPLKB55RxCwpiTz1hKB51MFU//rNrPGD2n4vQtYo
RwVIF6DhHIHYd6vCDbw2wMHGu4SLJ8xJ4nkStnNq25a19Xp+UipGvLtrbNltgqj9
qIONJpfjY5oFLdCXV9tO2ceC9bM7blgBD5QRNKp2n8WxdOoO6FWUYuPi2ub33X6W
nX0akpvbZLFvqExMGnYzqBe+HxDV4EKtMOBjr6xiMkM+Xk+2uw5F6DcCqMEhVQIU
8uQWkLm+1XH7SxJV9AZLSS2NajHDWVgGECsGlQgPvyx0awHuirM3814NA9uGTVgd
xe02zq0x9XGEvGMrIjsPbRhlqB47vh5DGGFged3Qi+2xeWhIUsEfLbeOvVdjnhVE
aBYLt5hFR494LucNDSdhUZQBqVyqWhlT3Uhmbt4atPa0Ktnv3lP8YwGH0uGaC+Hy
/+d3exuhAPAK8jnBjORESn4QsUlSExW+lnym8PDKwSX20nEJyMf0RK4+zaeHYou6
1qcqTwCqp0Gh4f0cFwTqf0RA+OJiqiT0dOkMeEVxZueM7iqVLub1m0dQMpZmpkIQ
G9bXjbrnKd2SIwZhbhyRM9J6gd2pou5+ofxqo780qsvLWjp7dON2RnFlLUnVpQNH
0zgLpzf+oY6HOPXFWwBW4tX/s1TF6YPleIhWY52rPlchxG0qjL1AI64mwtbRw0KY
uZO3IJjPgkwmoWDcSanoMOXYOj0c4pjHUDi4UmR1erZ08ZZKsfo8TQZI27K/xFRJ
klUckZXqfDUAeXAbHd9C/nF/jkwLlIOI1183TaHe6B5m7GCdpTPsfdXv8bMtCJFI
8GIsIebLrEnvvxE68jbyo3jffpkyX1LIiYYAXSsmJwCf8rJYjgri2j/Zym44hP/N
5TmfKySf7S7G+MfcmLT8PA1zsWOOL19tbQA9xPzmdeqcvZExke5gRy9ObCWarHii
7uzNT7s70a7CbXdnERFuDZPeua9zlAsqtabqVHZmljZox0ZgvO2jU9WVO5jdTaF1
2WGc9+loAc1Kj4g4ocDQG+oUP8j3hUUUW213c/l0UkugXgWtaL2plIchn5Y4EFQf
gcHj/6Tx6jvxKlaJXyoLGnarZF+S/bAQzjw07IlP4waDRM3lke0J65uL5qz+KjR8
GVyeKJBvgYsUwVgLz+Qw3BMg0DqTx0rHXPpcoKUNuG4KEiDY2ovLrF7uH6C7Fpfd
EVk5R+4FxNoBrYXmI8pPS2yuzAwRmdh2Ai9m2KbM9cYKvndVuaa8+6JeEGFvywFP
4lpQEtYQVUYvQT/4l7oVshOkZDqmp6eBTpFlExJ1jqiiTEV5I89zDedOuAqo9wUn
4TlSdsponepklTrqEniLjz2yg+JMxoWEvHQ01qQVqUnizgW8TKVxHTzRs309bVuP
SHHDw0UqTGvqw2HtxpgebcU40SD/rDW3Dw2qZdtmC9gxRw6AeYp5Lw3KppR7azlC
b+JqXO7QIzwRpSBkbe8z6DCsTI9S8NHiSVJSs54T/HL+L9H6iLvI0+hTzA+pgBgg
zGhcxpRRAR6fBLPTq2AN4nZcgsFfJjKBb01Moh7o2Pyh/3HIfB+C6q9/KXfsKeYz
7E4vYKUmunzU8XYKeFO+daUg8Vxv7OOS3BUqhv3ffjes0S3dVw2ZX0zzuAuoVgEz
0+yAxj+QXKBc+aQjFvNKW6tLXxbzECOwz6n2IJH77IcBhu6RKFOwPgTrOBZGrhKk
bAT/EVHk1b+pGBH+XAeFkNyxLbgrlz3q7DilwZH7kkNYjzYyMWlYrnVwq+8cJwmY
ooEwJzI0c8BQeI18ELNXPjth7gGmB99O95u4x85KMlvhCvDeeLD+3I2rFLDcL+hU
bQo7HPStAas1ZOHsZrBYHhsZXH48DkR7blmI7Yjgm7eSPcOAlsW/lYq1Xkwz7z9I
4TffaIBiDqgIVuudaRYj7rf42YQldaGhn/6qoreN2/Ul/EdZKfn7bjc97x9MDC5j
Vbv1NUk0qrsh1dStikntilh+fsSMmubJIx+YstDXMv8GLTupHv65a/dD6rvFPYGO
3yrrzpGJX399D7E2Vk6B7H/sOpb2frIdT1zESh21Bk2WVpHQjW5ib6zr0X2A5zDR
xKF7a8Rx4x+dcV5ky5UCualhPJMZtZ4Tt/kefTS43l3H+g/9D78ZIEUEQEa0m7Sz
AUoOb09njCF6P5IwxGg6DOTfCqmU3MytT6lkzaVfulEOJgyABsoESZZGO+XAb+n3
KHRNQvykBovzVilWiWUITIwT4Zhz4RNXtIRi6gjmrfxqs5Sl57pAgCIDyXsdT6mw
diQGRvcfodFJ59y5RWRy3iZWtyWqBG5zwqzP5LoAH9/0OrQ8SN5CUoDzL6vcpfTq
ufb1YMf/LmicKeNTrM3gApnBjaqHPE5WKSTf8CaIya8+VWJJ1glQYaWEcbzDh35r
pNvx0HO82W44b36KOjFai6nCKMS9tHO/0R2zeMqp2t+jaTdzyT12wShwv10+afZu
gMJ9AgvbIGvmw5Ow30V/arbLQM9eTk4v11Xtn+RGt1yFLpscXvHJgRTKHE6sb8Ed
9jQWKXbBomxaQ0bf1kwzrVWPfROfLUg+/fqM2j0T5sYKoZlvIsecCTS1xOasBa8i
fpYgYQGz86sB0C9VBlYDJesoNM5vrESZg5kVtffgfX2WCESjutb/jE9E/BP824ln
cx8mNbmYl0Bc0BM/V8PrGHCjruYo2xiO2qVfw/BSYfbGxnQr0XrggjvJtCS4OU6h
z3GAgsykv2GJ6wtDLsflbNZb9YHu+TwCM2ej8NpiNfu3bDt2aGO+8xl1Wp2fu4CO
7vbD+5eE9sCHp0OrmbArZ1cKixbERVqeRedCeSQeKro1xj1pfTlasLn9UsNKpibi
Cg9KzPtJIzdfCTfS95yN+3iuWSV87oIZWOj5yHTtffcw64VrmZHs1Gn00VpX5P3m
7m1XObUFJOzg/8nqr5hqtHST2a9i04CFFn4nFbz/nzMSzdnyX/JExa9Rkcef3B8h
UnCIz+hqIPNSlyXqnXZ5z2EjT4xjusF2P62cjCmW346IkQLCHqz29JFFhG/yFnAS
pfxpvkPC9pO174qE4BhlgttNp2O5uVuV+1mgtO9vKVDZxgsIzYYXYBtXFoJbWiWH
SbLQjGAC/UVhCWahPjc0pnSVDt6Tcj6YexvSrijt6hzi/HlWN/HSGAZcw4Kqgk9b
MW3J8Uvmr78G6HI+D2xFO27phqQ565eYNxPQoz5QjPSXk5j5deStra4eJCI0m6CS
vyi5wK1xAmQqgBalZ+5Fc5IGi3L51+lgU29lpM7zmzVS+jc45rSXlL4r/GhX5bIr
4yBHYAIjnvmfibWIvSu10Cn21OWPSO+cj9hM8EeXyJpVZgCOHCbZDLaXi15fbGaX
9F692ugDw6WacdWCncAc+EK2wwap1fjGB3QPC7kgsHa0KCzMUNESAeSvlEAb4xCR
qSBldGBBsRkP3gbgvOvx3QqJryjOfy7Xvcs+YH5OXqHfaP0oPbcYsZZJ+HW/65Us
7axT7HGj4gdvcBLQx6EyCzmsjy0xhnXRVSYDBz0+pRfsiDIh3PbaCLiw8LHuBntH
exjAmpu95Q6K0rmdwG5smoo75o3rkpZ94MRL7Ovd/Vu8cIeCh8Jn6UsBLbEAk2RM
lGNx9sGhs9y7Hum9wpB8OkhEK9gSQrM5GHBjpp0iwbUmFtwO3sJX6YoBiNko5tG9
jYrHkZLG6nZURXTukUm7K5jPaGeEpa6BdvyZSsrR2S1ysyzARVTjom5z5V17QOWk
BI9L1hZ4gd5sEdJa6e/TQ+wd9RF5BKwVn51wHMF2kjm9lv2MeAssKjufbFwQDQOs
Jm0c6ux9zYbEnH9R2NeCGxoTj/kHhhm6Th7pf51NcAQGzjOHHDirWyRMXWSdYpCb
lATdmC8pSdOVKX3+Do8gqzKX9NBuOOKSY722mncenbTJAC6i1t83A6A7Na5//NpR
g1r4BOafdHdECwvZqvz/DKV2KPZC6lEkB7GIqw1qXXSQxo8tLkd4YNz48JNHyJlo
2oN0pcFMnhcJlmis/ZK7UasHu9onJMK3hXw53aB1viKpgivrd1f0ECwalOOtIxnA
LgnIRZiahxqakgKAOUaHpaX0OOP47pKojQMyZ/k4Py7ADPBFiv8kfE/4i3HelX2V
tsWK7SLotam7jDUvvu2oUiX3PKnSLEJbnTjz0Yawz/JDF2qkh0z2mEBC54FziUDt
XiQhr7stqtyAf7/EcE91Xa70UFbgyqLCR5LXqcRhG2efdbCNP7lzzrJrHmoq2HjC
Bae7eZ8vDSVgF6GOyLuNAXO3t2vMnwQEbgPf8Dvwh4F1k5m/4qDyVDjhZIlRMQVZ
VfPtcKpA/DPzZ4mLa0gHuh8Z6z55v0IQiOuWwczfUEZqL8GNJ5gBztfd+sVbkzsQ
113mqKn6XaX9HINTDxVx/oVQjO0mgwCxAiCw9PX9c4DkTfFLNTEBGeXKjvTeCXY0
NP2BCyof5nNFiFNTbi4QR37mh+7grRfPzAwZHoGWxeEuBP3het6OZYHrUy4rb+Xc
8yLUTxzH3Ea6Q71WjFAb281IP7RaLYLGJFjllcH8e2sBxocSWWWv08KkO3gmhKd8
YMSX/DGE2vSUedj4nRsf7zsrhZOyO4iufKsMWaIZ+YQO1SDwM7ArIb7yj3hJyUjy
IzCY0hrws/MdtEu3XyYFPndmplInopvnn1hYP94Jd3yZvQvv0dZF/rZxfRV6JQC5
zZmKZOyuEwd1YgHki5jp2lGNTKEoUtj+VT/hRvsqRFKgYAfm989c+K16gni9QnON
y3GW+dlLzz093KimZZA6EtIdwwdqbttcgEUsx+RlgCSbu9viUgDeUOto2xmf0hFz
oqC8UE6vQdioTodGtKjwryRB03pCDYWrwa9SzAc6e+OHWp/aWrFj99RZCZN0R/NH
dPsOOo7gJknGD7fq/+Y4BEL7whCfaOF1kj62QUEePxAp2CXIeHeMmWb97YnhdZ4e
tJmZ7anTQKayBGh1Z3H8iH5UkMMQ3qXI0oLg1Qrpz7xwf9hZO7jXIrxVJsmycCdN
qhtGB53BOW1n4af4+XfRSDZSn8zfkRfVQ41rQEUb2+qwwsuC+7vdObBPD+XFPshH
SnWAprPvsgEIC6zxVZAS5ZUCnRQpb5VQcE4Ak1TZvLuRuaadNaFzGWSQbcc1Rudp
CobZyEAlwxyYBgeK3bhgrggrbuZV+pRNtcjtLKnEv+QPEsw5t693RD9zqb6fUi4a
61aZsGN+8V7N2XeD1+aMfd22nvDWzhyDz2EguwJavs0XCCi9mqzG44IAMIUkrscY
5SEQJo+VkjSg+8rkgVS/x6cQ++btR97RRKBSDY7FdVJ0TTFwpkbZNdVqY8cwc0fE
nzM+Odb/OcDyza1QXXWIZjfYPJG9pjDQB45dl4AvcFwIQ8ckUahtJFMvb/AlPun3
iHe2E2VFC1+eBVA3J/fLjlR4ObXJngJ18Z58XxlmF67UgDvRX44tPY2DtrNCN1bj
QaJL+I1fpjAcKzPoTbd4NMdHpHJat7LC8EV9AoQxbo8TMkKP3ZTyuHE3rsWdiDNI
kup2VdBSlol6w2YpQwQ45nsG2qvAHwtaZGvN4Sdpw33WmWG5ELInrfJGGy4yTjaz
uvjuRb05XuaZJKS51Y99vfuuGjdLgQWkUKxQgANTDyaur9Zsc+njy3XBWIZHz7TR
+i9eGfSJ4UqmPZUWQFNX2768WCslIckNRf3xhPQZE5pPo2Ohmt+njWSMKYNrt1EQ
jy5ogNi8HDDh10ewmR5vDrQ21C4Sjf8rL0xQaUHONRpqmwLY1u9FympeLoVylqiD
vMga7MCx2/x7fIWqgHfKkIDs7NU5roDYkqu2cTFjKjBadEkU9zcYr8ZjssB8hwKw
hRfqfYOLAJUbZaWDxnAlW4sWMZYPJPTQ9daCy8ahiHO0M9QTQsuhU8IwSCQ19cFG
yLEiJulkCQEHrH3ZHn0gX6KK6U00EilOmBKCqcadksfLzJbOWobI5RJcQLesCSz6
d7RfpUywElHeoLRlBQtXrFE+QKYibSRGoQfodsIuEVt37vTL+oWbjd2M4TOJ1n16
s2cTe9WIS/BYHcy8obuSh0JWTkze07R5BKzTvPpHxTHVf+smP7+jakxPULi9PKP8
/bRfVqN6O2QkqrmAUJ5vFNo5A1ogCdeI9OvqUFeJC7MHmzs5FfJWPkVSg7HuD06Z
Bd4Ph7/EDhHPCwUKa1IxOUbn4ToeCTf5r0YBYJi4q8+Lcz08eQyUzZS/AAPaM1gF
PsYeDsvcnW+Xk3sjuDUI6FPdXXxhtFsFMRF0U97vprx2fOd4UPiLDarnYwYoDbVO
17epw+iuyu0mPSDrUkCohW/hW9JXYJK+n6/0GM/GI20fg4sU5OJ6O6Brjjqvlucw
haU26rPkAsf4EngfunCC42YIsRluVsTvGOPlqsV8BboSkzwmFg/v7X+MvFns8F76
tTPqec2T+Mj5FwybaaSdsEAlMXjiMSz2bhB/MCL3IP9K+rv+qmiI3pBgP8LeKopW
A3rQcAMQBRC/DBOBnoHOPkF1WFnDUUQfuO5TNJupz9GgAsfC+IADfrQvFa/Asjso
KJHcDIyZlmsDzenW9NlbI9uMMKdXqSba2jQnBXh9j8z7be9Q3727q2O3ihk40OAn
GVh7fPnHfuvRth/rqFFr+8NdgVb6z4l6TCJZ7BtaFevW5ZIT7Gdvqg6TTmDb971f
xV4NhoEcLeRI16LB38Sz9umqUx0jSa3pw2UZtVA1kDafZ4NJqOOTR65gciLBQ8hv
0V3pSXa6HTAMAILu/5ytvHIt8xW7fYIRGU/GZSxMnzDunQjYeVss0HOxePu7JdHW
+TA2TGdW5oyIc8U0LtWYrF8lUM9z3eEFst1cGDYGTrcS7MbESSyRgUxNFXDSz3n8
QeAXA3qgfz8kvXOEf4TMdTNHaheDUIG9qXhRtX9qlKLRV0rWleVP4h1j77QvF0yH
4Pb6P24oZ+B2omNh9fnW5lBqLvEbAU2z0NrjA14IaZnl2KZ4cw6hQFIlsM37PCNn
jJtM2NR2+FZCG4IaumNNcq+7dbpUFbmFgra8c4Ltk1VpFzfaREJg2sROmFkxyiYg
ofYR85+8NPbhwgoVf7pGVIqAgFsZ4HuHGoNm9IMqcqDro+PFb49ajkiN3sQZe9RN
KMCFgCCLxbezXrdj+YufIh29ZEZcbkTWwLHB8vhWa/IyWfQuik+2XDT1CdrKMOPM
Q54GH54OqwvlNaAjQ9cXhbm+SMf4PrBYQNe8yj74XUo38xaNuQ3N4lvH5OSbIVgF
L+XixYVyFxP73hznG/SSe7bKyRm5OYIsnWjPr0rZmAppNgEkAJJqDxv7o6tiDQVF
28a4Up+jB/Yx4dzy+eIm6Hf72tGl2/X1m/5dA5JPUImfSDgyDt/G5nDV05U972u2
cxl+T7y5aIEpQUSMJTE8VSezW0I3lBOIAVb1s2zf8aNPYSsy8TOZge3buQ269Dkc
CO2LKk6ToeU0wJ4BMkRwg7WcwWCj+W8rRw8fK4tT6HaA6kUUZI80LKtinAQkwfeA
q4gpzigRbzpHSE8iTAj+DSaOmdcFWMbgoLDyhnVhLWC22dk29SJgfprAvIQ1JGG3
4PIzqTY64pLZ70AUWm3AF181F20tPIZunc59EgEqDZy2PrLFjz/LBFOK/Nz2IDfA
nHjIDt8JtsjsMYrDJ1kzes3oxc3PmL3qEuqBwSDDiqYkuaR5e9IM09cCstUGh/4T
JIyJpAr9U2q1fkh6gtAEL1kRKwzDSh2bo0CFACNYbYzJpBl2jUOOVjw4uY0htNEn
I53Wc+fNwu1+ajXK0jPnpjIn41sEe2VEtgQV/YG2XUKm86UStEHeIZsab48pRqLX
v2+WKf7u8A/bYSunN/qqtRGptqC8aykQWNSqKWvnGPxmcnPr2eZ0MGXH1aiad/w8
BBzTJe91AkF3T4n3UXAuJc+SYpAvpCHpKnc2kHgnorzZqHYFGlIVAeoYnjGWMhZw
nM09I8y/l38dj74D9a4piFTfmRfJR+slxF1+zaR+GsDL4BOjg4SGSAi5XU04uKoW
35U4Y+uDqoKmiG/IoAu/SpxKrpgmNQtwEaEB9NJ5gccSYP3YRHNg7XDpAJdEgYM4
fpMr1GkgqNNiDy4CsHFVJzcy9G9MSr6ShYIJPrpaEZ/GyDyI4CgPxA+qx//zS2Yc
SsEj9vrEiFDgIK3nlqWFiDEvjb1jeHZEm9vcq5+v1DmMeB3oUVhOPU47RfmVr4lk
1R5e3Q+UULb2M2SX028Zl/h8nEjmMtVrsb7ptz0v1MzkxUO8sZ8VFR5ab9qndUSH
1ad3QtBYT8wC9yLz5XHjwrTHDv9v5IaJ/odP9CCB4tkIHejrP6jdiY7/h8UleKOG
abRBDdPUsu0ns8q0PtL6MhOtdUwayKjWacgvhmJiPRJjBRRyme5WcmqEiBPMR1FU
JjQE4nGEFJCNq0WhId0TKrOsmKUfPqslzl0c5IW/yk4r29I0Ml2prJpfcD1+ce4o
4Ka2dHtdJOaqcNgtDxjMfpS+4h1o8YRulPZSbHv5NA6VAed5kVu/u2Ck6ckeMSZ4
m+7yT24SPHdT9BJQL+DrcPTBGYAMXqMYEFdrUvupq4mo1c7Q4x0wQpyUqmLE/+U1
mbzSg0Ts220ICcS3hBT5a4L4Bckw6dl1XTOsSYscvv4+cVoNpHFRIM+NxH8s7ltY
N8W9XZ8q/4jLBAkTvQQdn+ptxCNdTETdOYoxeG4mRciOSkloJZzESkw1nIvAf0Wv
CK6HtE4xap4SBnmB866JOBYhtokrd0X48Kj9XKaWEvz1gu6vs8iehKg2KYUYpjQP
jKfEweO6aantqLZZiZaS5JKpb2UzbBzkqJIcvPZNgu8Gf8HgNOu2ckthhV28p7xZ
JxnuzP9sWdTwJazyJMvgHmZ10s6KUuEw/YtMWqHdTBQ13wZYvSARqsT/VpqTCDa4
MfL35//mgX45R1NH1r+rVqKcVzqzVEYVacU7x6xWDEDgvTmFfXgAr01ou5MBrnIj
DiB/H/A35SoYiiLJIIk90ejQLuXryW9M4SNsn5OePp35GYCM7299VPCmsrHOlZFj
KZimv88gW3d26ffqsXfBQYvyTc62tQStRLiobyD9ubpwqY6F4unBBLESMNDhtk9f
xPpENeipmD/17pMtj76ziNms9MXT0vfd0fTx12LHzE50OfNA0IKaivUnUPePlkAn
BPujOJSqqvl7K1iuxNmbp9PL2G4sCm0uBPqYQDHJpp8XIUNxPqXIpCWQq47tyaia
gMAi9VzLdio/SChxt2W2QXBnClg8Lk87BSEOZSvZVm8IEzxyk/pt88Cl1flRCh5g
zfkKq305PxXm95upW7UcjjhmHHJyaUoq6q9UXure+PeQOVM82t6b6QWhJpgiNieU
tk+p06JxcatjUvBlNWmU1EogbF/D8E9zVeghZ52YIeoay0ly/AuRY2/shcnHaaiV
nMa3UgnWYMDvXtQiGNXTpHF6noSorlSn7YQMbx0m5hBQ4oBqSbgMD0uD5UoJ0y/Y
ufX99pVe41kLwpA9//feG52f5S9bFur0FlF974+op/8awAD42YPAlz/xkvM9+3UL
HjsizrieZiUfvMWSAvGgqgIj3zziOCqJWxb5lO+BGaMjU8bYiwRxlIZhC/QMkjvl
SWrqaLA2n5QeN+pTukc1CIh3YCDGbL9jXHOpjtTQqUyJLup5fStHTWf5jGEn/nkD
d296MC6Mn4TOj41LsEkv7xrM/3z/M5Pp0OUUk69g6xoY+PW07a2KHzlKhWiBsoOY
f/i796Uk5JP/2gREJv6mcxC3tD5FjNEw+fXXSk8RqRHBpItgxxws7KTx2IAQx2tZ
/ZwcP04TLVmoRDc2QBb2sObc/hZvQDCLHNVdMNF8D5YuG3NWeb5z1PD7LurHMwdZ
FROhFVFjHhw6uoq1lMy1egSV7UXPVwO9I9/VsV6NNQJgAn9hduMsQqkDWUsVLzQw
c9m2rZFkHScErzNKXwWhmIjNGn3NoTWYgJOpuRCJPKo5nHLvmstc58LMjuLhsA+x
kqaXi/YXJa37JJoaN2v5YP7mADzqxYdPCry9v4Q9L2q4ScpT3weZQKE3ztMMZk/b
SVU80rI7w/76jigytYhhkj9Fs6BYQClMhFAeBXGWBy3CjbmlrtdHl16xATAxe09I
gI1jGN2Ro6jzUrlgYQYD5a7F6XBgz+c5fTyjSb7alc5u8wOA8nA9fNVdMyuwIx6l
HgKZfiBzpNFfA7o6+SqUlwVw0uvYi1FMzB/jsGBGU8S9rSTkbLsnVx/eIbiVO4A4
mruHr0jp7glb0rEbPBMI29N3cUfPRi+FmGapaLF0VfJN7mNDB1XUS1ObcvXr7KLZ
YXj/p2MkcCkYv2XEXP+J3hkEDo3SnHb7HnFZzDwkMKqfQNtEHAc5TqJv5iBNjJ7v
logancnp9LsOAWluBbx7pdjQ4wAYBm5cPdX3+CBv+esuxv3YAL6urv6jxepV/nYd
iaN+U0+XcB7Yq/KAFQnrMfB20dagqXUb3Xmlfqpt1YOdDAENRUrwwK/c/xt/MNEv
vw/JkCudHW+mrJLbnWPZLAPiYcjLKh/xBH6nbTA0qTSRltWJ1OKes1b5DzhMZG/R
nMn262XUZXhSiMHsGBoiJ/ROGnAl/t8Bc+mDb4TRLWsPYdHGC/DbHj6GE4UpjZqW
2gsX5/3KsOkGukAE1xOsebVA1JRv/gdrpGtP9u/9zfCicH25iPDuT4wt9OVrgTfR
im6fyqozmS1vaPIRue2gqz2r3jm1J7jCHqXY0K7rZiC7zmYREM3OLBJz4pMDVCZQ
1FgCfeS0tj5i4pvj9yxudxm+V8I7zEEbenWVzXovlMoETpSYU1QnKk963dImVgV1
6jNq26fjNmaIC0sp5Abs2/zM7QLpN0KIc/sezps/cJ4dJV8ILrWXs0EkqOHVre1C
sKB7DF5CHsHE+ju4J+Cy8BlPlUiDPMY+plbAfEXda0XaXpuZN1J9BVSDdNmpOWo3
Gzn7P0UJ9pu1yYglKQdpKi4GTS2h7Vd26j/N2+zE1TigV+g8Gp0j+JYbWbmYupHG
NnEUfjlH50kIDAtg4hU64wQr2hlhBn9lyricQAdBWxucFkwCFDMtXhI8yemnswNR
WtbJABBqj8LDOvms1/QJ/mJ9lPY+Hp41cUeibDBI+ATBR7D5oO0KIlTRe75uxu10
F+zqwdWNi674nCfH0Wc/v48reniSwHCsYMq10Ns+uNxRK5OW9mqbfwv6sEFpuxp5
L88WRvtkvy2qRid4fAloOy9fNgYkkyxw1JOXMvG8Dv+efdUoNmXgKS+3wHylP7/6
fGczyMFbSFi8w8EZ3rpEEfFX0PjZs2orbeI5ar2hKYbsHsDOuJWVH30vYnAgU/Bz
ynMzup4egkX8zB0kZQsyXH2OvE2P41U/Lj/5BSIDeSlUNSeF3ZPzPJjW+YZ2nafA
4CaarK0I6mIvoc8gxtEo9c/3TRxn0JJO6kiYiIfDoyL4yefeCQOWl4nd9oFvLC9n
L7CHrLIkj/QV20opTiXFO6sCS55OaAbtHO4vMn8LpWfVCcTvE3CeAJxnXIgXn+D9
OVuPuVK6pM+7DPEOOKeU1V48c1X+cKdDh5CCOqN4ajwPwZF6wLbhfuFgZOF0Q2JB
fEM4bivTp7ANR6lGDqJBTRCqm4plexbP3S+XdXXBsbN3k128fMkLreorLlB6yG9W
gUQf/4QXemT0r7rGExhwAACrDViZVHh+TFW8QnSoesZ/i23PTe3xmWUe5WdcNt21
vEsGVME6eC15mYDYFIcOvmQW3qHfZ7Ui9SB5/MX+rsfivMIZSCT3hlwusAoOy9Fw
ki38uSFpshYWJvyEktYNcOCki5OM4GPz9FRHtF5UvMhMb7BKJ2T29495DzngkJ1h
zC5rMctcKnneZo/FLOl2hzaouIzViPh2zMQcKrLs8wLLKmp3RuHVBOCF1OhxZLfN
NqYJusww6wlQbhOb+hkHAkHcesLwLt/mqe/agBhAtFDWjGoYQNp7YIqpSC83EVMV
01UP0X5SRexfCGfwWzlYYNHZ4Wf9cJI7wjSG//d3HTCxlloSEvILLDaG+iM9vksc
xBj6nDN1HXRdWohvWQK4L0ZucgdYamrQb16UR885heunPf28f1AeraAlHfadQl8m
sUVxrg8Q1P05h66bD6s9vXRFP1h/+5k4VzMt+rStz+FzNOdccQ6vcAi6igverNnd
X1QCLouUJNZuGDtlXXYUBBgqrSP0pPgHkXYGMHB9ZJL3PVBM7mbyeYkeTCg0P5K7
peioXNZY8zT5eL8W1oVsxq3QbvRZvsQN8fDlAnXri9Xj+wKA448z/9M9qHOKIW8z
CK/US1Kp6NjZCTgUWRDt2ZIrdAQXdTx5MjFoxVKrgd1gjc3gchqd2sWeFc0o3auO
WIC7m+UykxABTSi76XehN/wuQN4ZWiBqKQ/FBjj9IJbC5DbtqwUwgbt1XNW93mWL
JvW41uS2rFle3v0d6kZsXfqoojCUSgVM9HbCguyWI3jzRXOWRFH6dREG9+Y7bf0L
lZJOyFjc0y1ahWgvNftZqOxq9ITqRjcuixxM7EhYM2Rd9eMDhhSOBqd2elgl4UTs
aoi0fi3Rd/rwN3/a4rrAui0olzIymztFJkidrvQYf7DPQ/xgH5h0hMcNimFnoxc/
hCaWB6EVNPq/sz2X7vClubPdbfcPKLtufKmof+oSY3FS+sAMFMZdHELbjH2O38kC
BMv3FXU9NrjaYaY0as+QOda7C+OHm2jqqXyb/XWr7emxXv1vqqpYzVgXs9w3rTg6
m6h7OhR+V+YR1YREBGXtsFORm9ScshOCcg5Msxdl+YPcU7mUsGxVNEJZhGiO/LFi
XWxy6gYORgEsLYiChSuEDHglwFKZCk2MiupZTK1cOXMHseSiks1gb961Z2ySy+ol
C04cmbTRny82yOlrie3i68l+AF5qDO0f1L49vN1VrDFS88xwEaAOHqGAcVMJR11e
edzplO4TyptZlomQQQpzGayEB9D/hmgr9bO9jXH78+97SkljT4g80yCEmwR3pvRB
cUIruMFWC6RtNoLtQFjSWZjQA3gvPpP7ws6ulDI4bFJOiQPnY0RRq6pN/9URXJQy
Qdbv5MbqADrPTieqDUDWfdNcD+fG1KE4h8tNsUTIjF24SQvOHZVFOOJfEFdqVq6C
Y23SwTJWIrvBSRz2kUxI8WqYrB5vfvJi4PR2BVXjmPOc660ANOtHxGUEu6UQRdZ8
VXko7chyKY2UsyHh1nH3X993AEoOroul1IV9B2cVlmBj7tlFkUnQlIrxShelKrEU
Y8jkhNgEfKnjEDbz53qU1Bt/itsR4JnvNhcbQfgLmRTEQlRbJp4af9GZLSAsO3IZ
6sfb6WfQz4xMX8X/nSbpsKJlzJoBbMmxGrplXfylJ9xEPT0e6Qycix4NNM2ltf9A
HPpnhHVilI1VF0g6Q8aPYBIo9gTmYDg+Hnazi8LuLIpZ/P4Kg+p2oOF8nedYS110
BkPXVRySdUJbI1ZIOi0UbWmWlYG1pexIx6yeopwkYZEYkVuFmPifgwUJeKNwaM7u
bHTC66fudwokUU4bPco46hR2s0QpCsxVhAaz/1oWgZBT/GalKRC5r7U+XclE0IUA
VyISgr7S4FreEInZlsl2W6MZKtLFeWYLBZoYL+ctuaONvC4S0q3jo2247wjZmYgs
w9phBZY8D0IB5Hx8NSj3jMSlklTOV+C0A0OkWQaZtJqXHPHSvXWk+AR6TYsjNUe9
1+UVaCey75HRyq038wTqByWiCAcms49MALkBkvL+NpgBhhlSB+m+bJxaUPY634ZD
cPKaw+6ejkukPPyvzAMjBa8zveqsQiLnLsypxvPIhbl3OApNWWC0UX5VCP0m5c1V
nF3BP6BUXKDrMl5tswp98Ai5YzNzkfBz3bEcMKMk6noaOZXH+dvzDso2unUnowaH
ve/XFht4Ok2PGcruj0nOnB4ekqYOF9CnI7xJ9DhKna2ZzkYquAatCuob9YWic+yV
sFK5isccbaNRF1qmBfBsAqL23QSlKkz06H8577+2y8/hlzIkxW3EW1xhLelu9lxT
yD73fZL2alCfbcvdedM/R/PFzGsXPIzmOQ/rdaQETz2fIYTB7zqU3QPvfV8uRUt4
ygeqZCZCS4/hEkPzekQh+KQSS8kqejTRq5kRrtnQLSlDZebzteBs+UcMIbkzxflS
TPYa3LzpbcZTaCXcL8YloCtoCjX3F0FF8tex41Bhjp1+QAhKMQGulMVJ5QCilz5f
Y+0dDZ/yJpIZAkstMVIcbUv13p7pnUmDte4tldfjffafFRlFXuceQaEAZtfgVnXE
CcR3DzsQdYld1M17U9d+ECqVBJvty86647WSlFfHxB8LNelpfxIliTc1vC7bsxZ9
dcK0WRBWljaB/hyIX+Pm/9NheJBQ6ZR5TDw6zT8PKK5JzYr0tCoKHSf8Uw8+rzer
xDG3A8p+jFZ40/y9poN/BiLYur8oaPyPBEccmvOyQignOeeh4xZgaUOYRMuSxags
JK9blsrujrLT5VrTMBsHtmIDynafR/WmAOvQ02vrud/EQ+9pbeRIcEz5AI0akyTu
HRzE0Jn+qh0xDPAZTR9aW/ZWxmkqWEWMkaLdL9hEnNKudKmlVuSXr6vlQwZOS5lX
kui+PJs8VuPnhoOMwATeujw9eDtwr5gPVpAebQLL/IZCRcFfbgHCrT4mvjLVshVr
+OuzZ7dJ1q4MNqSRrHtf1Z2QY0NUdOJsafTaNmuW1XQUJqYNJ0W0b2m2i37Cgq2O
vFvPZA0Y8/f1HIAv4rGLIZGth9DjlXmemLmC5yVUM5ll/PpUK+JvckY7ZFvdWYcW
NWnyvOmP+U10oAGsGyrkQfW/R6IEVDq5ddDFvF+UVbIBs9haNzSWhCoBxu0m61iq
R28qaF2xHFP8XGOfIbANYj5Ur2HvNsV3joLA5NopE44s9XdhHWYIisv2VZnUEreC
LgynudI4gwQ0O0zC9MAg9DTsS2TvfOCG6tN+Fh7qc2F/rMvH4yoNJmmgj8J3zfI+
qRp9F5K0RB6IFS3q+M6PD3Dh8gQgkH0wSmUCsT937Bk4wX0wijoYBosUbW4tFbvL
DenqlIywjB4do+IaxrjuILrf7mGOZXYKRW47189XXkKK+855+xfzheQlvJe/nI4Z
DH3pp6BXvGbsJukT4wqI4iILxB560fo7t66CrYkCLt0zPM56HuH4mX1IfYZdximK
iRJHUkcl+L+X0IaBbXaps0R3TjVa2pwcaUR73Qtyz5GzIWGSxK5jlZvbA5pFSin4
Lo3/KxD7BVtrJPEJQkGD6/7PFDwadsxUnh5TmffsAPc/0JFK9h6iROYF1c1SCs10
GAs2soynOxdDkE76LFfb9md4U/DzWo1G0xMZncMgXC/e8qGsvvUKHIWaqOAAoybt
Vwr4F655fTTbfEhA18/NPBA3YetIAN0I3b84YPHmCMm3o6MXCfk0VH4e6BmF5gKm
pIz7r/WFXDcWava0rfox2E7If4R1x5Ci6LBqtucAJi+91qUTVc1ZfwKmutLRNgKk
fp3thWmIuXQbXR+CCzj8AnfZXNhps16FZZosCOMCTiwm8QpI1MoReXOAzVBCZqqo
atC15fpQKZqk6jQTFyWgPcQuMBLhevZTSDrnYkKaTxjcnQelZRSDqEcjX8PUSS46
J21A+BE3bKqNF3VR0UMywGoGiZSey702nusZ/aTrumtoidN7SpmgeAmC6+bzgR0B
GG2pqgtCBDk9qOLOfykYzBNq74Pc/a00N1yDM2rbpTZXKBhCkI9+13gkwGWRm0VC
sFwVJquGs6LGWzmhkGKO6reMEGC7L3UUylxMvoIwTvvFmzDRjZpDs5zReRxxf7B9
Q1iD96zf1mnU7xz/4xqsz2QTjmSeRKl50z2iE5yuCz4aQrdEK9/j+/KSsMVvjs8s
p/3lkWbOWYn5Q4Ur6NtAGuRw33zie56J/10ixBTAtumiJRx0MltoiQz4ZupRjzEr
4++a72xBu2XeCiPnDJz7jZD4SBfpIMcbuXckf9sp4q8uupJsFy5ATTMeNipYoQXv
Eq8k2gZuAamJBgh5CZRfApIu8Lu65grls4oaTmmYvmXRwW7frDlYctEuu7xIX0zu
ldqyYp2jTkS280ArXypfc5Z4wrW9SAa1Bzhwn/nBy6gdcxtvO9J7U4wNYDT3ShWX
+3ZAPy+H7TvCBXlQ8tYenmD/jsW1iVOyXCFoR2sPQBAT+KnonIAxBXcGOa6nulwT
zr8cs8LI3KaPIm9WS3fSDFS9IrW4TNlpGtqKuMowXrZvEgiMGAVdnDCBkKUkstdX
L9sqGDUuC//1l78SH9wFJVuKlUM1MY7M/TsIiHpluu9Zf+jea6J7w6pkhstPp6eR
hl/tWaz0ZWcdEoi88I1qjWrEb4W8e3qEmlai3wUCk7etcpJVdrfeBGaEk9D7r3Hs
Aa0bUoPBZo1Sn4TDfT7T3ODvTQflNasQVYyZj7ZVJEr0k+THWe04FLQu1YIdfp9R
yhshEm18LsEk61sjNeAGtJxvKhcHE90HBeMc7tM5fqAltXTsJN6Iibii/h8AbsfE
CmtUK76PTRibMprViCSsP5mIVG/aM6Ft8v8waN6G/YUWnIEouyqaS6kZ35kam6MM
LI6p3nHJ7IH3zYTgWkKKmJvjXOddicb6N91Nz3RsrVp6bYOpxc9m7MSqJ928oRp2
qV0AaKPuFt+efRVmfdL3ZONIXJwHV9KbSuZCap9nopjVWrf20yfQlHKwcSB/wfCE
8qb2sjdLvlja8N+Isk+vmTCNcY6quWqfLHk4kILtRGIWXaox3E9kwOdtWBJdXeGQ
i8UR7iU/lp5PlL35JNTiMtTmToTzeKKfLSUhK/vxnVM+cP9hdXj2tXkICmpZgw1L
tVhuD/foah+LMrIJTre2x9ZnvovWcS+v4GK/Y9iDWzHOftthblYMOkw44F5K6O3U
FesfK9IjaCkh2btPDrzBMF/fT6dpRZom9Qi1cWJ/Qm74CDFxOe/YptRZlPVKw7i8
FrhoOQLY8MJeykkCN5K4ixY4w3e59mFgk2PbeopO6fmeKSvwChyGVkqGQ0cbC1CE
YrSqiWwpjEDCyvA1PyNPiQYQ8tNzNH4wu3XBlYpPsP902twu4cHQLdigqHHyeGDg
AM1U1ZkV6PxPqdNrszKAntmKQvgAofigTZoHynNym18u7/fTwIa25cYgvP9AJq/v
384V2ncs26HwV7i1OcJMUFtxokZOuSMr9pypfsrxixBm2EqAfcwg/63acMnotaaY
Meo+nM4lbO5uMYuRHT2O0XwbvYKsXCc5puX/aVGUqS5bxiTX3d/R2j1S2/UX9tEu
zTj4seLa3Yt8wvU1HmpdHUm0vNg/Igp6pZIrVr0d1OONeB56vs6ojnjak+JeCcf5
siHlQrqDOXgqsr7nslanJxK7ueGwAcGOTU2tjhrwIh8AIFOQ1y/V1A/uuOtXGrRl
A11zYlmz6LKPepPM098Jmpo7xifsMDDnqRPuaqWx+oFERoqNm3vvuJCaW11PFhMd
X2redr0PehDqC/YR0esCWqZo9a9CsTHwKPpG2315ivb66KdmRdFsGz5pLDbt23C0
6DE5okmWwXWs3qK6rIOjI3Vo+wf4ceZ9z018QODIsquc9oBOdf8h+40J9a45gD3h
0IoP59boyFWMQ9ZnpoZgQwFs0o4jYg+kR1ZPwvDHZiIceQ3zlnrdy4TPnwgizCuQ
l8ft9V5iWf0Ndq2JU+/TxWzhZcJGReliZ/mzMAFakIa1L9kieyX2BPp4oh5J0KUe
IcWYz+bpSg3nC6SgGN0m26A7wnRHD1TDTZjWny5whGLT2yAkaibR+GVQeHq8lUoY
o/PQKUF6C6q9rUi58J2PproCYKxnX+ubq+ja30S4PbkEJLde8wQTx7aIRhzhiT6U
n+GECCfLd9Iyi/tN+G/IrpUzFhpGb+fiPXQdDzRezG3HOseUiISB50PHScV1ybTX
7XKhoT/0qwwLrEG/3nzy4FeQIfNe0Vo0l5g0l5d3wX9vUwvu32ESBR2gQXRb5qU5
06FIVs6gUu6zc4DO+gUTrXYaiUeIkbGWod/rNmvJRtX7f+V2qpmwvfydApttOwHR
6YQTbEU0ORfgli1vlaR9RoIqmUzQSyVY259fiMX7aBCygh7CaxlrTdAIjAjlVMU9
HvjRC7Zp+n2f+v60eLHWNqh778GRWXtYtVSjAqN++TaHW5Rm3sYHVKyOCM1gqneR
+o9JuEWhsbc/RQF0Ci3CM7313ChfAxd9We01bXU48jvxjj9/UzL9F160nIzg+6yU
XGvpcc0vIT7lmcAf3zMDLuj+6MZkQTJjupzJ4oXfXf2qG2C8CROMyOm1GsGROjs1
JrrtrDB3UB0yNqHHKfWN3d3lHTX5B3GkeFdwUQNct7lXNSo3ba5wLAj3J1bphxGI
wkMKamB8nkUU20h8qfkvToEnrDQymbO3fAb2rw5qiO3d/OYP9QYBDjWpdW53DNIb
wUw+1XVw/8UQ7RCbSephvpl2RNlJdQ/4sfIdx8VPrO88c3WY8ZANZyIaB8pVamKS
nBA64dm/TI7/jcKYM9nCmaRz5pFBpk232IULvsPeChMFcYsRO98J30e+Lzk3pHS7
+8PcAJ8nTFm643aLIQ/0YxDa7cnb+x8C2Zxp4XnDVpSB54Mup6uNyN77wZOy8sv2
1SaKayPGNkZHEKNXJaabeB1UZdLg5Ad53HwzPwL6Zw7aM3kxKPKasTzN28CygFaz
2icOcHZArsTRVfExQoyWp2+ytTL+LLjBwp/DGT04zrre9bJyUy+RBdR4h/KQAM8I
gHgPtYvWmLdfbLU2GAaE5/MlIsY87krKYmJeMfbW3eDhLjLZXRK11BFsyuFvFUXS
bHTTWoaYbpO6ZN1VCSX1QKRigO9vgWs0x/S6GtfoHbbKtYK/s90nhDAjaU7n2tWV
qOdzXisS0Amc/ecDmnDOSofNNCJzm7KKfFPJJ/gS23uUIoiR0Y/hNy5Do1b4HDd/
H01pYY/8l1LAXBU1gxL8tVk+8rwvaLKfqGW2vAi6/683fm1gwMWKMsvuiVD7URrd
cM83Nh+nu13htpmOFOifGA9SsI3OEM0D0axY7xYROiEgxFgUvDjvDub8b9IlWPdQ
3YZf+nbZS5O+xQjwrGHKmiqPUvf0l+0OpX8sEj6jGJrvaW3+FDh9KFSzbO7Lihvz
F4bw5pKVYiwI6OFwENIeqcSPnH3GamUP9No3PBFJqUUJTrCgfbCerEvDzfwyIEc9
ZP5glLrsnTFcipwKaaAlbN2iyJeCvVH9k7RnPRt463sqWuoKia1QgZZ7tS6uliuS
iLByIY1orxrARs60ZFZMaTVcfFFVKYTg6OCwGB8UmAcSg0kXxUireXtDrf81i3iI
qyiBKSNOLgm5DOK4958lLaPzBodLgY8ezhV5cPR45rKFY0EWl24zft8AOdRTTVAo
l5BnKCO33C7Y8ZdlA4r+k5QoEgN+KGUsjIXh/nHVlDhkOCE8it8igL38UflK8Omg
VU5MYbYi4Oz9ghJLos7SFcMZ6phtN3WoeKYUeAf6kYU6HD/qFoMk0C49BQe44zM4
v6+1jfBQ/tYei74HDTRoLGy/UQmM7MjjYfjjHCYuKRWXPnSToH21nNYbuiWdu4L6
4cPpNZwVgC3kHQGDkTiiVsgmQiC83nKm/y7hsH9ftx7ndTRHpjgboe6+kLBy/SRT
az4R1mYOtu6/NVrhfO7Tp628YLUl2I7gYMrxb6wrlmjJw/vOSvSJzDm54fJMLIJO
M+aESd5p9Y2+U7ouuqMt+3e8KIWq3Ni4J3/dOwi95mQeZ4oR8V3+u9BqeBRUyq20
vb4iV9FHGcoUDSzo2B0dfgtMEFA56EMgcSlqT0cp+jQw06JqpRivrC0SQiipw6CV
py/TvPY5xzQY7L0AWIYB3dGvg6Fl4pMx+m4xmvZ6ETkTCHAiQuPB+rLTV2u1A1Uz
vCuEAyulfGbcI0y9mW8Nu89m8cVjojRDkbRdJjHBTrUTPJ8mXOP9ONC+DUynz2Kv
hSUXp/uSz0UPRoK0vKw4KzJkQRGKnXpXSzwLVYrHMouzGvUKmq75UhAcwP3jQicH
I6zEiQEjqQ7UYZauCc2lgfohT4/GZ1ufuFeeYC+LFJrZ69IAt+SaOzutEbl6FRa3
62eR2A/lPJ3+hPwvnGdBxG2q9y3perYT9pp7XRb7u5irH9UjuWuAq1qRJns1GxYj
afpPQxFKxn58MJwXyOi9TRyqdvEBwvV5d2dOXJK0yVKEHIOuAs9H/tBib2zkcK7U
aJ1W4w2vK6aEw49Rq4NnlJZk7bfC3nPv+PXICkZCAkwGaeD7Ic2w5eLY1qOcqgbj
0WK4UZJl5psPgTGLEvrxwuo4Ev+oKnul8zhrbTnEXyN2LmK+2GDIkasC6UEs5S5d
a+SRSWj78pT6cg/6i5Wfb/wME6rJKr09/cAYu9YcaSqH7tEO50CZTzBS9+MvahGj
/MWMnbR5lE5LBIodfpD/JLLM5YM+pUsRgr9n91Hg/sfjy/iQ++/PXm8AeFK2N8MI
7KCo/SREHzTIWHvnkMiRP9vT7i67sbwp0ahNduzOJZfhXRjnVYSjttFI93/Srp1N
9pgO1x32eQJ1TXJvwud2oAhVoJPKNWvmhQh3XM5xXDDAkjh/+APlG8wwRPVAiLD8
xKcXhKZmxvCvXjprzE7miCAYI54jNcN4M3fTpDLbhuc4YYZP837B2ZvydCMWkzzr
0jtfgNjpAW+SBPSR2G7APsok5QDGeq9Aj9ymZZWh7PUFbQFnD63abIsNxzOorTlr
pA3fRsPugkjOdb98MqwUfrMJCWZoEuGf7Ihq5d8qdZdRKxp1AUB5ZEPoL1s0Lj5E
CSy5/q6DvEtISn/B2d+KjnYbOrrprcEZajst9Ja63BWgeOyUd0aQXmjayevNzhCI
A1FAG171MD6mW99ZIolg4KNinc7FdiVFkh+w/KnLkbIE7M+OQhH+cbs3EiHQAb7X
ewS0Jd9A+uc6PhaclN7rWTFpSnDAqkQU7ymBUH27x970eSp4cXkG4cX3ig0uFqPa
613tH3etMT5fA6degF4XEHuY2f8gx+zFW/89h26TC5ePJJgSvP8tW/92/s4c+iDz
RCtS6Y0UxSFqjTg+Ed69KbkY5oAb/vbwI6jr8HQdVGtbEt73dsrpvBLIMgLRPu+c
gPeD15Zg7yHqhspLuDTb7wr/zedLo/uxVIZ3pap5wwr1JXezWhMmi0nDhGKOgE29
8E5r/4fIleweG2ylRIOpVI6XsbpZ1bE96F4dkWMyPvZ/A6i+XFx3i5wJYKi5WkNw
Si7/y198obIoYi+a0mup8MC533GI9haXAn0086by1XRwZRDO7vrTkbLYrdr7FLFq
lhnVgFf+RESk0Gtur8+SNvupOB1F+btLA9ujwNjDYujGXfbNLE/AuAjn20xfr+XM
Svh7OHdpil58X70IxpJTsjgIJcYwB4XTRhyJ79iaE1aINe6secSjb7xtFUX/05ll
Y6xx30v5hio3hnGE8FNzNraY5YfYHX+S7mJVfJVNnKffkeSPS7qwLR4e06dpUnUC
FdQLvDICeMcHJsr3aRU4qxM8kpXcnrZNATzr8bLdXFkyzpb7qhDN0QW+XNPCiSkZ
wCHaSP7YCUArA1WBVtcvXE62snmvcURiFcP0sEC1/IEognaF5APtMOMZVIcC6yLM
3Bn+Ym+3Ur6uwbss5Fs4knsZsTLu4YrF/BOCT50cc69mfHhVl9pl92J5hn2ZPp5K
IyR+zQ0nsURAPihMqU7Y8Gv9n7Li9Uf4VnduR/2G/TSiqnUWqZMqqGpGmt2UGTKB
4PuxGbAXcb+HKHmyCh2nIcsxeVpPm8nOT+lpWbf/h1L+L7zpa6G6B/D8Rp+NhhkK
93YViIihj0+boiaLxi7eEgOr4VndOGm1KCSQULMpFKKwALVSROp7qPQ+pBjj0a/N
LUejKKBJRbdpAnueFqCd0abaUXf6ud+l4Ganuss4R9aW6BHc3GRD7cncYnqESX7f
TZIIt3oUX60teGUBKSaQjAGZgWvbFBZiWzhHdIMonyZvagBa77sRdKkN/Ddx4xlH
l8ukPmchQ2qQPDqRslu/rxZsNisZZEtxQFu/jR9kC1DnT7VnpqQMrFkogB7KguNk
MOLWx59Xv2zVIuXrNZHssue3ht6z07JAFtdTUrgowZ/kMC7/FJDs+GQPtoywwg4y
csmk7tlSnguVT10LE8GYbWKczonAn5P/MyI7owpbsvGM+6t2Sj99ahonod7PboW2
ttU1rtqEbOKEOPGFvjGhrA2RkBq/fJpisMMJxJ+PREoDM/a1dlT1BfB0/50JhAot
jhFW2fRZqXQDKQ2u7yFqJdmDW/RclnEKA14RUVjwBpyXFlmsiCaoNeqnbA9F3KAi
w63spSyREj+SV+Q8QOqMPPdf7mQs9sV6DTGeozi8uorJuWgYbBzI6j5W4V+8vbcN
IrEG2zyXUXt6m+6v0XJVYjBqlo0bkfWjOUDc8JYtvm43DpoxwZopLbBVxqRI8CSo
cW5q5bRy+D29pbAF0zS2MWYB+LA6cK86++UKRKE1fNwCITW5BxLYYfbEVUHg/gt6
gA0vIE500irlXghvTY6GeGFd4oS5/sjftE7i/9lQQN/zqC6B33Y34hSDmABF9j5X
4I+UAp45zDm8Vc2dAHuywXr9z/5c/Wi54sLll/TTT3rKx9I3Cf3P4olCMIXgdw5I
aOB8FkAPz+dyGg17s1vXibPDf6zb9rBC1MwD5DEDorDnTSL19YegfKVO8xDyLSPr
dysyo7xVGFny456tBdC2LAg5nm+Cs8lDSTb555krR+jYeMnQSFOdRGJbceMcrTkf
PFKbzlaMz/WHNZ60spHLmfnVhA1kcrTBuQ3h2HcTBJ44qUaEl16Kz5bDqUdLtEor
xrnlAFhxaE7nwWGF3M9ifUYY0T41p1eXmgIQT2Bp6jDlVcIEBEdzlI/qECsc2eN5
lAeb3eh5fcj2FMmyULxBpy8U/qSCz1uyUkhqG2bawlLxC8T6HTmoQdtPlrsk7rbg
lr5G+r9Bjx5irbkcEol2RXUadMG4KLJa9HSr2hbTOI9uekTIvbQqJV/uOwdGfRks
yzAMBmWRM1m6LhbvlfxlEhqk9kBYhBt5ZNt+tDl28al9Xf1ROEE6cJJfUDaFPy2h
U0kReJu5hpzI8vdNOea4hShZeoMB5Q4qrLMHREHO4R3E8VMRIVDYkhFzufVxWlIr
pQa/Ck8ykUScU8SfucxHocEdqtjhul0VQd7QZeZoKL3v4Vd6teqFlst1+sXPhMJB
FzmNelXlu4kvQzLYkxQSy/Pwf0OgvAqN1Q5ZlkFynWNRLCBnOJ8J1lxkjI+zeSxh
lgJufDr+i0+dr52RZ/5GdA84C5vmrvdQniyDHqNOx/aR3kQ7/2pjm2hMaJMl9jjy
7xjwWQtZ7CR79JFM7ECeYJT+VwwsekbcBd+9TlPe1IsITIRbFqlR9JEAMscv+K/8
EINhkIwscqKElePCdZyxRX5XhDfAl42+qNrb/QkJgUg4IAsNIWsx7EGq/kcs5qUR
oc1kqU6zauFC/19OVS3vvd130FSbIMT+gmXGhyE3ES48ONbB5pmYbOsTibWnMUH4
UotoUvmiIFnYNVM7yH3M31TaFhUrVMGgAeV19mh8099zKqrgOaF/pI/FzluyEeYE
+pc5DddMOi5H+KbdX797l/CvKsoLmslU5FnlmVtZ1c5QhyNdictBhlt66o6wu9mW
5hnLe6WXcg3FF1PbPHRJ5VsciF7q0XnvrzgPQV6aN8nEgCiTZ1eAy4dkhSEpxpKW
v0TXdWDh/Z37RFsFm0nfGj66DpygFbKGr2Rc5H5FS8u8XsKKqQSpBYAT0YhwiY9F
n3iSW4kISwjWhkafYPnfXrbRZ+d8CkY0D1+X7ue2vf3DfkfUwycY3sRWgim0L8ya
JUzzYYHfaLLbwQS5R9CyQQMlX6rrWeuKWnGzZLgZrRCbZmXtevntWfkhM1pPpZC1
+s3T9nB54QYq3JFjfiJV8nmO/hs6WWQPD+jMUwEr949Cxy+PfGlFKi0PKS9kgsCx
MgYtGWZblrFbdSylgm5ENC+E/yh52VJtsP9bkG9089q8IEBHuyui2x0CTi4ZyGPD
bvVNpftEMF9TYS6xETsIG6VccWZiQu1bo8xPnLc8qxQ033QILuDKLStG5C6hBAtY
7QOQrN+0GUZpSTcEJOMHMmxr/2DbkuBNQs4hQOdQ4GsmGI3hdM9aPUPnLoB8SCZi
hgDBJP4KW3AouL1QWrYsTAHPqmEJJ41DYFRl4eAQk9zr240ElZ1MmNc53xXj2bBW
h/UFKTDDW5NyXwCuP+VMCHhptsQsA0/lc33U8DYlGPk74RRikKyjFy8UKvWg2F6A
JIWbzpGAULIGBHf5Kh2SKTnTGV66O55MN/73TGbeWZDv240yPDFcXKDZZWHrblpA
/9vFX6g0axv+7rAJI6OuSEQ+myqPz7sLXQZ/s90AkokI1qynxJXy7/mFNzmCVdI6
1eOld8OqDDWBG+gzRD+eS5M4fLO1WacNtoovbsGW0JliBF/vwPaopBnPbX+u2KuT
BPORMB6MWLKptTjQLrhSnctl4blG4JuISnge/1CYQy7XNfB0/+vZGZNcEnPdvdZh
pxV1pQRFKqykrgMBoZf+NtAGK/2pVfigI9bZu1FVqAkLo3Xb6vwIe09jJOFeuXCu
RPpbJBcfRN28wiYLSxi1Qp/K78sQcdbD70kogDbMSoc1xoalyo4qGqaKth2hjIJT
8CSkuElJCY/u5o4hYTzUmAcAxjpn1IQ7PS7jErf772S9F7vLDOjjrWK/3OBVi0y8
n4d7tGSKs0WKb1fyo6W8zi/xf1myDM2WRovbg+v0+LFtoVKFURZCxpB8H0c6tfwU
2pJ0KZr7GA/VrgChAT803PnJxpK/kUMTtN3eawxmf80L35itWpB/eT4XXqRVTw62
rYblD343fIknYfeQIneNPjGtfjXfZdBaExZtQuGS147wdkcxTgGyvtV15bXxOoPf
igExzqfXCbJyY5iLm8eXGXKE7QbI/noWB0Auz2LcPTHz2beKWqsVLxKrFMkzXp1W
E293AIZdcx16ioEnVG/3diSXGPai4NLOsGcTNAOvEAn7DXaTY/UPWlh2x0vGYk8S
iEsqxVpAh5DYJrdZTuTlU83rgsfgGiUGEtYeY2jmGPzqZ5b1CR/jMH3/Q/wn81gE
oeJvHKGa2sQc6q0tCFvgWOsxzWSkv3MP9km7o9Ow8x1epboJndyzFTXK+kmfYmoP
8fpncoe4yPa3Fr9x1337WJONlsNiXwtUWOuYxDtbu7wbTyQ7e7LKW0+AT29DwyQ3
+uhBjoARrnLyfzSC3OcreWQ+9Juv4GJuho06Uhz6mQI20NUN/PWFh2OXgR3sKOr9
e6BIhASWlV/fVxubDN49DhBHWs8Puti1euhqnU0ZuCyQ2vcPs9NJwI5ZbAcvp39I
6ibwdxTfVirVfa2HUjfLQM60o0MIvYKcOVOBeMRp574odvZ9tA3WKroX1Pu+FWCh
xdt3M/Huj/Dr3m6+3raCmKyfncoHqjfsXizr9JmnNdszkay7yH7bVVop6D8qtgvU
J93dT5XcI+4pvR7d0xYIE9JHsHMUbKjZ9uFbVuupBx5TCTwPr0gq/pTbUN1+pFtY
pUyHsgWJFC1psDQvcacV1+hfK+5Du0ntlc+TISBSiwU9FgFaJY+vzfBuHtt/N0JC
QXNzhsBzTSBphj68Yedy0Sppxu/ojbm+XU16sDYJ4UghX/JB+7/nC+IvW0PIUhiQ
UKCBwu54je5+67VqC6xKSunRwNEtE7vU234OemBjOKSH0FdMV8+z8KpnyHalBgCT
96f7WU1p4jzxDxkF3dd9Ogmud696AnkolPXMH8w14G/JHB6sjLULTO2S5+0OMPdz
+w+2p4lOWH9yR8fNJbuFDRqIjkM0sY5/lZHDKyuJk5Tu1ZuqbhXnWdR/QHinZ7Wx
mbao8gQMMR/K2GAjJ1sCLanjphEnTBkwknPMTlRJS7tk9PXRsf9W7gNzKm7IJ4NT
1BPC75iZUZI96JS8MvdIAgmdLdFCA2n80vwcugdtDh3O/EV0A68WDOnqavzrUrCU
r8N6lihqm9Yh1WSE32T0DjMdGGEBlFv616JVSd4hCgGzX90u9szC7qDg34ljlfdt
63ykhKeirxXvF18/zUZVooAqENPrFh7w+LjwIIMHtUy578UIoscb8OIm7+cjpjL+
y6xqk1n3Zz6h3prNmk87csTt5393QgrtAkzB+0uUj1eDm+4Zm2DLcg8FZqoNTAuK
tz0GX1nLW0YyanvkIag1o6z2TRuRj2rKRA1IJlNqDArh3X03iZzttKYwMgL7Ij0O
/2A5d+clPGi2yDaI+9MykJY1Fhd/cp21dtR2dFCCSfEmjyiqh+wF4emhfPMoKMre
CDA1Me2YLJIlvoT3hmQWhcXdFzAPJGtj6DDpJKIEML+G7IgPvzh/B6MQwGsH4IOq
p5hsHQjItltk7S7WEx2E2P+RJWooHnsphD+nUlvkwnWcei3iJmhm8N1T/Wxvmsct
XVde3zCPlyS/I0QVgNyUVM6kpXEpo6bT2mgGiJuUWF3XnbikvS9oCHXLqseNFWG3
wHIxDJmjTZmZx2Wi30G8Vcna50tYx8yptxX6pQviLXM4Nl+JG3CvTph6BjN7CEZG
fpeqbR1LhkMj5teUUMJ0K/PxIGwG6eFVYVBiDieEijWZTF1eepnWOXiZdoEwLlJc
Wajn4RZOFcF/nf59SRojqTYZdYDdnqcwIHGZDYp4tmszBMkm0BUNUVb7cjJntZcw
zIiY2xuhaEbd+k/QfOTB3YCirKvsA++rzJ4bL7UMWPNY8W36/x3mZ1SormH//7tr
rFSP3Y9RBpBPWQYvTQSbObu10PR7LUSRT2IL+vuAyAE96u1W3t4I/0lI+Ele81FP
VUa4xBcGv1g7wH1oMDDk2WqzKQ/+eaGrGPpZrsjh/QYSAQng4lywG0AdWuLPb3hP
gUmOjKGx8riu7J/Sg74YpGrZMSivgsvMtTNTfHm/gwZVhbG22lWT25CFgnnzZ7CF
K3XIj/yQFdm+m0ng4Rr9GePVu5n5rY6mb4hRkPNhHZ7UsbFFmMcPmfRpsxbel5eM
JIZz3VnVXGsWGRP8zhJ8I29yy3xQIPQHgHKi/BCUE+/fCnQZ5zzyaVIap/A0cImA
uebQPWc8l3QKiifjGzbo5Ho545FGF4soZBbgaq3Ikk1bp5bf7na3Tb8c4J/ESGC8
NNhLKGGBTgf/LHR8UW7udxo/EitUI+2wLbGZU0qhKoOUnf7lwgNINd/GCr8JgTkm
taKKavAcSNgsNYuKDwiS5ULaQ68zL1fkVxAl8rATvjQEdHpmbZPwOUkubKWZbFmx
esY7U96VYaLKpNlfgtiDaLviAHpikgGatY9vNAo7vujeb+aAA9J29UfJiBjHkfy7
7gDoUTbWDjfI5rnbMXzpTDMVU+Te4nYsz200A6p5mWyUALXrJa/tX+xj286G4pqb
yNfv2HeHADm+TN7TTO6MXR6LN/GR8zuqb7r2K4lqgrstjPwgJPlQCXL9+Jqb0Jyo
aMihqcS9iFz9TL77Xgx/8kK1riiKU2R+Iu2blMekQToTxuyqp0gJR1Oe4vyhr7Xd
QLwMaZtYLj7rNBRfBVs3iSWJ3sBMc8uLI9vDfHjmAZXbtD79mHh0GlPVqpV5xeJK
GEkMkZSLnOedTfMlwnXxs6j0FxtufdIX/MCv8+RKFwMC2ShNXFH/yRoW2wVDWzqZ
eIfL3slqv1W9ltSoDNFjwLQaxWg7xeo7rSpMCdoKF7WpMa8u3//ZugHLNvBZ0eov
UwWKs68szTC9OxgCMc7sxMSCMaKZoWkGQPL7aCGUfFZT0CEpVmqli6MzzP2Z41B7
SISRyl5bRxZY3SsI1qDHhIgxXslrxHOpCdLsr/STiJPhjgMre1VfgdsPlruUN/G5
nEjyafiQ5ZWsdQwuYd+gI9wVsf7Lc/j/ASSPoJEG6BRiG2jujify40xIaqGZYSzl
F7EFWaGyUvQY9h5cFXBawZVD+zrhnn73eJNHKml9piIJ6aVrozg9glN4tn5PUVA9
QSepwTWM+Q+/HtE8M49xO19mIu8BboxQdCgCu8ggaV+WlvbE+60sK5KDC5pz5eWk
UuwbVuzvlEQnJNifkQMaiGQJQMBJOpmPoPISkxZQf26ZC/g3TPF3FxUR8AextnoV
nEKO1Ew12kCwMR5e7KHmxbj5EnShF+cM1HdMQMlLYb1e/LnsH2gx6vpN9RBScmct
6tPyMDtGslyXHbLR/ze57EHg10lV8fKg7QfwdwSf1pAaBaZfJjfYpXZmIVLG39DX
OVZz/Lw3K2rMSdVZpItg/OueTzjrZtv4GCxNfLYeWoo/AztCY2QiAtpY+wq3x0J5
u3tNeTv/xkSMSK9iEOOC8gQxI0miD7Txl/E2HPQfQGPFHBBlQ/fJ+pZo6s0KbvPt
lIvToLlNOjbHNXPTgARYtFjM0IV0pEdO0kM/+lOHHUMWnmvJdtIqrMwfaLtINGcb
X4zjsDyhKjoYo7D1bciuaaNtaKj18lcWSfq62Su5TMftyrD6EhKV+7VdLECmDgSG
YGZoMgjRPQQv1qowTUVejbp4TfIsAJC4327B4znaLW+YdBUdT8O72XGWa9lH98FI
WL8Arn5SlpqDDzIPzS5yyAbtZ0GiWv8OLgt6SD+Xv/WPMMdPYEAdtohmNrQuteP1
oLDbfweLS3ZQMW4/nD1vt2MbxJ0AEPIFs3eNbl2PE/51gBra4x+2QMvbQy6qHquX
eEwcT3EW3bqXoAmhldWX3ncsjnXCbEug/TyXD6TwFZhI/euUdBoEj2Y5xkSUHk5i
oKl0Hs6LWiXcRgMdi0EMludo0OEmFqpdFkrvdEqKe07t8seuCmicQu1zKMrbqJEw
XyCHTpK0yS1LzfniHNXdiwxDVxZbHI6YgK+cFyOa66JsONSRa01ALGla/ixQZxS5
dE2D4u1xPHeQYlsesRm424bOwwFfejfZO5mUSLHjnHmVQ9L4tx8Srrg94WIVpd7N
f9SQmkmPQxCZfuNFHy16wmCp6OtLJ9IiCzIQVBoMYILO+4x3gIA6xldULTvu8OOr
TACQehHiTODclkZf1gIqbI9d6ukQ99s3TU1hrHfHJI/KCKq9gKgGX9zU4nbtdFqa
AU08Pt+D9mSNRCRXrZpLaZqCz6rWzbwylt+iRcGl5fexQalGqlWMLy8TTotoh5ML
2Rz7CK00k6YeIFLrFo2+1Zl1TGtjMebvse0Y36tS69zifU+8GnxCBtOJnDAGdz3m
2phpCUlZwMfXigOEjchFL1VRt9oSH8OlAf9iOLfgIYB0lVE69YaxfwySOA+nIZIO
jFBOmRyNwM09np0inNWsQBCFfyp+3RkLTv8SstfuJ7FCR5QSJtCkYz7dWVKUoPSJ
ZDX//vSStYZ8ZAHUHNDs283Kuy/1Z4pQGyFcBql3bKX0/5q7IRwmsvvvafbhBLmK
bPR8d/eleKu76MED9YsEfxRLHHFgeKYStojhgxmSo05FMHsTNnQathFa3IHRY8YG
nO9E1tOcXAegsw2RJo38ECSwZ+pM09BgCWmbZX7rVOj3h11T7Rr3o5lKlQ9EFLsa
/mDwIFx1c0oRzGPOLu+0e2Xqt5oCi11b6RSssOIsyyGc/VRuzJ9zVd2KsofTeN2X
+77x8BCM/mWHo3XedzeKiJgFoM1gN9fgqVwZrM/yfhG66zbDaLpNfmBp/Aza1B6H
DTZOUdMT261XyBbwgQuT6KHsaJXu7OYdizXWkKILL7Gtp9L2nGnEEuGWkc/pWfUD
wtOOejAZYc2BgB21k6FXNJRLiVAnLxlLCrA2ZdI41cwkviHAoQbbNtRpc0z8cxGU
aRCGrU8PJ/Pvt+1mS5Ogz9Se3zfRXaOIQ2pfbqnyrqyEbF0B1/SazqexXaPiZB/o
dYIRoFqr8Q6XgMLalcJ2vurcybOuy/y+jCLPW9zCxQYlUa5sd8Gb1IZnCqu5YA1o
5mkoC7BhN3k8w5IyDoDXc2uHOsjNJJiaBbzHOsDDOaEWcXyqMfXlea151qJqCmSs
9KM3jOiEU5x7ivMG+UPql/p6qjpyGeA4kh6ZaXaddjxXWUmteh2EhiX9E2iaGRQ+
7zHPpX8YANRHP0x/jcWetEN5we3RQrKUgCmQqu+VNBcTmztTNzQa4ZG4YF8nI7xY
AcmZ+sz/S8Yr2bca6lwzcOZg1gzKTGxEzpV+4yo3+nNOcQwWCAK81zWBeEWqvDhI
Lz0PG03WnLvM/8w6A3i+kpUZLMMOf0PGBHeRuXOJXTcEj3PCV3R/7pnFxUolnbwz
xDeY1Q2OTmuylcG54v7snvcJNPsIbKeLDWv4TCKLrpnLBwCWIrEYx1+LbsCiBEgm
umaWYCzBTKNx/0JsLvz6ps54idsiJbkmZ0PM3ReIMJfiY9GstEaQc66n4g2bSC5C
KdxilUw9NfDz5TZ31Z6pOQoUmS8GL/20adQc+lwCot4SGDm9S9JmSrvDQJkgPoqK
Iqj1EjXV4oA/pvvCoz5zzJN6vsfQKz0uTaIhkKKhugsuO23U+ns0kjbXVnLCy5p1
tpTL40OqmtV3KM3kVGDMh5s0XIW09fk/d3ybcHIz3qFMyoPlSDtU4zOxgLXFbpup
ix8N0ultco6A4zErwyQPK5uOInxta2qtl6j4WDD84x8ygeg/QA3OPx6ugjCKT2/R
4qSbpfgKMblt/ZBlAgl3RlwLaQHKoEkwDemgW5v16ZMnjRe+bdbwz+8VtPFskq4+
tFuex6txqhfuA8yJ+WcBqF4nuDSaOjf7EgbihoFWiJS2FlFj8dSiLJXb0MmCTm6m
Vrw/rk0mBZ8btkq+4ld4CGs7h3tMRaz9pp9JVV1QrrW7aQBnouOQZVdd1/oRTA68
CbO1BDzmwz1zi0uN9KiUqXOocZyHTChnOAFIfbiKYQ3B/MaSSTCEsMSDk6aQNgRT
MoelLU6hw+A82m6oyde75IXFl8OaXz2X2Zlz98xVkKJs3sGI/C1pKKgGhqhzk3y/
97PXn1e8ukrscZkmt0fZd4AbvCPPMaojdg1EqjkpLoVpusKX3mp/nguYGnLZw/W9
Qwthu3bxRnj40TqdhGLqJsE1RAUmuVTkXorBGpTntxLm9OQaq7l2PH7iLUetH92f
PPGuYnjMWae9ff34PwvYrdzdnEJFuU1oDAuXeWAAEQ6BxM/oaN8j/wk3btiqsmcE
iO97msvpR0veWEQFh0pfe14xE/xL9O+/M3dw7hEVCjKZJbcTLk1v1WQzDeM4yu34
hDybpM2d35FZ9QkB2JAtwdN/TD2+eU8QVxe/meaNBLAOgKkln3kWb2y2j5/HdfFO
OmF8Bw0WOHv+eTZO5SB58wWGBlFr4yV02ztKnZ3YL095J+t/KVGXx40JD2P5A/dj
UeCsNyGjkSEXF5ZJgb2jXkL3cg6Ox45eB0+Xqa8D0QqmdJjYR9SXmqc0se85RTIf
3ehZNjAKOaBSa6zqNPp6qJy+VaegeNGfGwcyphNll7BCVnzB2hckAJ4KxX2XyCKB
J8Jbqxbk0pub/f7fMSJJiyogSGnYx+YaxPxn0PvPmM61Rm95zpXc6697ruve3jY0
ftLLAF3rAncK0qsr3ijxA/ge5BXUlV3wBgwzdlV/VztR24MDfowMh8cEgUmlmJSF
AinaMdpwqqPxdQi7BeXho9RlI7iSGvpDjoFQS/J7ib4LflCkxu6O3ykNiRqi37Dx
oGNAUxv1OWJKl+q+jITaCqhy7HWFn9I+CECE7RrcMbVs6qNN+GdRWEInLs2p2Xk3
ru2ajF3XQqFEdw5J8ucYp2TB3BFLHe3hHWDkr4+VM0tqHBBoFM8cYHU0RVPS0P6s
UB+8RVzHdkA9L5bs7dT79ijjELBqIwTQeqBkWW+de7jqYWXnpBd6c/5YBdgREE0B
+aLZORYojXJ75fDUkLVUmcAuwCkAXFfkU0wbQX6id+rUkwJEXBx33XMkPJEAR+XM
RlUyNV/fFZ5jRxk1wvuDoqtlE4uGuMdDCWnurc5pPHPFT/1qll6gQjKmWHKj8Wjo
sXWQ4Pb+No4pDxDhtnoWumW4uSfDBZ/kHQIs9/zAD/sHToS7zSoF1Kxr+i/aikEA
hH908HgMM2db3SH0oxb5Pn46S95vmfcGTIZ0wlTA3aZ3s/Z80RTolyICsQtqHLvp
WMnZZAkFD8DTLdCBqKf+TVkfnfgfAURD3tzpXRErKIrGon08EJOB+PNcKmWAz6Ze
stFmFmJ0IcPOyBqrBzBev/BrHYa/VMvCpTfntlb/mPq/A/GC0ldcaAZuoVW+1pyp
7imbTJ8Ymm34Lc29FgtCdBtpTfhjK12huQALXTQ3EcTcIOEwBuW+3X0E6O7fiOVY
1NbAzMh0X5ICf3iWz/+XUqxxoQbrSlrK3On7xJrGsA50Ov51hmm4c+fbxDhafHgx
HQVvSia15xYZpTyj33qoTNVeXFfXunGxsSqI0T/C/85ISv0sXLplEuCZR+WBYb39
n4w1i7xVkEKIGrQluna+/iilnAdihJR73t0ZnoeTuAQZvS89xyd53Nhrf82+WBqo
8vm43W1q6sCv5kWi5SG7D9MnnheV718fh0PsfY+dZtCyMR5Rpn5bS50/GPlwlMSY
60mW4ciRfs4jF3y0dPE5cLhoLwkhTL1U/a6s3b+fVD4KFPEsL/PmGQ9xZajDFCxW
ujYlwTl315Z5msjVGhdDNxVzQT4J2azgtZpJSTUimaWYjTZWJMFDW+HNtrJX9Kfc
hyYksRWK9Ng0vO6QW+I7cSS8+DRivWJrfXbtmASzjbW5PYNHnnBfbVbYkFVK4JIz
adM8fUkhnKBsK7N4s3Kbbx6efgoHou0u1oh/cqbMEX3amXwMKMLtjKYNzT1LAAJc
pY6s0S7+Y807Zk/benATiMASJuzeIv4zHnYktscBanCrlAQIbEX0GWeSb7Y988wc
E4b0jLvxyMUcPrcpuqvr/HnK5nWV7OxNoddJZf4dr1suq4mMENuZeOp1evBDFgWC
ZFGRM8EiSCD0skJglbIEh4vsYcTmPY10Y0Lf5+okGgz8xCBOPHA3w+lCftCAXubm
Wukr2gTe/codHoQfShxyceojGNzKRv0wTOS3NXpBYo+IJ1phvv7bFx8WpaKyPQjJ
cPk/khUAXHWUuDcF8+6LBpfUovFi39qpIFU//WI0pNeZ/ZeYL/4Yq4dOmJeDlOK8
mJIxFEz/9zHmLvwMAQPERUfDELBYnccnbqXVjN4bef7HtRPpymVESzuF277XJE5U
gJDbNBxBeOtRPeQQZBzpEm+spFK3QwDzgrtqC0Hu5wAF6QHkKgE3SYFM7zyknbE1
gVi+BtbQGhD72kvWd84uuj74//uRSfZfc5WNmqkfspUE5rw4yU93ZO0lWyVWRj7X
+gfkZ1ZIiu191d7/Cb6H1mnViL4drQJZNxwuO6PY8va/zS9amwFDYXo/jp5IizHh
bebL2WHFBr5fNZTD6Qhp5h73wU/RRLR4uSHcKYmkG2t7DvLwev3BmdQxIujq1yh7
OUGMjzx4dbvnoyBWrKWowLsEFrwjF9DGp/2kOlpcrC8hAv9wkuTSzkjxXaKt9aX7
rNcvoIKQWUjNBfUjfOvDFzU3T+hcrKbFguCECtSnlNM//rSb4GFfT3HacrYvz0xh
z7qx6QwfM1z/xjFzibW3s1jEPU/VSz+gVkDFrPtw66JpDtCukY7tTqgI/ZTxg2si
W1F0UIpVROr+47V7x2gbN9bREBqWod8I4fc9klBiZ1S7zbaX5zHBV14kt721VQq5
55M/Q6QEdi9l6ulOMUMw/JMziMSWisPyBFwJhFkBAfVfpTIy1lv0Xo5fofWER/4W
QznWq5GrA/6HYxOP7QPe4tsEIkCz7LxsFk2ObbzQcq2EfdFaGQFg3V87IQaBpgHu
UDy4lBCQutOcyO3BmBRThnBUoX2x+8MP9tDsf6SK1pnbCNwv2vUjOq+SaBlrlRhf
/j4LH7Lff9w03ntZT4pwQ+6SMsLaYnLeyylSFakaCjUP7Rd84qch/v8Ngj/9JqJE
oWzFi4HHkFWf2kaE1sZ2d0tmRvcZpFhMdMbRFHjGt2RcTZqqgVDRJuIadF2OW9By
u/5fgitxTFFWbCXoime9NAXJr7gGmuso+DyG0Wo4h+5gZbPCTfj7+4fBOph5DKiP
OyRHx++oPIoIZGu5k9RP1SD8djVlhw1LKVsHpkMxV4B4HEXSf1Sa5yJhpN96ZqOr
ObyTufv2Wx8pNdH68rCSPz6rdtLxg12Eaj94tpQIrUaeM3IDI/kBJsnnpLzgMdEK
qoI5UR0XTxyCo2v0QhpIdgHQ7HB4ec/9I2vpna6XR9iAjGhXadALwqynSeb5OxyX
FDeLwAPia2hzCdf5LNsMOXmajzV2daUMjfY6ug4PYdBwORUF1jqZCnSUP+yTicC4
vxhLQKCeBv20VoQU5nFfczRGnb7ebwO3Y44YciTbpUfqUb2bPAdGstKYar8EuqF3
jDr6uzeGTs4oZuhi8RW9sMz7uMXndzTWAKcpFSyEbsiCHHQXBXlsyKccZx1OM4Dv
ZZiu4Gg62oNKdWmlHCCSKoQXQ54AH9TKWwZRdVdsU3u4Arwdt3m3y6Ly0q7ssbYu
lnJ5mi3OtexuwE2OXzKwm33bfPkZgooImuDN+h9Qv8XD8kjI3LjDkNga5aB8rw/b
iiZysh/soYRlDEF2zbtejywuBpaKJIUfDsbYZEg85GqM+y+mfrWa4xfya/UtNM6O
t14OIqZD5+oh5FjSs3c7QuswDBz6FQNyMzu3WeaFibl1/zEwt6Rk7BaYLVMfeS6t
XvOb4LAmFTYWjBOWgZoEJxDeHEs9q1WbqNwppqtNt9cbjspQE41QJmXU2BknnPTh
KwayGWukrnG/K2QUw00JYXxbwNwkGUtAYXht8Ns36ucYpDyd64ci3CdKSuBuhaZ4
SpyCV8P9oi3HvP6NjS9758biuLZGBeg3oFeN0CeIvFv5wBKrd1gc2Njja1yHrv2t
HyVavIXNXrGaVxxH+GyOwZERwCIwMax3jKBvi2FL/T8i9dSxylDYjWWMFp3cOnwJ
FVjd3fwDxO4jIif6v9fcK29OXO1Q4SOR1Vre9b7I6Sc/n2PeuJtojK9oZbtXoTg5
N/WG55G5Qy9m94bzc3qemcN8prgowNc8pGWi+h6FJsu9UrTwy3/tYd1RMpor0L5z
glyYNTLFp8Gtm4fDRvhxBtsOXG6TNKlXeKWNVF2WVQJX+wtOxNjGrRcdbhZyYe9a
3ugQnrtCc+ZoEXcCIigTTxmZ6mReNVeMfrQTyZN4SihUklFyEynMC/m9lyQayQtG
6yw+FyRNNwxCzMF4vT80VtMvjGn6Dy0e0zqm7Hi1yAS/NHGggYWs0IDYfxzUzfhQ
M6bu+V91org2aSuvgxfOYhkQeOloou2iaeTBdPyPCl6mgyxTEnkeqfk5+FH1l/uE
eOuOKjDHEai4m60ux3/NduWei2m4kyQeeeTJj8I8LHzDOn9uo50YTcdHD+NxpewY
3pLX1Wj03/frkY2XhWUwItCvZpibTbET68mHTJytc64qXDDQ0FgQSv0x9qZwVfwB
OHvQUhQS218uTwAD2xgTJqNhmvP5+Is8U9uEsbCR7th6ozHD7QM8tLDLslTL0gti
ofNMYpNC0P/DcNdcPuyDk35qxWn7CtSws4omO1YqK6Q1PUf9dBMqN2XU2co4/OWz
LGZiWsUVeO478Qk8m3uy3R9rrpEzKZrEzYjTIEY/8tswWgNNWIrMddPJrZu53WH6
xcbkQATb+pWykBQdqQm+v7wPX9t4o3olnKAFCgb5ogqkm+xe+i1cLIvUyC56yj4B
/TK5mHZL8uTqd2q+Dl6sEI5y7svKo5nZPbsvwK7BtQG6rWDxNbYj5c1XNDa8NZts
YN7lhW3wEMBHjAjA+FQ6EEKexaJtV3XmLMIDIbSyvotOMvZAXqqHEo9WYeaR8R+5
6HoU7z5lbXmOAJbgSw7DL4x2Xpm8Co/37n6joJj1T4Qo+ETtPFLvdh7VSrcpaiqv
5NjYfTD/A7zNu7whkFr6pZxtxo1UmBjSiSkaJ2Qdwcs/f5D2N7y1XmWWENCCsQqN
8WHE2eGHvP71l8M5tgbH8QQivXwGCmbO/Ar8SelcRqaw94CabbtnvhiW3fMWkUsd
oEPdBau14444D1wzNO84SYgVyhUKdx2kMFgFSpipa8cCbx3A5bM4jnboxHOgyUwo
JnfYePH12553i0WN2d2qB/uqfcUcWbj2NKrqadZUhCrsLevd3+fMiNoRDzueLhGl
VRnU1N/FaqHtXl5juvK6H9COGbYCryEY0SI/dkQ1bmbd9EYIwFMNSdMjg8j93T71
pLi+xbMbxxsSSr7EIR9UCBQYq5S6SVAJLY0ETihDpHN475iBFQ6hTZOFs2fSeLLz
SqjENpASk5QdjzPS6+I6GSi5aHg8Zpklmek12eEuQ+KvPArDckub6vvwpqcCEdug
dkwMd712JIRKSrV5B4A2yF+D7Pnl4ehC850V5OBuFE0iCuh4IAld7f5pilWx/Ypq
yFHN2OHWuwRv0xpsu9gwqxpwfxLUTcp6Tshw/epWRJIPWfZYX6WxedwUwtkGcAgS
Ki0rlRxagle7YrTGKJfmg7nwJlyy1z4ZjkEjoD3hhNUBWZemBO0N08zGqfUhvhmC
2shWIckfu8SaioIFLpWb4zMTusY5S8uTyNTooKy1Jc8VMiNKxLPGpNHxFDeCUcGN
6UoPTr83C2fLQvd++j72i4HR2s3P+uUqZYQmbSNOvH8vHnsnyRcKG4VT8cUb+y+R
hXYTy5vtvalWzbpqUs19FqPVh1UWCGwSE1f8eGoKkBUMmqr0r+vwce8enH+iZAU4
LxlBP+TNRbvuF64HQLC5lw6PmPF19FYfEBTDXrnc7+ne9cVEXRamMKW0aNY8i+5t
ODkP28rZ5B6pT+FIuOkGYa8No1hqSFmUQOEqDzBebkrtxOYxvfxwSu0M6JhgNTuY
1ym6RdaYrtict5VVp1fuC5WAAXiZVRHAhBOHmb92pmw+WBOBF0tiNR+ZyLHC+upE
rXXDDUG7Y6llLYipqXxtYrytIA+oz4np2k0twKsiW7Jyi8Tgnimi9+RfZS6PSE7M
Oj3g0NCpT0IFDXr59O/itvK5uSdK6bX5Kv3erBk9qOPzdgBRD3LYsm0fNzjmMaV2
ZddN8JMvemjYHw9UVwjuZiGf3+8b2tIcRgu75Kb8TTnRllUs11MHlKx3e7Pw/a7/
q/UA0EVAbZ4TUFAann7WOj8xd/LztIQ96MqsHgzSmaBFnj/leFvz3do9/Z6CGzST
rmDl/SMkERGcnb54psLMReSNesbWXDjw4HrfqZ1cc2u/7teBx4e7PHuqMVpOiu0D
T1By33yxdBwLDQ02Rr3IUpiDj89OVGpeOl1H3P6tC6OiAbysEQdCQJjn0kVY+i4+
ozsEwQp8kGsKeH7MSfNDDmvLovwRGDUh1r+7Ns1Raop66EivnTPMKMqImhFn+Y+w
Y8Z8FMRBLvG1ZsUxD+hNy9Q2d5OIY9QQaH5CLbG83K6IK6+drGN4TpKQjZMuDFB3
oMl/U1hViDhpH6QuAatPy0F0aCW1UIZY+s0tyowLbeb0KgqaN1JQC5SlAMRbmflN
FlkZlnWEROtFS833A0J5tDWNfzNAsdSnxc8loJib/Ceg7tqtEnmnHMsNx4Ck0frY
Sb+9sBU8V73QM7SVllhdbGNuxI2uPBMWQafhIHhDrGRzXLtqkZ8ryjP8WMYiBnOo
TGPPmrGBG4AX9wa3enByZXhOyVDRjDnYc3n/450MC0zP/6y4hN+iC3I6RYRHLxo1
S0kiqlrO8HPqem1lo7EE3WXthsc3VAQTtBK3nrvjq3MwHXNhEzH9pPzgHh8EMrSE
yyVAEuui79vPjOodGaHsZa6dCLwsyVRc8F2svkDOfTHW9XS5BP+Mica3DZ+Xof4S
A6p15L8pw9/qRRDIcqjJndDhhpoHzO+D1zNMZQ60X/RemvDLMj1kbsAiVDRIWu9B
oyrpWUCkOpIDUXJ5gDvKxrtJZ+JL96PdZVO7hL1Cw/efxvmQUr4cZyWGiNmslW2I
3XzucHrFacu2B7ZLrnFtKyRPUrfj4GcA1AaJq9aVKpXhsHN7tlhbJiWMsdJDbtzR
75tubCOBVujaNAbbh2w5ovZu99/vXY7t5k8HUsvW3xsohBKwxAtIKPa2kTgBoQuP
az300h55ALrGBZ+gwCAMJT6wfoILo2f1aa/T89c98p7+qSFM9aMpy9HESJpkhiB3
lYkWMAZtKu3DTfgGhgwnwt+byzaf1yRA003PXOmAeSi04Qvmm3Jxo/IjM26cXOOr
M63i/K6uIxI5JHXc1rvEI7bXqYDyZ6qclxF5WNFSNR4DIIJ5y4Segkmp1+1sZKXs
P9p8btaBshz7D5tK/FfYPqAixqmEuPrIZTtv7IZjGcVFfD5aQzk0fqPse72NQf/P
ErfeO7fXbe/S2mVyXy7R5a5D8GbZISPD5PnytCICga2LOaitWC6W6mH75oWzt3Bo
zxyVJwu2KMakr4TDx/qagUgGMRQ7xJ5Za3T50vgQTNSfmHDRrcG/gdO7uUUiV0PU
H2Z/IjsIqyQr1IoTggGp0tzD0wTXLuTy3lqWuGQLRXcUakhTNOeLJoouCDjYMRAC
VHxo4kKAN+cjZHIQcxWkBKaOoV1yDf+FR+8NQdd6Imb3gDwXEFmZaglVUu/BPjL/
zqgBsPriRfH76lf4i+m3slhO0zZrJo5zLECYrHW0UweyrZS98b/WlbonQ14Hu8LJ
PXYrqEVx1MpyrzNzLdT/luWd0XwTQHGKRQ3slCzhZT9t7XgFNh0DeVfeee6L0TG6
wCC9KtCJAefHzdI6RcAfAdU7g9Hs8hjtHDtWaYYT+pafsqfyI0wDxFKolZWOwxiV
vUBpVXdOOH5EB2sQxRwMkVgZDMwID1GTxpUMd5dCmkLQV7FZ4hbh627F4P2B0Yq5
W3KUWfX7NPVXXl/m7M5GmEMy5zgH7+LKXp7ttZpm8s459Ngfelg36kYWkaPtN7kA
kvHYcGlXnXjx+KVtmYp75G/X2fq+0ekIezL4l39s4Ivis0jQC3puiCa5q/ThSPYQ
1EFHEo/vU5/z0xU+M1dFjbYcbBJ13bjCp4HCr/heHvs2jlFtxqivggBB+QoTLsQi
2RZt9clytyjofVC+bOUQ+6e8k4ylHxX4rT7cs5zjAvpG/H1fJz2JA4W4D8L0FQRs
YY1f+QkCIvPK9gsaiKbGdx1PabDex9K/D/X4uDZxku2dQ5jzJngpTCE/EkdQr4g4
FdJ0lPvMF17YRk6cEPsKyA6t1Y1h/MzMsi0Ul/5TaqfZb41jfR1N1zH0YtTG84kf
Waj7hG+CpFIkNM3R3d9IE5xnf6M+xuR+Hi6O6g9v+RwlNKVT9Y1NIkaPdnkRM7Sx
KcX5Wk6gmMZa8XNeQB48PV4lBMFmdRIQ6mrdIPM6yUt4HeHGRJf+rQ9PtpG+8oBd
PiK1AXGV8CA6RnEYcj/+QHJ6u1PDeUirQQDcLIJttPM1WhqUgKyQtiGV2LuV0lLW
q09TO1j80MbEaITt8xxATSZjyuLhh1vbBMbRSoyHqNwTLo5gG0moUVNdVjJmLqwa
h3h5QolKAUSzFz7wBsB3G8XVOWMi8Jgq43eDz7JHw/83WpuYcA4t5fS09X6r1oCZ
w0AXzu5eASnKCMdh5AMqXUMWvraRKbZISyJymeGLhmhwe7pz++dXq7BgSAcWx9SK
K61rm6yUw0B5egvfmfjVoljIHzPSz0W/nOOSYU8fwl+C/YmNzbkHLMHnY5IH6VSJ
o9WOYE1Xd5wPHsjaXHmwhxq3JW2yJoFUPhBNrqo4CRLIXg8nYeKbS7dYTyqIRlEk
k8YUYYdfQRK1DLVlw7IuWxLtPCfzanZt/kNqpfbgRrSPB4BOEuXMhh/mgY7spcxA
oefoO4ltWLpe9L4tL7Zdy0IYxmbO4gUc2cbFJ6hghB2X7XVr0js1s7QEjeFTYyep
X8/vv4ePKDJPEuXfw4p2N46nQYUYqOnwa7jmIY7xjsuMUbAKhfsI9c2A72Rngo0N
VfggWZHyVrSXg8BWQntBSbHB0Nx26yO+XhLnHyEmmzoQgarHw8xvIBp8tzHywFu5
oiWXXhHZ/mkNBqcBsjhuEpbrtIaqpN40yda5KQWhS/70JMdCvZhEv8dg8bnhU+i6
qCa5AbcqYPYJwS/DPrGU/kLJUZKy3+doXTFkSf93TusuONWmeLoUFVgnfmlQFjqo
Z5hV2uePbeCLKDf6kD3xCnZ6zWJvjpomTWNOmdhQUK4sgE2Y+3gE6omzxC+395py
FbS0NnhEkgO0+4UrRq7U/Q1XtotDrj4e++CG7tTTz1OblTPYVIIUmG1BIdPglSEG
+hBWDyQKowfYx4hYB1S3yEWPcgtAt7ZK3XRgMFNqVI05wF3IccymIh9LMoQ7Fhod
82G6qVKlytkQV1RKk0ePyzBERZde5s/C83Nt9LWQWIFjVf6URo7DacKv9muwng46
DN9yP3FJmNbtu58j16fZ5sr3S8FDj9bAaYBrWUl6vV+aJ68QQC0T4W7VjosWaAAJ
I9u++eUe9J3NPu2HEK5YfEgYIDKeVc4y92BLX+Gu5mSWl7iFrixgGQ0nKBGj4s1E
x1pnM583TBYYFKZFtVeFeN2Gu4pJszS9NZsM9ts9EyxYUjHoZjSQkQ1exCt7nC+c
zq1nJcDtnTRGpCyodxzmB8EEy7q/SRbmL/KcXCKKWBTsy2pYFuVkT87cVpZ/fj+7
3v1FB4kCYoKlOk6BQCpSQiMSgj52le6aPzvfAFLtwWgtJlb3Hqx5n4J7mwYgNXWX
k5fX2AFa7MNr/JAJZOftCgQyi94j9YGJqc68rCT1NfLTxktMST4c5Y7f1auxyRTk
8INbZo2ZqolXceYvbb+WOf8nzIZ3xCSoAPjVoOdWB51Fdue/g5YhVa1xHAxIQqcH
QzJcM/hRxu/sJzs8qWgkLdi/ulwux9yNb3sLSEHADOaLmULWQJC5uBZfKf275eW0
JMdvHrBJZz9/J67cl46fwN7NeSl9xFAHkvGUUPHRZfZnERA+KakP7608inYIo80T
tfoSGw/RuB8Osr5Ex2QZ625H2nDJu+SNMfh2m90i+l2Wmf69iOQrTN5ckK/bW+gD
ad8EkteHsGOIh6pWlaAkmXHDxwofkbhVsSmiORr2yO8e4hRrDiLKcNR+7Nmhfj9Y
bxNqD+xy6OAnO/I2g1vZijZuzch1GnRPML10CFM4rUAsxfzXeT+dMGShKWgw23Dn
GBQKpkGrK11H2lDudzGPAXBnXKGlBM9UmedBW4hfoR+OZF8tkfqGjNKbmKHhuCQD
N4/Vaq/luvAJs7YiMJJQaA6DLBIQirYlodyOFpwdP6CTFJjhIUlc+3R2nttl5VCQ
j8I6wAPgzn3gXNq2ObhtANfvRnTNDbb0yaVa2QYG6dJRX2UZGKPuMAcj92dBkyDN
bsC3JnHC3tUwpFf6RSE+ICpuMt0lFtQgutXiFXeUmrsKfr/jpF3GnEpU38K2XeeG
mbjslBYevN2IkYvWtnP3R8QoL7E5MtIIOkJadi+fuAXgmU2ffDFynRizInpVdUvo
P7XZPuP8m7e6THELJKxy2DZbkc/APOdr600nt/CMFhqUngVOqfDYIkyDOTpbfCeW
EEm80h6eKmRlYSaR6nxksl7M7WIA+ug9mFonawZNoC1ssBQUWQLJPWxtLLd6YIgD
1Oed+5dLEZJMgG1sfekNRg4rBDdblCRmU8aclMZ6HTBN75KuXdIP63wOLgM4oiVi
FMun0Ft1I8wkRdja0487VcBaipcEpg88+A0R5a7PEJuDnm4xVinmrmnA6Z0p342f
bjPaf1t+Fu+v7HrsNxuo7qm6qRlgTbzJJ9DV+Rcf/ZCDU6XhdML3xE+U3xXF/rFN
foFQEWXteAJHlLFEisqO8hQlVGJVTKB2XG0PEZ4TdGcJ5pWhkumyH4bCkeh7zLmu
L23EPl3fjMNtAx7silGqrREIN5OII2MdeDQawoAEo82Q7VUKQomV+GIdVc535/gS
pmwN7cJ8fK4e6k1diHMeDO/T8V7SPSKPeRS+rhyqU88z+3s6D1vMlAjwO2S9ETY4
3AysIIr4PHX0RK0DyR1i7GPcwHeWroN50MmgooNlReHpefhHD4I5ljXAEfO+hca6
MKoGPa6+/MUWMe7IudJBiMbxikzIroQoRY+b/IbXi7IBDZG6Hny1C5K8vWsiOe5X
VUFS1D/9wtAAiNTEOWFaOUG6+Hs+jJibfWbLEFOH7+Vzzv7A9jVCUlJgTI2Rw24u
khB8mQhx6N7KTNU5cxFpBxLa8XNfxYsjQ/BSkMXGX0/VNlOmMOSwRQoFMBQNBn71
XhN3TPIHK/hdhkqyMeZ56trBeYyOrhfDjOpSrbGd4/rOQM8seV10XpPa4vt7bKn4
6iUbMhHAb166tCymVPZCfpvShRAIAwmt4IihpacQ3vLbL3sz62npfh7Yy4m+dphD
S086NdPzLYkFsV9Ei6iKyru1GT+mLpz6UH/g1ut0piRMI+fJ9JTESB5D6V7h0Aoz
sIpMan3CVf41/V3wx+b8Y/e7bZ2oUo5WxnHokUQevL/XDPIZt0Abh1Jw6Q8Zwzxe
4nkXxBL25KVlJM+dvygDoQv/+vlnZujz4Hus5RqtfLodinwd4xH0Ziqsufl0EXWV
+8LKU9urSxRkPcQOKfklssVsoKhU2a2g3l2TOS3woKWkGZQ8N8fsRXEinq5IFAh2
Xw2dIOG9x0jpQBuDXXLajNTyaxvLYPFFqNv3OUvXuD8rKvLm13dHLtcIX2GQK+ei
CVV0AWu+usSaJYsQTwRw2tdx4CKEeWT48I+B9veSZpTsS6ekA3pDuGhXgLMoq9lt
d8S3yr55tOcrnG+HHQOBGgUOMPmjdE964h6t1j2Zkr76LQVtlEz5zSpgG1jlUH+z
Prg9mq4pivfGbzRZVy1VDOE5ZiNP//d1KXcKj0rbJ4OOAT7FthkHa6AHlQyLLryI
fswDt+OIHmzC0gOyAwOCjoIEgqj0pmleqI5ASZ4BjM7zoKcMNJa+yR2bm+PruI2f
gNPLT+NwivBF/7pR4nOj/g/X8b3XzdPqjr7GOK/kJgzn6I8BTtXMyAXY6uyOMxsW
QRfFti/cLsxI+oalRJl7XyCmQ0NIU+EPzvep5c8lzc5gmnPXm/L7iYWQpxclcXBK
DZwUwB7RO7C6lV9zXNDuWoHnnSIjfBCyRcmS6NABc94GYGC5MVIU+DX2p55iwSHp
G0YcqQlkfFp4qBjqyK6SCoFCo5njFXQqgfx7vSt5S0puqfdYlBDLfO2VEqi+fGdH
cTWVryxOI4IJXdPX3tzxGrqzzJfanGAnJd7E6Mf/WAaLLbL4fwOL4je4uxna8C4i
O6NpkmVIDiXtCEzQnG+oLgL10dPdzau4wyiIvfkhK7sSy0yNefiN6cT8feB4HCsv
ubuNiYsTr5lcumIQcGTl5IwdnN9c3ymDLmAKQLiShDTmUV39ufW5ec7R129LPAl5
SCbuvsFB2MxT3R9seOVCtaGKV19T+9hFcFvD+0mnPYSnP0MhsjEJWb6o/8+VtP5U
26Zbsyfg0bbZ/Cs5QDcZpSNBzj2P0NybDAVjSf4WM08BHnIJBJTAhwvZByLZvnG7
+fSOxwZM2IfWMtTRYTlvJQhQav/YllidS+CRoD7LMfEMYM+s0N0oh4yHCQxpbzWs
etcdCTOO/stVCqt8Sbt+ScKkdKQp+LZbJk5rHr9WabTG9loL32wRR0XLP+qJJS/g
o3VDbyvaXeE69Sy2wk3QDDACDjw3vhdtjtezKKQG5sSsJWv9n4pednXGErRihEUy
zeTCWPaUzVxEXw54eYEfZiNeWA+0O1mNgyP+118xzLTzwLONkhtqMwD1e7NhNjCd
uV42wVvp1sSbiJXRmqhiCGXnyUH0ZQdj64r8ST5oaBiVjlhwm1/Y8R6wX9uDtrDO
B4gnJLIWk+x04WZg8jYm8Bx7Pvf6+COjXpSI4/C+Qr/ZO2eb70908rlOZB1flXpI
QA7FEMQjj9HYeDGKGLhPgjxx411iZTbLOuWSIKaO9srAyvI2D39TNzOwQhRYy9aS
Kakp+P7iY4Nx4MTohGuips8cid4E18Z98kTrIRuhS64lz6D/uS5j2vE23SrSatqB
WfgVxct+LpKPyrEOL38hwG4NgMhe7oxLfT1VtR4pZicZeD9ynB2yGCYM69NbLaU2
rXS5g25HRNFbLLdzIA20n7MqvjiJy0Se42iSIGInLuUslG66nAxJ4jTr8G/rFE/c
I8n1bfMktKo5gAOtiFMqtq1wYUXqnKPDd5RdwC7sja1EWcVZHVfmk6aRcmVKH3aV
hJIPrRP7C7suuqLkxuvk8vsILQ71HLiMwrQf583cRT54zR9xy/yn8d2eg42uMhu8
jI6J4YypqpkDoUUgN/MV55jO8OQzxthe73JwIQKeFv837Nd6i6Kw0tDFywKzIWBK
FXzcHbzDeGoh1H+oGpD0J3doGa4yq2DqahgsIHAr9CL/UtxbNb4T0ZOh8CounrV9
xHVqc0J5IZvNOlnELnbWiOSMcE/gMM2ButNkQA5LomT73c3k+xpbpMqbh5g5SprN
lZvBuKrEBSolh0tASBJ2zvBQVH9y8zT3SeaoTB43XXgR0UyAeEtPUCvqzEF5LOzh
tCLDwv3k7L+m8XiV6aMXsc/y8zrqYmwhdYwBGEWSiaDXETMafJ9SAyg43bMsQqLp
FeMiEamFpqnKwM+7uBSHJ/sPJH5OWdyVXFjxAVswL3VvfPdLBWetUTH6k21jLfCr
bBEDYrLJpWWSSchfyumvNelBRTR+MeEgPDENsY21yzskgpLP8XzPfzUj0oGePP02
pBl0pgu31WmrIwCjMzf0Vjt0ZiHXURd2XEOM1lpSsrBTH6k1DTBp4G6A6YVxJ+VS
OrXFwpQX3kAOIyRXa9oGazCi+vx2Y27jyfJoQxy3gx7LHQ17RLatbL02yPpPPjUY
kyi3q9zUN2laK1WEZMLOH05ybhzl3XalyUL9P59Nq2WlH7dEeEPRlTHrwZaCla/F
9BMja/0OWMvypuKY2oNVAbjAexw6+KwWDit3bwZfch6RjEMwLn1INeObr0huJAno
EGJp7CO6OIo88USq78AhXUEP5+BRaWNfohbh+E+Y1+z4YmappKpedC/N1GXsqLMd
gaMgxK+RrP0/PzUB7WAXHshKeVn5hwbOjZ17T0Ynet7V8dlylFICUf4RDmGfEpem
Hgjo71I06kys5kIaznxoXveoQRfTzxmJnnGEwTEY4aAdOs/uIYLFIqcV94Z0CVdS
7imu9Q1e2tBhqE74tn8UHWATTXDkjV8CtYOyo0GRxuiBM519wk8imFZr0QN0dgop
zMPqlVm9BNWVpLsbBWEAai8ZlRkja3Dw5I6fCowLzKnsKqRyUEstEcrLG3RKYifa
zZ5+/Kq9tWXl35oBipRI077D5Pn8Jr4R887rge7LSrD7gaeZtsD+qxrTIfnvXHWE
Cy2GpZ3BI8tn5BWHvQNCr8k3UNP1VXSh+Q6lXnUc+ywmtrphetaZkBsGfB81cirS
lqFHDAHgjc4lGvtYzmwl/evQ+eELpQmc3RC/6XNVjKhH+JRiY42bFg4ouqcb2wNP
JJO1OKlwz1r0sDXysPhrESHsJHWDPPygvOQOI7bTtdtAVll9axjmU+EvSce3M118
mnsg0vTQxesbA4ENwOBWrGkalykIwH0qGj053SDhxmCrR0m2ODlWvmrs/cT5oyyR
iQqxmPNbepd+n4TpjN5GdreUkZE2+EQXuBMdQomeW8r7ACM/m1wjWSapgbOqOEgb
BEES5I9jYrrHoLBMAXYigEaOyUVhIA8Mmb4Co+N//u4argkBB83EqRJrcjIG9UK3
3/k4esOcR/Sa0Ev2eVus04hZX8w97TJsCt3t3cZJR3l9AMX9VolSSWsjOYtRC9iM
pKWnkLWfNdEEa69MpmLqXiQehNG7gShvTKq9xKI+fxb/qnbGd4Y48duFKTLcPiWS
bLgweEozQb6qrhtiM4Gg3/bjT4Do+MZdjOmKDIe9+8QiL68i/Y7mIw+k2AbE+qgC
3qc2XkE2sIE0+gnGCipihu26CVeSvbweZVhIYuo4/QFHC7OJh5Mg4ng9PpLgBh3E
zTASj6X/Fi7UsyM6z4OLfKJnE0urT9IZWTdY/5SHHcEBtEwkhwDla+u5BEZs1LQv
gURnlchG9epsUxbP+Hce78fPzJv7gFT3XJVVPCufsEvHiEyqy425Ki6G4wKGixC3
hPCDGka2HoaPvGw9bgFDbgGLGdQZ7N5Nc0G4F+4J/vKBfc0XnWV8YV5EDTALCfjL
Iw1HgZrcgy2FbBC7NC+BRFLE6nZ9xwRJWj2BkGg+YbX5JEsg0LxBS90VU7S63tWI
edIN5Z6cUV4WJDn2J9rXShz3rRGbp2IN+V16OI/Uyrm8QlIFPcBwShVPHGd3HnJ2
9GLlFxCrTt5UnbeRfFVBK8G1mXJ/H4YNUw1QOV9wMhQPnhj//1J7Hl3Ug1UYxJcE
YOdaQaKirazE/CgIAzWYdKO1rt7dhUkk47d+ZTBEzIX5+ZyZUSTJK3/EoxU+hufR
d3ggpi+iDJ7rZ0TfJ3TBW6/uwfjVQTJn8jfBA/T7uR7sCjrqk4+JPV17zzugNTpe
nPB+jCohZMjh6Tnr2xK3EebCaqwNpuyRj4fnW2oiMnsGPgwLTmVQ9Z4eMdd1kjPf
y+Y0YYNGfUdBIuhpcKq7wnrZrqABQEotdNUzyuh7NbiHDalW55D7fhYCsXAlBnk7
rXlMGF48rWsFiiUO2YTD1ZrWVu1Q5VA2HIeM6M1xFJbz5An28JtbjI6g3d6YVYeO
i6GQRqS0+BxyaN1PED+DZbWAIILFQdknl0f+Fl/6xXij5q4/alNZEaFoyTT2wQCE
lcSzbWlR3ranGjw71QHGor2k+//yhuqktcv3S12rgwCQKgxT4ClBvocBJodlcevg
S9gUsAetHfWc9Mj577kaCeovhB9/wkS4Ajjp7It2LzSsk+QK0bA5ac6iZjpMRQDD
GnHt0exlrMhvB1fE12MoeWZwPK2w3rA0rqptlw3V7T913wHgGQxbAS8EMCUaZYHN
xP3MmmOZXxNfY0tx8r9pb8rwEV5RhDSFF9BqEZypKY48f3D2u2n0LMN7RavNshQV
redLLD6v+S7swDbbztHpXrCD8bavexgKyc+V7NXYjbFgUPFV5ECTA2/HpMuYdWbg
zVBGEc6DUNylxBLxnGjt7ns6M9ONhhZ6iZzZOuwO2gppMTJlmkDPI5QELil96rR+
IG2LO0u+fyVEFFtFlNdApL65riCT6K1grSJjNRnaNfyyUwoao7QBSLBeGs0NtBmQ
+SPpcx6l98DZc6o/WeOXCY/0CvZAAEe9YQJi0Ty2SaUyCXPIxA95kP8wyjb7LuCT
6NuHlJQUYxCc9NGhrP4h7XbqXqn2ZB3rxOuFD6Lg/YJspNzbnulBb98le3GZ2hg4
iN5YeyJYDX28tuhOIYyNhDDC2KIb7V7gzagEAuB73Z39FI+8c2goSmbT1/PANEdI
QpGyOrDCoegAiRhTN7/K7mtpm7+mxAD/eW7mUokawO1R5+cni+s0U4gcUbGTefO/
w3czKb9ioFT2LHCs3eVWiUuekomhZqugTONdgsmRA9Q7KufHmj5NZdMZSOkxglZb
W93QJCD5Bg5Lywh6PttaqwrpSbb147LcbCg6LWFOTXuBJHgRUknZMTAT9a2VQxyX
026UjnzJsa0C29DwpOiX2IaCa2M+DcQx0yVLM1UMbFP0ND2ESx036t7uuQUwO2Dv
y2qWDZbSvJS2Z9Hl4OumuC7CD7n3cMH0Oh+mhHOAMdP1Na3VXMCdX3BZm7nu0AK9
YpiV9UkE0DQjYQf+B+ZjgNzn221DRq6H2Sy20bPxMH9XJ1ReQ1pTqOj2RJ+H81+l
5eNhPITCV7/EwwxKBMDoI9U66RClY3tcSLU1ec2HibOrzCMqiLczdXYkjfjLnBgz
h877Fgw+5IC4g1JHv3q2yVMomaNA4GHR6KFfIdyoZFP/p3azKfhwotd507114Ei4
ET2fh+Trz8xN2VK84FFbqO/TzuhIFL7kLDVjWx223GtjujeVDJnkM6Tdw6sc9HUZ
rhw5EzEvSwkYu01FlW49MpLcn0nghZ+NIeMoPnbqwlyMvIg7nQMM8yJQIrXvAFA9
0iNsMo6mw3GemcoQVDvTWFMoeLAznqNgEdVpA03y+r6vf/t0LSLhDuxSDrp4M59O
Hzf7t7bzTfH7b6cy5CjpegaGqk6F9myIndYmSzevqwHDP98UKEC8bN3JsgD4Pgk0
nuvQTdiwnpfkiyNgeTxUBO09O25m7TpcBeqNKgHxz7gN6yz+imoCHAascXLAqd9n
pvRGdIv/YNaEv7ADstBzFOwWUaRKDXAtR4fq29Te5o7A/hjZB49FCE4tomYp2sde
/kB8mx70xZAkoa28YPYcIbi3GIvc7wQKYqkjzxNLMPfept2gsqT1nNfPLFxk8AC3
sGsXqzk2XKbL0z3aU+zzWC28g7cS1fSAeCm1/xfaWoPbMTnNsmAwjBpRr5TVsNUr
PkMNzEIXlMMICxkWBLzBZZM7jPclZCuoARywHhCL80sZ72ku3xHjB/zBQuCbJC5O
ivYCq8bWPyFR9nnbkv8RqaKUVQDu2ned4e2mthYDGFY0qtzIAgSMDm0ZDp5v0jIn
V9ahIRIuyIgRlm+jiHm7OYq5c4/A91j/9Vyc2veJ32MCtXlkKYqd+oXgrAYBflWV
bRcnzY8ZWky0NIgatwjy0FzP97/OgQznnLXq1kF1at/ssCdZGN7jK2rEURQUZgtm
CD8tCsK/wT2QV6banG/+zkLzVZPbpJsaDeqAlsr4p9g6Rx8sJHU9hEEnKzDJ603l
E0zBKDZaw8Oc/wYP2RN5V7QrbOo60oaAc/7nyXw0bYDRUCznXXO3Bvc0qFeXq/is
aTUCcge3NmiUY5hEyGoBJuI35jAn3ikbkNPjpKxZgy1t6XYi7OgKdomsF43o53+F
r4TsSlLONGTlWifh0kyCNSFluXHJuifKYAAdHnEeMlP3g01MsEq/fOWck0v4djd2
MLIHol1UEBiA1P4/0+/thEEFFi7B8+Iq9/JB198/oUuMJ9/egGeMbgsgon8DKQgQ
Nu9qHXzLU9O78wJGX/v+4mib3n5GquqB7yfOrewIagcYSZpElYFJCOhoQIpudZEK
ek6F4W906LFierKAqDTIdqLerPgfTV2qWgRNq8r7RCevQVLaYWy9ovntTyqJ6Urr
4r8OKmguA/JO3tnyjeDbnLeTF/RT9BGqM11ZvPki5YY9LXkX5yTJcPqRym4/c2K0
N+MyxSkbo7eIv4S9csF2zyxhkZbe8gT3N4YgS9JHJFvqKuuw1r3lb2UitOS3VEVi
MY+k8VT0TXbw0rXeHXH2fM6WOQN43AMcJGCoKkv/vIS9wgqrn0oE+GVuWaLulJL3
CiW1iz+xwufqHUmfMR+doYXG+3oeJTQ8ailTBwcgHJAx374ZevWbuHceK5KVmBX/
M0JFUH1vuTqFybdVKW+AKUvHSb9tPKfo9RihCGm+MadWGDJ9pVEZ8YTeNhA2Acs8
BIbCgYtEfD6miSJXUs5jjNboVz2m/e9zG4zEComxkGksGKwL+xBwNzaBE84fM0MM
IP3k4t2+gYyFte8AF11urxOGqNzPqdk0//F+y3qvLUjbiAhNWTIUJvCs6KOrVE5/
BtDVjZBqbaWAH7uFieMReaL/9HWoV6aBIkKXZR+rkrP2UDbPsRFaqtrJCV5nsuzj
0eJYamckdwbFu6jFkTEw4YpO/kx4lwDS8qk4k2tARc+eMORFrGzTJ9ZSVNAzoiN0
MnBtQx5OXKlPZfE2rWyGn+rCqIB58JyhePc+NDYM4DRYV6JjKbQ3r41Rozpxy0t8
iRoHGp2yOSW0zheQmmu7oVgH1plwy/3o6Gmm3R+PnM4P2HKcn5wT/aUCOxrhGcnN
oyLRQTfRNUFz4gRF4QnLMdr0TCCxS+uo1iFHtmyht/2kaYE2o+8lYBnmpyYTyDSh
ueLPSHR6nfZTzPiy+VRtv9le6boo3aSkgRBoORgs7A2jX+x3mGwtTMhlkm+i6ekM
gzJSH+vgsIeIg4ObiJ12mLwkqfbEc7VScIPCSn/9W4dzgTwEhHnkJFgRSOxjhBhw
NoCyMg8Jf1leF9auHglSIO2AQvzXWCUKvBnQlFkpkytzBqSriFu4C2A7CVJ6mApL
a8Vj+iPjttmIhGYwmK+CuZhKg+4kBt+QzeQ+n3j9gubf3ZCJE8i/JqSvpcJbYK03
sn4QKw2YZ8Bqxg3G5IX1aYCunTc8QAAF37yIMzhAWxd31LxODk3Gk/B/KhUzt/yR
CE34EttxWfVYtrYes9IcyAZpSdAS05TEw2a2jtglSXMIAeN7qiQILLRGUR6DVgEh
Rcao328RClQQVO/yEfupL47+dVp97pwPQJzugqiY392GgsPjzGg6Y5yZTdv4Vm0b
8abEBp5l62X5GIWAjf1jDgYU0zV00A89/ofYf/6tiE+euerRS2v6QiyZWg0xCfPf
ifTR2ZpJ/NqqnHr0DmHoW+74QlNRo/gwgxSMWmR43hZqRPd6twzmY/nNEeYcbU5z
tQaN3rc3p9qJaLvXEvHmUaL3Wls55BX/fxI6kpVO9vf5jMSQSpxTrEOvshDHAHbB
vxtCLnFyyqmsjRugRuEUAnqYddkOu62qU3QYzQjs6H9vAkPPbfn0RIgi36NmhgS/
7WKNARYzdcYWDU8FrSCwJgYRh1gAEyq9KBWdx+/tiobEExeCN8sTgu0WIibuJi2I
YM4B/bScbmDhZnUpxtUBtoteKUGwd0aLsbh9Uch7HncRcelFHV/DuN9CylESJx5L
L1VFP/x+NRc/3vHpRUGvzNy08f4yKEWZNvck/lyCSsT4zkvOBS+wviqF4jZ7f5ui
9jKbFc7d2aqajluVrIew6zxUiWQLesdneZ8KuUCkwiZB5oRwLr6Cz2u3GyxHwGm4
O2xQMag6yxkOK/wl3asXGokngRgNegqU3kYPQj82hHeDmCjuKmLpnytCHcEG/c3J
tUWGNjCydbKh/XdSPml5BE8uhdvzXHWH+oF6HAPtjlL0ijim6JpGvmuZAnZyjeqC
z22PIyt1OgReC0SOsTsxBn4NAP66sPiTOfZoC6Lt2l+UjIjFZePc3lJmlPOrsyWP
lEUIoxU/DZ5LWwK+foGHgWerqKbZqKnzQPBH9rUCmIQE6801pRNujXaSa3rsubvc
kUlhBiyyZjffCVlyL3RQb6t9mN7WOabqabWM7SIW24d8AZOLl20bSrz7vhba/est
ik9A7AiX+Gl1hDd6IF9mQJZplMIk12qanjwfYp0mT7h2ZbcS1psAejrOm5zOTovj
7+6BZK9pSth3nlYZ9agqGfex9AmO7AGRNtpSiE6igbgwpxAONpG9nJRKCerlad0T
BZOSJIdsIpgvQ/2ff4IrX/aC1wfm5r3DNzvIFUL1GgemIEkDfBrKZUGbm6/csPn8
fR/0ao4aSMWXYA7j7lJ5Jdv63VoxTzyQKuEv0mO2rpAd7sVfbbu8ugY2BRwBkFy/
1JTZnXaL3xSqkL5dayyFeSVWyCCSWiRbSFCGsqE3QcnGGN/9Zv82EMtiVeWta0Gb
WCcfWFs+SmT4fhCkJuiPY4zJIPw4eHv0J3Tfc6VgNTPpdqlVCoxLWzW2qAyzPglw
nsI1oNz0BVGdadA/Ly3HRLB/Oaq/G7+DoJvSBHvVegsokVlsU0lxxO6J1UIarehg
ga0UugHYzjoqecAWRDEJg65Zv9YPKicQFNaL7Ulbz9PWIfQ/kKSDwqJVzctRFsSA
AT+UIk+qePdyN0dGySQePH7teXtr8aRLtW/Ewn98vklVp1azaA+OPKMnNv39IC9l
V0dMC7VubNTTIa4ZF4ssiSCVVE/Z4JKPyutddQ2E5ssgkjR5aaa7e65gAKJj5OpA
tpytJO7AK4+BGt+J2aiQHcgBa5/2nkpOkjlp2HfW8318N4e29jTYU13YghYbtSwU
SDwQ+X0nJ/FOZVzPVy8IeYhC5ZXnCAdDUCxBUmJMWXkZIzPk38L1QIMXqlyAsi42
TTNA5TNnlpYBNOg0QZ9ZyZ4EgwxLugV9ts+YQiobPnLYi9xVgC/7FZOu59JRw/Li
ofOIoyMJB/nW1wLove+UTW66Xxu0g77kGV4RdzyqT/kZeLLaO3xAxUAWfyqDGOyw
a9AO4PoApPuNOrCtiQTW5CPVhzo01Ntg/3OPTnMljeKG9LKjEE6hvEPGSmgea+sp
2K6VnLbb7RtRtVEj/oz/9/pUJcu7JfNhdOaRRtf2vABVQrsHbSJEpY7DxROQvzWr
OM0sX1MSJpuHA/qX5APQY7ORqbr137kWl4S7zA3QxPv9JjucWDC4AJwRiOLcZISI
iDrErr2ikW551xkh0my1BC2GP7sVSKJC6rrvG665RIl3x+Z+EFRXLQS96PZOfZN9
0HCqAyAGZkRp0aYUTxKOgeMbymhpET/0VKXus4EFxLQhfrdQaZQu9iUYV4d6I3BS
b2SnDfh0WQuZO0l6JER/hjSEB/hFg5NXqq5RsM7TsbdQycuwkJz9GpmoBanGdA61
En18ku7H6/T3sb1NixEkj6ZzNFEDHhs8fkm4fXuLRRZplh446/B5hdVMdhxf2rYh
MiR2PhN3RXwQRjLswV7MEwWPWY4GFEH4Vfz5ZwB+NPLkpIFAzTJ9SZ+2+faKHjIy
QkklgqFsb4BOx4Gp8FW0gog4VeeR4D/VWHohuVi3J+eInnW1LMyQAJk4f8TaDFhz
tVK3j6fFlW+6nOmWdgRIY1swsJo9DDx0MyoOLPuTzFVTjSngVxvr3q6mRgR401zt
8s3qnaKOl5WEISAHrS97Ma55nS/6Oixlq9mC7KvAgOc9sD6SwhKt1uwoNa2IZaCk
Hkyf03zuYbUl5hmnp61iz/uY4gJCSsWC2SU+pjddx3REbKHNj+CP2G5pKDhXFdea
flsAreHsO+ZdHHHiLoT44AWLNfSDS+ZABByyz2sEV32pgwSHCCFRHb4PVe6dIP+A
XCz377bCFoA9AmFob3IgqnPtSIKMsyyXcmbzSg3xRPLubxeTi5LRgsenWRLATt3s
67CSEaOuxLWxOtd/tsrsdawnF7duUSIXh71r9Difa24xSUtTOYSSeuniljhNAIz2
9fdd+dvlm8XwTvpM65t1/EeutgL2oISLeSmQR87Xg6MGx3wjZP1yuOBsN7yJ8J2Q
9KwKwRBwsBEM/SjKsPV5eqJFk1FKk7gskgMsk10pUkSTrT5OupWGJHlmld0A1Xsh
TDmzu8ZBwK4g4DYXWN8rnx9QCV7frD8kl0pmFSa4x+a1t7/FmrBRSV+qaYvxT4Fj
iazwGVGz/qWbsBbFUJQEpXQliqVt1liqp+JJmAXJGhVpPq/+B6mRO+Cp/sXU8n+J
XL1fJAhkPB6QYaAy7Lnmav26qY7aY1szbeMLwSoTiSjjximQMCoK4VRKI8dXGI/T
wDvA9ZTtk6wp2sCgR3/WUPWnAzfcj6AxDfPuOYU4XpZNsO1V/NNBKXVZREMXldbR
J0iZ0FixtLqMItOv/nfRHG3MgBCoTGG2EtUOHBGc3eUoF5/S+rgjUb85G1VbFur4
cWoymWqPmjW5D4w/iYxFFF/WRTVNk8jCF82b0QAfHXeg9N9EgkFdrfSbi4vhwweY
lCGBeqTHzOEzpl2ggpVw4rNXvEZS2N5yk60OcSru1zfLlBZn2FVKm24UvWpSkT9T
JmYbRMeZIwl+MHtVmWRqCBKTlBDExggy2bPXTMX5OIDiXg3rrPvp1eQOOfiVQAkm
og+eosRngjg8ZKMevE1JRwIK6eychcjDJdiO4Yf36NZPlHoJZ0Uuw7/fCXf8R3nC
oGdEN+l4F2OpDSULDVZpCGLBYvVALfoCZKAfH8VkZy0N+2ESOvqLVVGXqk+IbTz+
/w2AVnTpcWCeDFFuT7JyqeRhK34iUHKxfgMWKpAH/3GRJu8kCSoxbYwSi1I1/ai1
UDJqEt4wvKffkbpmUPxDEJCrGEEHFeB2FI/sqqzo+e4Gs08ZSHIR93F83rRzsiWk
NO2nbX4neb+VbZ0BcvhbtIkvQ/BicsE267/Pcv5+6CSD+//xL+0v6nrhA7s7ReHj
tYvNTQWjv3vjLePiJURzCVVQuxGascW0ZaFsh0reMFjgO0ZzfNLeylGQG5VeGNFI
/BDmCFstv93uv7wXSg5AcLmoPLFOTtrkVLjduqs3Ix8Gx0DmOJ87UkA9fp0AG1/a
G4eb0xgsoVa0WCSAPcisIfYE5/Mr31FXRanffP7LfsId7EWnVFdgDWM5WctdS/8x
UmGcYnpZ/1vc36A3b2MiIZW8dinZgm1RwW8bILvj1JjEP2jzR/TdoQtlXVpcLUR2
qtABM5rDfHFu/vw5Xu4j5aNQ1sGUWCTEEujMniyH0ZKeJITde2AQgyim0OK6kfX9
fyIXFjGLSbr4klj4lVI7fTVN3voCjbGv9jMksQlOfaeID8g8VzEVBXLTfhU0sAW/
MBeQLzAxK7ZrgqAKyOz8jStmDDmCkKd+ZR9XhApXB3X3UM6CTIGO9Ol4pQfmlwSv
t2Ae6REw4CTMJL8ACa0dXX6sWKdacZ8p00tC+BFRLEfQkUxzHdrjQYDQVKKlWq7y
osvqIIJW+L4JdvxyDMpNkEfk82imrHTmlfU5cMgfjRw7BrRkWAzGL5jEweBdSJAI
H/LiSmCo2T4UmohfSiHHyMLBPTLYel+uzRE06jYMkp1zgv0RzUjmNeTu8aWKExN+
9yC8zszZgkNOiqcZGbVVQ6wc77ekOZCYXChIYiEc1pKAzyHaPUYFE2ZtRZPIC0Rw
metyKjpncq2F3HR33N4psS0H+FSQH4zmDhPTQq5sy4TMKOYKFJSjj4PuV43gzy0u
15NENxMdrkgIuvYaWks/ovEXILpk3pNkmCbAhUF2Afd3LlmXCAAddgUX8q2b6SKV
wEUDKUcTdBwy3PT+GDpSHSYKDbFDY7LgjSI+0/Cd3RZEABS3Eh8n1cnNfCS5wcgX
WpD4/GOmYvijCY9y2pD/Ad+IM5eZ+CZFm/upx6wAHKZ0f3lbaT5rtv5k10WoXYsA
J1J2Jto5Qc1hj0rrXLnIJWQUFb5uSkXzFQEJfclamjRW+uRHa2tFj7joB2B8VbDx
OIaslkmOxCR7Sa4TXOuQ0cLab/ZRKtQt/Ve0iJEt8ZN0Rot1gcoRMcSEaB+VDrlV
VOj/leHZytyAMlzrcr0Pt3hCLrujLqxODSOzNmaA3EJNfF0Cl9Tj0mS5gAox9yX7
PZsbSE5m1I9qesmGBsTuemlxVBV5TdeuhlWRcaIywODySVgdYNWnAiVYV6hr1EwS
aoEnmrVgsay/3J69E+CeHDYamSlh2yIzfIZM19ybDJJBv9eZuTAw80vp8QXck/cX
/qMGAM0ujMLUYBEXojxgMrnZHN4AoBl5MINa26hS1ud8sfAIUEttmztESMwcPAVk
mUruifp++vNkwz7Nkn9gomEYzP4soHJT0xSrBaESVNzTNp3SIgtAhIkbV9NKb6l7
vBb6XMPlkxufDrYTmTjJ2l3WX0HaK3/0vBl5Y2T/Gj/0iotpb76hvNcVH50kAeJP
93BD9Tb0W/XH+O4h+OBad+L41fD1PtgmwX5yI1apXTYLJnfs8dHeRNNpaAaWcgC5
OIlfTjFrsfiLq2BxA1JmLqvbv5AzFFBR1NXkhXAgB145yD9SWotqCM0GhpZbOOPz
mB6nDA7nAOJgtBhL+SxpLB9Pcb8D0qB5ioexLi+9l3fRmgt5KIx+sntVZrrhS5lB
OZ0ibcGIGpansreqnl1gzXeSUNa6en9wEKyCO78BsyXd7YioDZDfj8U1hh2nWb1h
8tEGUvpdXaRAYhuBA/xuewCeLVJ0aHuNq4YeZZ5VXvzUyZrWsXh2wU6B/iQfwKrW
fWbUQ+Iqmaii87i/dT5ew3m1SNmPrEish875Pnnuefb6Ij2ErjWEZcSSsbS44eYj
dum+g287PUywpYnggRMmTKxyX9NCThJhgdXJI/G+0N3PIMjgFmVEopTQ1iQmTOA5
e5IO1TxeMVG7BJKgHYv500Mi3zueOApLqMs79DUQHq5dk9IaVnXuPmNKQ0NtMT6S
+HoslmzhgxppHy/BMabjqu5lYh5lkYANBWu2QpkAqCw7csYE3g8P/gIUqjX8klY1
TJVSual0v6lM/VmIh7jdYkxAoIBHCnOJRDZ6qxK+YOZq+pfFlQlcmozVEb75WU9X
TPL1Be+Ieb147f61KWIo7eTtH4XVodN7WEi6pd0KIRclSzG821YoU5HO9dOnxzXR
dycOBLDPl+23WKq5VGXiz/63YhFyu+bUPiNBXx6wS+KCuj/AjOzJPD+NY69mupZ/
KVSuuYGD35jMHTIkGmn6za4yW1OKKChqbmlSedR3PtYGEWXmc/xzjIP4cxXizrlf
UYHSssX504QcuipHSGiquDBvVUS3frNsc1iR+8fEc7iCfUAbqtbBcCBEmRXxcc5i
NExwHNCY+L+Nwpur3+GwxIdrUkWF3TZ4xwgqP58BlU0j7EtTqdz8J/cftEQKgu+L
WuTy0jgvNOHzq1y69N4oNqDBh1rXka5A8tz72Gid6Nmxchs18VnQiq8/Lkz8wJow
gJUE+bh1/ACJDpa78VTTLdLLx/opg3snGOHGOj6FAGq/HCcBN23kAHqCbDc64KTn
g+s/cVgl+4DoLMJuy33HDjpW/zIJM1tPCc9pPSvy12uC1KxbxpcH3HgB2NrQiKge
fmpynAlop8eQIvpFzo5IIJ16k9UrtG+fAoOfibUTCc+vuSxgnY8BHFrng0K3RhEg
u1DxhZph+gNISkKuHpa9buMiZT+h0LKWDuiL+0TABmYfYlM0fJ2tlURO7XKFLebz
lyjYm9kb8p8vBy6YURd5sQxQNDKrtkURu2exVY3VKhnnSfYKxMTfP/DJ5zeum86z
HbMh3acB78Z5MY+EQa4FR9Dd/AzkM49c7o9jzPMBpNUd4uDUDumT8FeT8BxpxZMG
Lg555DgHEgt5VxsXhB1UfZTZMimK15Y/uJxkDncp6OfZVd0IbZ9kl5ukAOMXFbPZ
lC9Q19yQi/goIYr7TqSG/tc/ef339XNjBZMy96c96/Gb0/QNaK6ZW468Kklw7h+r
+/JfYByWO7mU/JNgJVfILkeVEjU3DRZ44wbJcUV8YuitOMBHSJrcPojMpViAamrk
USBrbM1JV8tFLUDiLCI47vfPm67CXLQNmwfeCnU+M6f89DkUetKU69uBE29vaSwJ
xRMxrtR+gU0mKsm39w18RJXj8cHu4rLaeKwKokJb+zKZ0j13vWOMB/X/cE7KtNOS
gJ6+rqDeAWIrnkeUWysHYwznfHqKHj7iTC+cPXTTYXSjnvTOZLkMZiiK/+3tw9u1
t6iNcwcFiZjDM8+qHLVGcv2Kce9Gpo3Ox/ahP1xtPEmbfuvJnzcl642zAT+jIggx
WZR0L16o7MvuryVt9jJTjLIQEWkVoduoonWt5NZkBQHB3Xx2PZFZ9ysQgpyfksII
APW/p5nYFEIh7lxsQKbrSjeKUOesFKRf4O+PDWuqBfYBDKWQoLQ0NQk71zLQvVOn
Y56lE8GAvvMLi/0KznrUTs1Y5H1YAAD1ud41pj7CeXYA2tWcAixHwTDJHI5DRaPv
EavXCra1Ll1VEZRU8A+x2Vz9VGNndmCUsal4O7s50ELJQGHh65uWhjBrRYC/gMe3
IxosPw+vpI4YhWxuiOH0+SMyIPXQ+32TAcMepSMofSU/5FW2+2KVPDopd356jCvO
vF5rzZOuYwB8ia3//6IfLitHMLXyR0gE6bfdot7S4L4KW2nU813eBIgHz+vec5Ip
uE7sTAfJhEzbz5SpedIvn9s+T0ekUnaf9zkbDKXxtObnpIlD+r5F/G0HquUvc2xi
/WDWt2QIRSP1lzXQIj3/94rNeqrPS4Zq0glHyrMdQwhgonw32hwO1wwyhbHVYVL3
xGpj+PrPcUEvR453EYCajAFmwMvzOjV67a/6WSJd2fzMT8sD+jXnJLsNeWLcJWu2
yOSFDPC+oivmzaiH2C3iJy1PS3FcYjPM5EswNbsiylW47IKDQujFV0nNHpUlC2fV
t9dX/fdRSI7aua6j3ST8Qt+Qx4gr3E/ZG66dWuQg7LqX3zqysTJWU7sUBBHbeINr
GEEkNrTPzXxfhEtiFmk9n0BLSXDH3Q2O/2t+TV9NKrfh2lSJI4jxPY2A7QF1tW8Q
bTIIMvQlZ1LoCftIPa3JI5yKl31e9TZymIPIpoT6wyfeyBR3dzbJKzYHME/ye3TH
tqHukI4IAfIh7BR2yd7YNrcmTB8GsX6yklVPnuz7hpWi6foACZo3CHGszfJUP001
cjq+5lzX+0kh+BL/HtVF5FCMTLSshWAc8gZfxQfD4GwECibtTzRewy8vkyKffD2M
032QGYrscA8iNkAmpmOiz9tCS1NqtEGfQ0bMkaRm4yWPgVsVAFgKjaSP8VWb5vi7
iPz4aUfnZ0CvGf1YXWMR/s/fPD9a91x/9Onv1AnO0awcwwReEFKboGXIkuwQT9oG
y5piSwTNbvCYsGblg0C6D5e0N88mmOWlfIe0ixX+Z97wctu7kbiihl8GtaWHhQCV
SYC7x2CszFhG5WzKH6QDeK/4RI6e0IRCYUM11iYJ0ppSWUuY+KB1tHU4SmQv51eD
/Oh10S7BrpUdwvUAueKFewKwTp5HMmUt1hmhnoL8N8hh94gVYeUUv4xnnCdeP74J
o5LzbDSRbtaJZJzKwCeRTJuant6vwLeh+a+j9w6VuHCFjxnKBbR2sTKTLshzIWVS
lrBMJhxr/W1nAPSMtflwBzh9sZ5ofv+6o8mrQEWlC/hUy2u3d/YVBrD1XiMThYWy
842IZR+8GNopTRectAr06AWnnm/xQg8NicE/ZlOM0zIdkjiI7ErNCDPQApoxq4IT
dHzuAG4AE8gkBNXbQwogi5U/SUOg/Mh/uBMdXgVSBMP99Q2SX9I8krrxaEfx4rEU
74U6OZvy6B1L/WrNe6CesYmHVkYLZ3VMT3NmC5itsv1uTz4+cgfs1CiO8kJcKc60
pjMRW5ORNaZNMenSkgpjUM67xFtZuYHymvBGjqlCpdlIQXzlm2RDKPu31nXSV03l
bX0HcGkWs/Kgk2WrOHzVrTNFWCaRTjTS6+lZlXJDa19yYHrU5tQpAN9dhHWgL6Ar
qeFTasaRuwxpHkCTsame+fZCD+Tq5Az7nSiCNLLjnOrUDPFBXUcipI2lymGwK5/5
IyX59EdXEEU1U2Mkspt/I0Q3CIzI3+jbDXcNORSz/ktmL7dc/CCFBLFLRN91Sd/J
QGsXrUrcU9DN+c0QLdjLKRyez/j0IePFuuQ6esclHKhNmmpiXgftlNCn/tbHmizi
Sy5s71zEit5zSGmOEQN49/khEhUgzpFxeHwY3AeUFa7LwOzWzkO0wtI83E7r7RRr
u/EqUxC4elYBWrb3Oil+QU7qO1yia7TbX8PsxUhtg0tLOz5BlTB5hj0kp+DOOPYA
KdmIjrnhIWc0l2xkSAHeo5CWdZxrWMrkCyktGVOxhgZnAdFrfIi1+m87mjw2a+lU
SHXgUxrG4UtBHZ4xfcrUWiHKRk+fyY3APbes3TbimjUC7G+IFF2G/C59czv6JPcD
NbHVVF9tvcspJsAXZcbFU+izb5SUig5Y8tCIi13Qfo+wBHNYQwSBymHzOLnHMpeu
Gg4xmeXZwaGivxRqKwLBDFkhU3z3Vs+5wFcPS31QZwxeFxN75hQqOupv7zi2dgx6
aAsRPoinxQfAT5MGE9pZJV06EvlZKQPo7kjNdsiZ4LTz4F2FLIhwcgy21sYs7Nen
rZGAfHnyLz6wu7GowirneojZFF7Ul37TG5a5DKGb1D2riQGxNp3whfteag22VIrT
uofW73Bho25A9kFWV120Nwx874eDeuMkXVJkakYjdT6YcI7r7WjrThOV05YhhRdk
/i34AkDgzXCTMjDKGIZA5U5pm8XtVG2++S/lauM32yRpgwrHgvlFWu9ugOQWK/kU
ZtWcB21BqxaEgytw5FNyWwPcFmQgFzD3W4FU3Iy0y865oLsnTGn0oQd53I6R1RjE
r993rpsON8Gm49T68He8X0ZVGef4egj1n9T98YRpuwl3Bv3SU/C7KOZA513xyhS0
g8qoFgNb/NHplFo+HaExiB9sYAa3ZTIV2E7zOI+dzrQYIer8moa2P05ebk9CqtU6
OnSTFasW1VcApi3VFXX0O16q/OaGtr2dKrzYAGf+UxH88Zz7ETjeW+hpqAQfAihP
jL7fVBIxemQZ8anMNIW/pn71BtY3Bml/M+tPfgKmD7QvOT3a+WGva+BAN6DXkKDQ
KTK4AFi0t//tO/Qco8XhRdHyBk9TIWDLqC1meVusinrEqlalO3Nb8thQcHaeI4h/
t2KJF0I9FmcH6Gl5IZebjD/KppX4DgENZ4NmFyhF2sFgSbOszDMRp5/iCAcDgxSR
3NKffbXyJb3Ss1ktryDeB1AajCUGu3W9aEZ6MeieBfUfhp59ClWMIKmK0C54MUtW
+2iaiLOWJRq1pFwDFatR4OYVLJFMwNd9VJdZ5wN2iLU0qBZsiQsLL93xlB+cd8ao
50Rk7zRsvKUg0ueXYb4Ybh2r03+fXp45HDflyIMGeiKGkVjYqNul2m1cO8cryF52
bdjuOBu/BCtIdqP5ARn+eWRw8pkjf82Pnc12bI4HTXsOyd1hQjriJcHpWzl4HMXx
2/6mUETfS+q2SBfJcBIlGhkQIFi46S5jKmw3o/LCRRGkFdbqh5qEhXGR+F9gMxCE
yh8Zl1UICmLa4GvS4V1lhKgDvFXNkjk8Gw/lLsYo5gev3xxjfA8aFH2UkPzsEGg/
93PLTlAsINWzhBCQl+9n2oI/mRnXJVIlKdxFSqp+TENHH+dKhpyvL0GVNb+I1d29
uL1qZ87e32zPCm42Uqij6YlapccZ3o0/AImid53qRgm2zeH0w6FXqcbOU0h9Sce4
I9KllNtQX25aV7YOSbGT9sjvBMMvvCab1hWz0XfnPFmQYuJdLS7o7pBj3vZA5YuQ
0pcQrJjfLsOIVu0ezmhArQG52vrzEAF31zx5UyivRljH4FhnsNDD6p1pKL1+G/SF
AkO6lOU1Y+hcMUcH5u5o7H9rcVgpHM3PVdpIoOfavd8tWSS22pWkOIBXrEXwyHIr
0HBzfiCilW/Dqgpfayss4XozO9GpUuzFgBx1mtiOlWyVFGa2V3xc6y+dwILKnGs7
dHjHo0IJdABXZS1NqesAK3NsXrg+n9u8usfx0QR1LGzAeYwu4JQ5BubyxNOxO9tu
10L4EWvnFnOcRjuE/aszgzJkUc5kAgn7KxIX/smyvv1OfpQUxTGw7G9bpvUUggIB
CyTsSKW2rzVjLthjeFXggCdXMWeDwPevX+GLTLmMyv/meGelEaXveXf14EKjkmqH
s2nGCs1X0dUewpRYvvx5y+yZUOJ5nhPkQNzDh52TS/n5CVoWSdR92wSGbI2HeDpO
aKB7j4yxGwVbya2wFPrF1fycU03ynJntzoN2Lw21WKLCVDhYRMG4A6xRjOwLi0GO
6u5g2uLQLToABOBTO4gt2HnMUVb5d0xK0+6aDarPv9RuFGiApg3Es9prsACVK8ea
q0N2Q/BN2IcJv8xxED7PG9S/cGxizOBePb4XZBLVb7JP3TL3oQNVfOqbQi5cAFEy
t5cnwAGb4atwhO924ypo0Z4xvcItliGVizrIat0yLUGwDlvd/oir2KMhWaY8YUEe
TuwdgHJ1VdlF1agT1nJbXBscRK+CB+BXKkRzSeFWy2cNu9z8L8gfuv3gP0QFjIxk
pnA9FbwDsRnQX9ArUFMkZvuCAqOxJI+EW521ltKY+5SzRatAa6aPw9uRMKtk0x6n
02QQDvUf48WLF67hsxjS4OG0tXDMHRIlLQkTWbZDQ5EksnM4Vq8l4km19A/HHM+d
HVJm0SHWAMh3BeGtbtDV/gttk1+BUQhzQiTy3Xr227O4NXzEPv5l5aiKahc1fCSc
OFh7KwPY1S/J+dUdp6vGswj3I7bZ5Fn2E7K6Kl78+E4OXSrEhFxFFXLkYPgjmTZo
avvA1qzAg9UJafd1T737WRfCfoQKt6Z7hUSCX9dHSdoHEw4VVMuFTBwZQbNLy6rW
8mSZcTPrWTZijfK5UtN+TTw2nhfqpFglpU6031ZurctyAJPG9QzorNhXK6ZUrCYb
WdUIY/QwF84qc53ju0x1seiIsbUL3MxKnO5dT8KXZ7omH/NfjFnEiK0R8mDM3rc6
lXJ0b1z9Z4yuuQq6tUVJBzvf1k0y7cPWOYWNi6B5gjpEddt0U+y9e/cf++bkpaNC
sv2U9dSg7JUcroNBl3vhdJSOFdkRt/iy4V+LSt2WVMbR6iG6wNoywaIvC7AuIXOu
8v6WYqCkvH198Kymyl/R9rQGYC/SFSkef6GsZ8CdQo96kiaMOrmAbacXmvcera7k
D1F+0eW3p5wSWMQQR/AdYIHJKWHJIvgRAsFVMbJt7LgSB9NuprHHUsw3nMrcqktW
SE/O9Na3TghzOZs3JazvnRWPZ387ZC83PkAj1rDcah9bPUv8dir9EdNC5sN7TVXI
7QQAL3RVzpqEWJ48KDmbf3gqKqdo7hpP4kTmklM0HeRx7gAnCVOlWnba1XAHHmww
AKqRuARnARRAmyTBXWzTZrx06wpuqsePp7nyk0OKOvRoGXzWKCtqVnCqyX9C2Ifg
5LQMvmge1SDsRhZV1/+OEtra/kZ2jXLMVVKtYsqZh2WGapQF2EDddqeKgBNbS0eM
M3XjidAwS9i3HuVMb+krHV+6BDnSpRQTFdIarJT+mnHj0b4YxEhL1T++2yM6XE3W
hTy4ZmnunJa8WclYf48II4G+1hTnfTJ9n5+kT8JiTj8ngKLPQqawF3fxVGLiI0zz
JFR+RTwqMg/tkKC7PKS+2q1TUyYUbZmzYuFTpWIkxqH3Xod2aWfxcoODm7cKrQLR
Vhb3HHG6kYUjq5XTNqL4PdPelLqzKQNU4TLowuZyT+uSKVYPBEIuN1TrV3GFDnfQ
eSqpy0eKOuOPUESdygVXaPG72DWhRIWFUaWRFUbz/IK2kIYauuubUKrQKJwSq6Tc
LuPezx4P4Z/+lff1e6UhF/VXE35pzgybcZ+rZLfvvpiJ884fS1D5f1BdB4x/HIbp
m0f5DVL53EEC2s6XbHL9Ep2tziHCqJICNxbeULS+QJAYVxJGkImvR/7xHgwvXFjs
Yj0F9/VjEp/JbKFTxKMnp3m3HonNsoytJ3AEJ003AVRyYnso0uwByT6Sqst7oQsr
dzAWjIebeYj5Ar7svA3mth9JGulzdnZvtZl2cwtiHRJ4a9ao78/rBQUmg85MSXxo
aFsfa+ulKpSG/GXeQAa+l0DUD5NZ85Rr2WMP9Y6V8LXyTQ6SYvl+e8TNkA9Wjobd
cpLBqRvmeeKARO2YQTzBnvbVvLZgEIAQUC/l0PVm46okP5Cqgh9D00k9oxcJksYs
4AsaJIBlrdTjJKMEdnAZskUYtjRzJFuyJ6Ev20NbZRaGXx205CRvgT4ftwP4UhNC
Pt6n39NXCqDIxPkmuVa1NH5yDLRtGv7MFL2HO5bVMy0Nz21XTZZC1cvEEmt/aeEV
ohNs8B1tityzPxlo1kEUCeyfY+ibEIqFMV8oIJmFUHqWefnOSbxbLCPmwQ2Q4Nv1
gegIAm4o1T5Z2ElA88fT2QNGrSqoaoQOD+DkoqLHyRg8a1vJKhWZZ/X/6RN7zUef
JS9hMK1hOKvj7LIEUp0RjtnIk3LWOJOO2e/CM+NI9FZ8TDMBcxEIIG3WTFhMdiGb
KzC1QvuatWRbSZYgpZSi6dY9XaRz6N5JUYVM4eHYu5WamjL2l8q3bNNXcPG8Q6nQ
+uqLiwlMA0pEyXwLQYUpSXwdNonXoQ/gzUtBryK4DnhmWb5QyxxLHFEsa/dEAFTX
9k/fw1yvOr4UQmUnh6J8aoqX1u3M+F7/Uh3z4ooJIH20I5B7KBJkEUk7dWws7vMq
PDmlPL/SzmW2+jPW+tmACsjkpPDH4z6amiim0B5l+M/d7k7Eo9QtdwPeGeagkPIE
BSYmeO+CKwv/O87bzAX41Utk2u7jTtF7q/Y0flRy6ReDSHX80cUFOKV2p6P2C4Dy
jgraQTvFjAIf1NrXutQkFOf/C2AZ2QIIkgczKa2t3cJOx7+rKtjk//7Y0p06gwUO
QlspzBggexXOMZ0AvbybOHu1rSt33Ndg9V9nzyYxcGCgwajBXYMQLdJr3w+V4Zda
/H4jWXKIlrnJIFg0KkKQB/VMt1CgokiV6ExLIKxrsQbpFcDjsd4Pl4A1s9gzRlBB
lOtnMEddBQgJkMF5TfCkAtJz+EIGB7OS71NUmrg1gfRLNRZmztFl4XjYupVq+0Ag
odfThgfaQ6j825w6kzo4gpodsTNy7S0T/xb4Hg7ubAPjKyKEzpqxXerzOGXc+fGT
MrXc4JnwC/VBMInjU8DDPkV6XpRnSIMnjm4lxZj3FTV0i8n7Ijn/TeOl74ss83pl
n9KMz1bfNH/9h/9QkSxxyk8VY55/Y4RqlGk84ZgOZs/SPaHjZkOMR7QRyV8YNSCY
V8U5Q1YvvZaJVuRNTJ0K4T2nwQbq/64DZdX2LqcpGDjVKfbRRzjAnAGTS2g55O8K
oqUu70y6ttNWNjdsCuNS3zwMGyCXi0yM/HpEqKDBsMN4IK87wgtSA9FjqFMngRRX
NchVmkt9lTFk1vHqIMUtCTtqAHk+usq2rnJGS9B4YURcGu8BPTDYPUEw0KWHFi2I
Qm7yopdbrVVHHjW50+3mcudSbZ+60OUUu96JZzDBkf2X+KUsC3Bb6ikxSuwWSZMG
w4FpX70qxHhVPxiwq5YVbomU7M9QKmy5e4i/GpfPAMGskMty24/4BpCho9F3Mg5t
ONdacczKRvah5TlSw+EdW2eeAwa1i1hEsD22ibK6WMbUmgb34QQbL69+i6iup3Zs
nmZsIOrrSRc+VddiK56Ib0HBLBKS9qZ7zrtnWignKXBbs9DVfqckf7m6qofM8ruI
+LkfAQc/bgcWNUe4x8RPq3EuqesJYGxiAANnP5eHqRvKgvBl7pMJSDDd0UqNH1/U
tlo5hqoP9C7PG25W1WfMgtA2hiKbUtVcPCkrttStRX8QEqZPT+C4c0/k8Qakh/eC
gFNlq0IXg2WNxTg2bAuogWda8WN5HkMNRdp4Z7Y+0B4kLeBZktmksdzfjVlrcRIQ
G24GWby68egHC8+NQBb+6nKEo8km4nYzof9dbY398oFoOkbhsebSc4deqSTVHDBs
yFGsiydE6+TpbdKmjHlxCQQTXONKvU8Z9i8itwoC4P9+snz+8DHI50/X+S8ZDmop
aZB9KTnPoVZF8FCHZSJnF1wn+h9g+dTT9MFLjo2Wy390MTNwtN3BPbE4faEI6vRC
L2IOLnIWVGoMbZMWXF5PHc343qZgF3xRjZp9oVN8xAmE0Q+Hjt6/MAFQkX5a4vvs
Qp2WHKmf4BM1cdAgGlzFHTVgbK48ibkd8AF2PWwdltKUhzKhIpYNJKQv03UjAH7b
MpYsdzukkl9iYc0nSNe7JQsmIaZkbxjXwLs+GghtQqaWcDsc9ifNGiQZIjoWBoLy
1nhYM7PUN7nbAl80iyuA8HHxxFHFiq1dbPNvjZrHHbf3FS6YFQbkCJGVijvkP/rB
Q/lVQl35QFp0jCY2UmsMB820x7wsNKQFd/0OX3Hf9iwfVFSR1ZfbC7y3qJLAUmVd
8Xo5+N9bRDynQuEf0iFz+54QLzCAKZ6Sfmd+iWS85UfSLMnIESqKVQMSccDSIwoY
IvP4nUmVCzifcA7MiGo9th83+gn/6ENe+HUsx2vdq7naTMpJusd50AdKt/+fshYy
Ff4IlFKfm05sQik7BpowaQIltyiC/iF+gYdtiJCNyJeVhr4vN3lB7kw5AzaWdHr0
RjRsXzMgHSB0DhrT8GR5GWhgSlqdZnAkz5an6Rv+RMP6DmIyH15OVXygdl12oIcU
xhbphH9wmu15o0MNIqONdl99kJmE8IbMrfbiSVGXLd8/+Vv2pnwo8Kug7tf7hcyx
xraqDx4GBbQcwAplGpKY/Z3ZbxFR3lSV3G5c6YajkS5ht8CojQ84jTHxRl0tLFws
Hy2nZUy5HZmQbdtdc6t+NZzYu2ZHxtp282FPf8TXFVtB0ocxja/rnsvc1+G1+RNC
f74qRAcZOgH7pftgpX1aKdqv7+ePxcZdfcGqGVu2v6LgoFQclbxpZyAinMj4FXAR
fVSzy1n8dOBVeOw9Is3npHmprWw93jzihAcWeoE14R+/vYSQIFcPrMh4sVZIw21O
0TasH073U+SNQ5hbe5TffSQyjuuwZv2fqO6HlS38CsjP9EMOufIToWTjIDbty8/2
hDlKXlDkC7CyEcwd70IVaJX8qHwfiXIXdzcEbJ+5Uxn4E4uxOX7NuYa0fREoKPIQ
ouGHYr3/yf8d0zsxwLGYo7Lk3uhOhOhL5JipZ7Q9DbAgyHlG4SvRMyoLJJUu+LD6
W6Qo6GH9I45DddhHJMGebtmlyVUuUX/0oMPFghDq/6v2tqm+Em/vJg1ujI1u9BOK
CtaRFZZ/Hb8Foa6Ojrm+zcWHWCl5B+hlKT0STplLMuyEb6tyw6ASsCPWjNhVr35n
9XiYNNHsZy3EozR0BKzTTOtNMIyOVNtVEms5qluCHz/MTlOSvM+PC6zpNNKZCFGS
hUF4XF+f8K4fhQDHEuxNdd5Rn2H6GVZeIoxlA+EwPh0EmVpO5cRUBn7QnRZBLWWB
oWKYPyj1CJ5o4cUXNhgLm+cc0SgElhpUIm/ieqzdTCsjpWYbsJzufrf/2Y4t4LL7
qfnvKxUcXGkmTMWcrXft3j3nvFpuneIlMNMWd30JSUfPEbpcbTwsyiqYlgVdf0Bp
+Y+PiTgncMPPqy6YygHs8bHLAKs1MUTAQAWId/Zc9B+TmZmzR2wi0POCxSht2k6R
K8KzzMCdoOMaBSvWUOIqQAIIWtLcaNEpYuhdCQldfey351RKJFOVz9V8fpkcE7Mh
hhIqyv10DYUXgYo89H58IQzQ7kC9WZSojsoZtXVaTI9NCRk9tJhKM1Vt5TgUratX
ZakxfpYYp7XsyAVxWx0w/QFv9GU3fPc+h2Gh3GWHkrlbgc4PbEjyalYRhwv1XgNu
ei3H8IV1Mgp2p6C6AbEVVlqvh3X8TluvI0Ui1TxNymxH3htERHCJr9oDRHSEwxXF
xSqagvJ6z6UvcCG3bmLVVLMuY15v1yPMfhdkfzKxCsUbI44yLNwMRkYEKd1P3ONz
89qKi1Rd4jGSTRtZn6IJD+HqQZOQpyQ9baJLHFXB4g0qv32qjjjayt4j3tXlPxiT
bshyK2/Maa01MmEyscYqy98T5gMD+EFZ9b9b/uAMXMdzkWCQkmCiumw+r8inNMbZ
aVzJZTmAVRbgC+sR/9dtfUTiBSpSaEca1oxzMsZhJl9AKJ6CX2nfKc4Al7WX2KSW
mOzdD8HkgJkwix08e54krV/AVelOuOyvBO6cLomUpo1LwOpsQEroy/SKX65dmOry
dJ8EtUtGOMk5TugmiAF6ZERY5ES185xkzN3odCeKRANHuQ9UJR9OD36v4kDTaPi0
oYtIskiHmpSA0rdpPnJ5hiUfizSL+fkId4LCxdGIzq3dsv6djkKXJRwaS1YD1en8
LVIpgNmMUOjrRSWoZrVSI4HHKMATDgg8BDqWTMzX/XIeiXPFF0uR3Tigfgpt2JX2
46a9WjEANo2tEqmZJvg1z3fE93BnPdZSm+tNKGMq2MAldl09HbSOJNDaKpHwa1rF
hI6wbQ15mFFWZAXfn/EgPZ9dye9dHvXdyh87Qz/BcHDebKhdBBpmcZtt+O3Lh8RF
/saSylKrufFTzBooQZMoRiS5MwykHfvxWUaDvZWWv256DxQrJuLTLJJ8n6ARZgd6
q2tU1J6envFkJRVyHDqA1foHhVWTNO0Nq27cYj7J++BNtfDqM+46LMQsYPx7lIGx
b0EjCdrm2TI2bTsu7DqjBOwTIWd5cqt1WcJJEWhZIAXE/xYlw/0zaw26mI1kpxBZ
Bn7F1UFwLSYuQFMinxEmGFDhfOnhRwtjgefl6njZosnu0VpM4b51uGpnrk/5HBHV
er1QLk2NTlVOc1yanPPbHe91iW35ThT4NEj9C4XX/4wmvsQ7KYe+QAx10tCgcBfc
uakMxzvfxW4+8jEU6VE5s/JZrQCUE41XGuZyorLLxX32tETEjG7dvUPlnHSWU6R9
98Ot1xQlSlX82HoqyfxtgBHp+6NOVPt7FzO379MnW3Dx0JO/Hzwe60IxazCKtIuo
tgomwJxvsKiae+Lvavt+6asVBv0ixTboWLNB9eEIU3aq9WwoMO550VhIHRc9GiFh
3ZBLHZ8k0BXqifFX48SPyIZwe3rcbX8LvJwMPOZhor5ibDHdo9elm7fxrr9JgrM7
OVfvX1nxYGJ26hg4O31lvbunfyQY1RrUlWxu5/ECaRzD756ZY7ItxeKKW67PRkbg
PklIXQl/JlQb7yuInBtEnSbOJzkwTACw0KJPEwQJfazGkXl3guGkc3iCHBf4OR3C
kzPNmfrhBAHtNHB0XHehFT5MsLRV7qaASew5dwpMjQMcXFSWrk8R6wt4d2tewxRk
hU7sEjlsf/ruzEfg92vpgBBi56uEMikwicMZpcbmFpio11nfJwHkV1qn91Kqtfry
psiTHe9oj8Y+OizhRzD1eGibpVKx2r63xjQ4krs88qcB6EwiNb6frj6jyrMAb+jx
go1Df4+GM0EgjEbefDPXTh0Lu6tuz4XAaOYIhh6jMMABxtVq3VbsslAF8OwLSpNY
iJe2SmfzQ2x0tjZ47bsRorCuTxY4BBQzES7s2k3sh36RGLWDEg41RKiXGU8f9bag
HcW5ZbpGZ+x/tLIJcWWsljFMMwP7oS9rlQDp7l51cQYRxaLf/5c8+c6KHEErCO0e
aKL85MkKjevRfMrfYrGPbUtcQjWrQidR2EtlWueAQvKFxjQZjPTPEz6CpwQ9p9zo
FGTDBF3ZiAVja1pE56BvOKQfTVwDKy7Zd/cC5deJoFZ5kkZqCS9xNZsDlmC2ZE2D
YpJnSIYGAavVDNMAVqm0w0F0/vJwXs6d+gpfJfXe2QCutuJb0VWL1ginW9EHbl2e
ndBIOhsEKhg4kcAafjEbj+B20ZOphcdroBLj3r0X5PgNnn2cf5Z5hIJYGTSO0+E+
Ky51coev1VmK4P5ERoRJT7cwxFbtcu4QGtn2nWYb9Dx10Jsk0W0N6TKsy9HpmiVd
mqv15LA3sHS85QvUwNsrZ4HtDitGYoLOmpKAqo6Vg1FmLJHMhzT05m0pIrZeY3vf
8py9yPkDiif2HS8d+vmFAkTTRLTRr22nzkrJN0HUtPEVMhH0ApcJXsmpXLvnl66D
/2AqSlXx100bLNANNXX2907vQp7Vke/eJVs9G6ACyusBdo4EzDrw6AeDCA0OruTO
h05ZE/by8+0Z3MtvPeOISk4J/IbKC10FGugP95CbMjXXGHfuxnKcRXksgiHpVml0
AZ9zpLM4zUYAgPO9uEr95kiSPZg8U+FPnZBN78hAFAsxurvPMsx4wdBgiZkb6Q0S
V+FSgmrRTzxF5kjOof0HCN8hyoo1Gs1zYukJ3XENFLfjCilzRGdJHCAFO6pRV2Fy
LJktkqkZhe1hYCVRvA8B24ztWdrqH+oPTX+bCCzf6BtkpLfgJyh/+Cvp7BPKGNVy
owAW9AMbhr70zzq7Xp970oMb7IxKGr8gkxSuTJzTnkdnzW73LJix+EITRo7ke9Y1
I7mimBmpcZdTQb06tl+Ao/TwmjcpDO1cShAQJkSk+eme7xd5+NJM4L5r5Q0kOE4N
wJsT5AMKsH+XfVp2CnUxdKtwPvOSRaAbp1iC0MRMER01WHhV3NaUGnStij3FKbVe
/C4ZfwbYAyF1up5qYmul5aQA5G2/8/Y7sQXl5xZBAZbGZINzCz9HVmqM14g5DK5M
ja9JqF8nwu3NQ2vHt3DOIXFuPQMzmKYpRF6ihXBuDU52QVm7bnrSzuwhAVVuoG87
9rtGyEwnoHpjieYkcHNGFaU+9u7mIxN8ftzZlPkomPFrg3ffPk7+bXpygNq4sTF4
eZyaVYxaqF0k8yyBVAUNW4keLGT7Ky9TTkQZEztuHTiLWfhb1WSakPeyS2ajU0vS
S+JlxzVV7HFYNaWYdF1dBeQudhr0SNEsgmTxZkcmVONItATrzRquMe9QnT5x7B8e
XI7aQ1bMKOGKQNZv4wVniE1Uqk6zZNOyX94w/rPmSlGozhZyKyRGKIhSsUKsbs+k
EuXMffhYQjn3YjGIwMpnYpQeWYRKuMKUj0cB1VMOkT3VmBP9q4XkkMlDl3lsQO0g
eThwntcWw0eRZvPzC2aLL/oq3vliSnlDycKN+Yz78EkB5L/eQTxgpBTUcTOIrhXB
/jb/blHsjhtUIW6hxKO8Xww2ftO5bf4wzlyzsBpp/HpMRRia99Sg98jKudFPPo9B
blrMX9CW8WW/MgE0fph6PRU3pg1g2cCisNC/SPE/SvvD1fqyCzHT0qXcf5RAxn93
PbTgBXlV3nG0XDgwCAGncYjE5gTfeGl+hjc5AN3/BFm8CoAaw3QDRHmY8MedQsLZ
RSwo2vTmEiPdpHwp5ZHa7WJFNA7rVagzAQsTIg7+EXmIWs1rBtYeEt5T1xnJYrkM
7N74b1gnzlGUxwqpuHIfaEeljTHvzfaW+L2HCbu2aPc6+1fFiHnCMBMrDgStOqhd
VEZfMCa0mdge9hAui3AnSR5vJbNk01LqpkMY2XoxRmlZ1I210cdInT4rOj+N3W0+
vg6Z9MddRfCmmz4PTVV3xKR6GHpBTVjpGlnxS8VmGJu1yIsOgXPi5qiYGHRtf9n8
DyBNvd6kcizQl2Aay9zeoCY52JfbEOCh3LHwI9J+sHTR6lG7bK34yb0c4gHDVzXC
b4IXZdGKG0UwckFnvB4zenzSeKw5u4wGdaQGXpVjGCKL78igJ4XxmjE/z/Z8YMGJ
VoKIKXNd0y22qnGrbeV+z4niknlBVMLFWEGA4r/Pvm1o3ynhm0fw3GQFjG5Wuf0e
W1sppMHve2Lax1nZzkmEP/7IFffFUA8eTtFOkxQ8yAeVmEnE7rSPZSlSzEmFNiCb
4weeG7x7EehftVxzHiAlRfeFh3BAOFMecLbFo2hQzxY6mHIklcXTopTT1fvUR7bi
QboxdO60H6fbNk1dGeZ9eYlWHjE7L/nnm7zcPBlYouOOTF7RX8TJXjgdIARVDnIh
BedvjL0uILhEvRpuqm7KKbWEMk5eJSvrFP8m+Vs2EfYm8oF/TeW0WjBqSNblsYPq
pdFdiTdA3uUQ1pnWs6ZizjuZT7eGuiy6/b+wWshQ3NIlykedPczxA7jMhGw8kSD8
eBR1oi/aP4iFaij6q+lbkbsQUbK3cnMt07qA2mcZicUfpE2xb549eVrVb/E+LvjF
+17xhaEDnQBi0PJ3mfd1t2nQSnk+xToxdTP1VESVJg4HNhgGQhpBGBmP0qL8gYhb
pgsghb+7kmYL671RSaFCTkSOAIa5i0+nRGu5LEWtlfAa4jWlyF0eEFXuBxDaFHRU
oLhf6kO+Wk9p4TBBKLAo7vHJx32yf1juJrJEyZUpdUZA+cdTRVH9OQrUFkbiYdYG
Oapoq5olktwfiEBq472CiztmBbP9cHejn2FEnAl+H2keKwb8gmwgLbzlaqyYN8jD
InTfTXumJulU9yo7aEEQXSbA0PWBIzLt6LZ9heXaVaOVIPXneE1S7MXA3AlBoxJr
vvfDniDgxKmDnxAPlsP0PMYIFSS748KQWM3hHVFKvF0uKmyGtfc1W4teWcrWFlUg
EhPNTsH5wsNzFG4w+tSEx+mdobhWkL9dhnhMr4uwzlsEWNfFWkXCAiP9l+1IjXYS
tSS4baqsCZL6rc7hwiOhN69zK9UQwyIrZMGGSseSlIJ0K28RI6nSHVQujyULUy/f
ZOWCn/CV4fYF8yuwmbgbLXPilotaYgcE4PMDbqQoVFg6SzkaiLY3Kk4mjN6FA2Kw
ZfV2+JW4OKBFLqpNpmhfKpip0f/VxILn42K5QGCGvUuc/2lLK2aYbTI6XQNAGpWr
K5Beuh82BNe2W9JB+mWVhGuPc2NtiCV33yVhTZ4jgwRAzO4HBaLdCRmOOrP8ew0e
hF0lrfeMHp3FKLB3Z+tuuIEyD1QdHm038jiTuxZanazVR3ssGxbNaDTKcvkzh6VJ
sEP25ou0sK6iOjgJIEJ2+2MqqyMEbasvVPxzlvS0OgGig3r1/IbcKOSTa2IhOJXA
3XO+jbF87NcEYZtuJKOBq45sqNMGzerRZ/pzxEZ0zrfcSUfEu1ZU1MXOipnoESYo
ZZ00xRcBj+tr4/0Xxs3/pz4lv1y7M56tCZQfuYhLQIRRZSOY1LNMlPwsfNZw1pbc
dA+TYEQO5FQZ29KxgXKOxEGrKJqQFThZc8wleKh1K4SGOSS5AnrdcN2jzQ/RMAsM
WvNY3/TzygOJkGdDJ4W4J8MejtvxiTC+9rssgdgg/EAGYyvBIh5kXxdfvCpM+V+Q
TtjaSg/Z7dhLOtMRnXaslYRmddDdul0MsMORFt9Xsoj8b4PyA0KQgGOIchITK08X
eGwzSQzhbJ6AzAUNGlO3N3aTUEC/LBFntQXAWpvCgEHEGMjRiC+CuZjCfT43IovQ
UgqrYC24kxQ9SpGtt6I7WqD2Y5M4pFt5MWfUzB0buKQfsJ6OypE9rb/+KDJU+kTy
pBu6Eji0p2YgZuVXIv2nlx3eCB8Oz+L9Ay9uZ2H44saOxEg8O6GEtmRlDkc9hSx5
w0ow07AQCQfbYgUxVPeobX6lcYYBu1veMXsLeCGtJwKRPPJAXgcXbNVhOI2ew2dQ
U3rOXwDweL46/x8jBgm9pDAmeTtC3cNhwBSUcJRDHk592X1hNyrwvr8bCxS0KLKP
6uC89VUAEZ6Ro18vUgiKAvupfiIQBO3wsxFZqB6l6M1zE4LP20G/IXKlR8kqVzIZ
bNYJE+iUibflCwpE9UlU0GbFvcAhyjDk35v2LlNBomDmhj6Q2jA4KRqiP6P9Yiyh
u695UsS4jQgIX7oHRLoaLJlh8FGy0b49ahNbqGuQjXjR1XfdqAP/rF9eqihlHxR7
fQsLMPDYYSZx2duX9MCpgd9P8YEpmB5L8ZheibqnArbdsw4Pt7Zjxo5xcE1R7rFJ
RDi2cjiO+u9Bre0e/IheoXuyptZEpM3M47zsVitQ2cZaVlFXwwCyusgErlXxu6Gr
EPXCCFqQeYehJ19Aj0hh6B07xB9BDd+2jWcMDetKNgFjWSWjtcKkpH2DT9bI3U/Z
JIDkXAcmWoVvmHr7TbB8JvNWgPNIn92Vb/YO60vA3vIip62DfSXHZtHb8+RwhErG
tkGlgMJ+ebqQjPm0tsakLPR9KbynuaDTPJgqpN771n/zy+2JggK2RBStGBHTS7Cd
zHGy7HSKO04kP4n0sT4N1cs61FYPi2CEtza2W3EAW86R0UyU3vbLlGUtkYl+Ajvr
pP7hJ19oM9K4lLVdttHRIVvPrKk2NxwaOqSmWynmJhtvlKbhlin/BJkXPNfk1m81
91xhTaiIXXWy4J8y6QekLsT+8sJsA/PbyxnL6ESRE9khJz2ciNP75g88Wj2okOQg
wmMj9OrnAhj+TuINc3B7aWJmJc0d2nrV7QnG+fzaQJUE54iRw1PF/P7c+p8r9k5i
F4202K7twUnaBHF9R1y9NE4wkGRP4e2tWpchcOYQtiTNzqcLpZ3OnObrFamiKEgs
glqxgqAfVS6I2n7IApOJ/2ss4XM5xxpVz2ua4Q9/nfUqFUlRku5n88+cxlKahQ5Y
82YB0waq7zDPFV7J7rNNoUT1HtZ48BRo/LoD09Y2apJF4Rbj9eZk2pzfhytR4+CX
7KNoTt9ivlI/TjdAWfKEuTKixXREa5uvgK5IkFgL1obb5zRdz5fCy2bV+N0mH0So
1flzpcaDnNgr+tJYTSjoas4EJDkyVPOZN0bjRYR9LH1iNmACAw+5SmjbknREj8hK
VV1CszIxs/rLKWkdff9oM45q5GqP177elZeFX5iRTkWjTjjdCaqXTprFnmoFv4aN
4yEreq7hKd4L2+wDZMVgJeb/ecoFNxlyyH2EXpNHLyaPOSCGtanrB3wVxx3IcUA2
VtWNCq4iezB76JaBm1Rd5bL8MvpwVjAJepGvJg3navaZLd8YHVac6ipoZ5f7MfIF
Rlmet3JpKAohNExB8MJKH8PxGQ0jI7hcSl608aGFfdXoXHrqlJgLGt/LoVvfJKG3
0A6MQciOpUTq/UE1erCxQdND50cIFzv879xe2RocvhvgfoQ5U5IJ/ce++eemKyb6
x4UTu9JYtCgLi7eDx8Gh94/vktYDT/LGVoDUt+7PLm3GhGTSnzZE0Snc28oAC94s
FAEghxYTV3Zi/rSysXBPxihRQrbwtaEh9sNotVtgtmJb9Qb0XYXAoDCSrlQlTjq9
80xjY1c50fjii7NRw4VzUUwGuGhCVUfSHmg2weNGVE9BUI4uh3LTBq686UwFlx+Y
WYnsnq7+e5NjrPlk1tYH+t4f0ifPlmMcYPZFO4EXpdtaboPrfo8iYawPb1ivF4kQ
i2fa5/HMavq3LMBmAuwmVzytEz1ZV+DXMhtmN4vuFUxgiF8m9uRo3PHIB2Tt2Ywk
KKC9zLzejq2MP4xQL9hSp2jy9WjmVU9b0y6uZeId/Kbu7kxWqZz1rwFbDYqZVZSu
ECYLv7sXsB6zoROgUqfqr43p53o6BRXfWPm+qh/2d3segivatX9T91aONw05sLNC
pq5lcskbKEQx06F3X/bz4gY1FyJ/hpU8vHflefDr7t1oRvGuMZUDa/FNC5lNLOSg
8xRGmSzOHcfBeASEz4iuOsnQvMUDCi4mgLpuVNW9oUx6h9g/ABcO8+YrQEsIhCYl
D+erzJH44T1K3U0FMVLBx8hqP9VN+DA2n43QWM+qo50pwBDkhc6U7/muqo2dzZlG
owyP4kDcmnOKxQAI+6gw5ekWpk3zfF1wrhVe21zz+yqy+NNao+Vh8uio6Lldd6n8
eCfKTFVheluAzFatT2THiF+kNs7f5sdsqSGwHdTEkzGDs0PgzFZGupTtKAux5HnK
IfbMCDjzIKivS25Xr10mWERDVZC3lAm1JHNmo3cdNwVlxhyUHQ/A/Iui/tX0KpNF
NjqRySpsayIxeZeoqFUvKGp8YTgnzP2BRPnwEGYSiz0BMBpWQ18mEwJOkZrDJPv4
6upYlrohaI1wVh0+6d+JBO3wEIAUM8cb8oOjBxH7IeNrCA9BJ7K6vzKbKpx0S6t2
wKrNfJyQFTH+I3WjtPO+hFR/aLDNyyzTDPLIsTmPJwjLcIiTdR4jRAH7hq3OVGkJ
qBRafIhp7QoA36ANkO6F6szrVgREJ6kpOO7P8g35tbG7vmk7K8ivxR1+xm8IKAr/
hU/24/7ItPvqe1vXUbrSaHOubpHlDGyu9OQ87AIq7k+Vn9p8UsNTQP3C+ac2aLEK
kbR72q1+NBLkwe12C6QJLQlnxHJqYUhAeeBE4HSx0KyrGv42dVgsyAhW26BDp7wC
zzkwajcecVwG3LkIDx+ZqjpK5vaq/M09Gg42h6TQVmfhA4wrPvfdl1Tu3WjFdJDl
4LG4uRaDQrySIS+Ka3Ngtakcn6NUijBgcFLiC/Ib8K3bMfx9NEtA8/4r6YSgSnMt
yhXGOUyC4MCmXfdjxo2q1Hm+fi8EbaTxgM6xOB/AmbatqZqruBeUYa9/qQ4XwwqZ
kxA/vjFNDAqHcyZj5BCPSIZYiyjhbxipsuhfx5kHFKVFPoM52OxtsAES/bFQ38n1
uWCnwniUnMUTxp9V84DZt932NA7Qmx3R4Tnjk3Szo2VaXiXnBvD1Ll7mAEH1NvO1
W/Puk0xbbnbAiL9hSGJHyhd0AJpNo9WXoPWCVjIs5uUBXIjJQeTagzV6DNMaxlGk
rMi9PlqqQUOIHIbrafXWCpaiPjIyIDupmkxVtsZ8tgiUKolIqj+kk4sClpXJ2neE
NmF05ilxemRy6Q29e/Rgao/1NkTZ2KDYxbENJfvomejJiWRfvuCvZS+hhdyXGe94
7w0/Qym2eZt5C4nsNncsQyHFOuDpHjgdtfn+bikizV0ltEEDehm0NVPNuvMIf6f0
e5TPk0EnAO2zrGF+t1mqF1PdGtYYtpS8Fa/S8RA02M2ULXklruqrpgLJD6HVbMLe
mPVMC6wCpUEiVMB9D3CI7kdhHCieb+YqPQJJvPNMkzFmNH6GbTJWouQ2WCGDAxpm
hpP6Dc4gTBgzwsatCapX/sPn0IeNPmpxQuG9dt9U2cYhPufGwNqnMfUPYWJCPNyh
ZMYXaBm6dDrPOeo8xOZfLKeIQgBL442RaK5zMHkFmpOhelp1AUqKf35EC2B08xxw
CTGEugxIv5NdjDrYx9Y7Z1U8ggh412TXpvHFUPSZig/pAbDP1xDUjEjkZNro4kFs
w9Vb+28otPMqCCQ/3IiYCdiZh/6DqfsnCux2x/pQhzSxWCsw/8Nh9OfSVn7ZLxI2
seYE3XtcKAADB6HLIunPkpZuBjirqeIEFHrDv0z2aFVcwPW89qRRZMDABfd4t+O7
Vk/IrFr6AEaOCmMuAyHmjIfcXZa4SqXmNflCuAgRYaXxErb0U7gq3pxTJN4RY+0P
4IydiKG34yAaEoBNYtQDWws3E+PIsamygU9gd07BNlim4OcfMUfOyX5mrEL8BBhT
Emfg219g1Rw+PxtASMfceHABsowAz5q03nENHeDVWZrSmHE0ubrM+Eej0VStHqvN
LOKOabmar4VblsftxaVjcnGVWkc3+taEWvrRHTSGNNyvkeYL4HjF0WUA4x9a7cGk
eHzCU++by11OaW21UmSfMSPm6LYjngjbed9QduAhl4W9+iMQljknkpYC+UfXRf3a
rJo0EbeKTE84UEI3KnJhU7QpsoCx4Z3OLWm7BImqpOkssbquntNGi+YhrqeVqwDl
keFsEjZtJOoDtdRb+A6QY8huIZ56zWCim4PJGrDs3yKkw5p3BJ5oy6OlqpokwOaR
SWXLPywlNhSXRVaK4zvQVJNt9TwS+DExdvP32VuS+LQJuUlE8kRAPEDeW2x3Sg1v
7lzVh/dzLD1F/xHiI5Qd1WH9/WwLmIJV/oSPU6Jzi8k9OR7RF/2go/6koRCSRAzm
WvlwC1DZd3cA9IFZZ1OzW7W1MtQcLRrgkiQXnI+v5D2ioN5C5+QQg+WEGT+X0jcr
im94p6UgGAW3C3iMeA8It3pgibRCQu9kui3r0QWlrze8mWT/1NpIQ5VpxQNbgImX
tKVqHRC60ijmpx2Mz660imheLmCooNDJfvF6/A1vhjVHa7hzYma1RKzTkM8jhpi3
ZtNJuLO2yi929bkmJqJ6iZjw0EC3k4wNCFtzaT6LwD1xVINq5iJIr4Bf2s6Z10DH
kOjG3/QBcU5taXdJreyeS9FFbqUzIh3vj6bKyLFfxbJG1zgxGf6vHXjrB4NuHUU2
mJrD1KW/UHsJSR/4VQHIr0lSVCXNn2jRRr6/q1LK4wdAD1Tbe4JTZ0egX6nvUO74
8Jq12a+JhQbYC+gtgJomb2WmJOra+g+TNaN3EEL85VvsPC3tZ7Z5CLo1Ii9sHDK2
IA6d3oBbGwAhwSozPZ1IhuXbPSdnpKClY48D4vapKdg2Oxtgp3/03RhCd6ywNIyf
PIA1HQ5ANyiVpRK7q/mrjvbAKtARgv5Zk9n/0bZcKbxVim4Ru62Ad8X7olVRKUYY
hM/wfO1w5RLAJO4BeT+DbJxtqEUHwf5U3AfHv9VwUK88fwVbtwCoWSvF9ab27TOY
D8nU6j5+GXzaxwbN2zgGXKk3V2/NC8bZ9WdbvB9LjRPA7t6BzgLFRvDAu0ZHjher
7pYHmCqQ/yIfcoKmxvqMQLm6xAgYAiuLz1pU3HHmQ4wNm0XqIzVFxpIHkVfeZF7w
JVxv7vtFwjKmcKPJd6cZwBH2KGKe2tOYnzWgruamgml22i49i6Fq4JJ9DnTiWTap
tTthFfQ6pxuPfkh7/igUyScVyMznQv3DCUIGw1CcKQbk8QZBPL1GFUv9w1A4jA68
Rj70fS3zlGULb7trKhPn5l5NqQCEHIxOV+gygpSuaZtZre0vXGPTcupVHbae2oYa
rmcrC6YH1yEFqmAtjx24ahh4r1k612SBPw79ymA1MvM0Ipha4JlMrm6cAypeftre
CBa6rM05Lwu4HvqDDSgJQmHOlDcYUkohD1dvRnZgSe1pYUNuw+ZGAojrQbVDsaAX
4z0+QjhEhidBcfH70PyFNY3tYN7yECPn6NuPFN4WECHf83QjwftvdyvBwSGTpIgA
IyxxM8xRiamBmJA4sROhEG7xEboNoDZKsbGEzGLH0gTLhVfZVIz3L84SWhctyq7r
uXGM0Gkjs4p+oezCBZ37fsfS28gI/8IimZcM5jqzA6sdA2WMf3f8+oztPuItMhP5
oDICn6VhEOym8OV5ZOw6/WlfhgKQyoZDRGLfi6RWnek0OSJ86OJ51PPvS6Eq6cn2
06vzPFrTM7o2CuvIN/NGVSSYoI5f+4c1c3jODkbeBh+0PXMVB6j1e5xPRIyiCok4
fAIjhPrxMpasuLhXOF892l8tfQkg+NXujASV1ycSVbev1ZlGgQCHzfoCthdV1dJs
eGRiLAb/kVSHE+EcRAb5q93Mf74YOX2ng+KjboEcaa/7e53K6/QMBfaY0kRgfjdp
FDHbsKHhnP8H2PipaTTRbWJH5Y7laEJeHlPA4fxUGjHkUjtUx4avx5k3S6CqW5DF
HgJ7UTaYM2BBpp4X3UYEq6GvV8NYbFvIMmzBI55WLIdlhtDMleNPwawwFORBPEYO
pJoGQ3saANft0JHjcfw3q36Dd68XURwMXpS0D/jpy+1WjfXBTk19hsiNNQhlWa3a
ZmJI6nm0ewFxV7NrUt/LO+zszaCBvd1ZFnBhKuTOUDAkZCRZk2vPjWQdzyjYXo80
v5x64bHu0EsteprRPeJRRWRbldz8B3aN6QGrJ9d3BVGzAWb4Olr85fvuEgvQegAt
OCHlvm4QYqH67poRxwDDZyVouTeKNb50sXTCZQSMupFM9MrnCRdxvkEPnissjSZn
3W81FGVkG98Cild1IApiZ9nXS25dCt6p6VCH0ojcSencQQEL++TQzOL63Ld1MoBU
Whll5/LqMiULQb7DvYeifqPVbC58NnMK4d+KZ499kAISSMUvy3l3vv6bTyoitRNE
xOdE+SVgJU2fQAL+upxWLa6dGuw/yLxUdgmZqIepaBdO1fOQEyTkrmIqyor+vfv7
Av7GcBF5Y2ako/ptlB9CaT/LfcGdoO5BiB6rZF45VT1eCNc2NEP6yyFZGMQrlmDO
qtBV2jfY7GCaX6FX9WGsVe3ZvRbUF84GZvuhZ+wKWF+U3pl38gAO3qHSHKwgMyFj
zkCyiy+f+yeq3X0cPS6bdP6jmEwcoG1FrbQn+A9nJb25JnC0VE+k1KRyARuzUpWT
QOiI1UZif92qkpNjjuBtDeU1VvCtILliNoV4nAUrPrZjJpFBWcU7vRnRLasmJ6cl
eV06JcrJp6aHjLh90pYCZmLMew8QL97Y68n4kP0ayxHxLqOiWo7nIxfYTH/gUPnm
cpUL5KOFwKiyORub36awvVa4vAlO2/toiKcs7XTpqAI/aaRFwGkh7uVQdc3iZEzc
qMtZuhN6CMh9dYZoHzmmxD6FvQ+OcrEP7MsCVmoLjvDCDpJN3Y0K3zAl8nU8cNyp
6N0wbYDl/k/eyw0hvvbll6dIAzoGhnEJDtg0MenaOjJUVY59vq3awv07paoI9H0d
ySeyhYYegE08N5HkYwPaykb/w0Ff9TqAgO6gUwZ3RD+4+ERRvFbUA/CoxbprazvX
jJd5oT24cPkD+s+Z6zRRyXg5LplUza9f/gR6E7/dOvjwUOiUE1EyHFs/Yh3NQtQu
ycV5HJestSzNz2qMitJJhtz7xQkxKjfOzlqSKHIhsSdy6hqbDsrlTRBiNvpioYvE
9IXHo/DKHh2PEE0dVUaSJUifpvbR7DGlZ2V4nLgLVSfX4XN0B0HqQZXWmUNgs0KA
DTxsRC39xqGHP05ePV81zAjw5C0XLgR0gcNZkBgJeBGko1YRsL/o6p3eDgjLGYd9
d45hZ49wCvHV99MNzdYXaDMOM0I1X2hwNAQpcLsx2uc7NR+BjBc8scJS0W2rDFma
/SGvBSwWPLkaSuDLV8jb8eV4keT97aQD664ENR8INZ2jS+jTro4+eZerqQ86mhgg
U0qySPHbyvoAxGgNmZGkw6XVDpU1eLV5Osm/685QGLQZETsBB89XO8UX6vJU4PVs
YfFDMCefhpGTyDt1jIhL808g4GY1n5rz+8tw7AhYpYdYHS6ZDUXnPmiPhYZU2f4O
s97QKrNy/mEzVK/M9m4CVG7xlcrAyGOIeyt0tworiLirFyEgnVHcs/L3F4ho4PeQ
aGjdILJy6NhB8El5pMf4gFLTeMJtb+RReXy9BjmOQRybTeaSG7O36j7hw8EabVv/
PNHMutlLTQqh6Q4G7/ywByuj+/New3WNNHFpjB7b4dGXyOPv8AJ0r4ZJ0/AaVqOu
8xRMuSx7lMe8nPaIC3Z6CvTUqX7YICZ+lOfmZa2lh/D3g120diqi8uqmgeeiNT4m
Fh/Rny0iYyOroEn17o2GmcuaNRlSodcFyTBiPwrlkb+Z5TvaoXRXozUhcxC3emDe
5t+DQ9ToruhzJNu1S4/KA36OPBBJLCeWWdI/qRY+jFpXBBK3hvvpdBMtKmX+RpZ0
7ED8PM/ULtU0Vx7184YTRo+K+nKdSC1/+kWR3pO7xbRUdS/DvHrOtTWIh7rLgmMw
yjI365eDlZd7jkxv/wJEF8CNXR3rHexfC1wjLCCAeahdIWKnhBZoxM7wgdW+QEoU
0/7IkjbcSmKdO/kxdFdhjpNUvCWcysRusfELldRQabe5PYoATjgotO+DWV35/aZj
YISD5gpMDypkh2NzeZTEIUBU/acI9BpQT3ihaKkEgrajKxVU0XKh9WbC4z4JpSMA
8I5L6L9EWAIBuRYhcEl7WOkavoZFgCmzfHBaccJloyy07W0bNV3Nk1IDvHHc90Vl
rm/nVHrVmvqjlcu7HZPId8j34VvlEELOPmh6BSnnRAO5Fs436B6CR1RptzkbE2Oh
hE4tMm9X47tNFAESn+UwDR2MgoUe67sRrz0wModblivj2rx2uhe32+AY+1ox9y5J
PYJULS8hwp82ohJO6I/gqLKUqBBg6d1hiZ259EBEPNBeSiwBHbp9jSOM3MMdzdfA
w/QnKfbj3hjvaA8+Av6ehV27RZueoKV3jJ49jO+yG5Vn1Qg3PZ4yoP8iGdtIDfr5
vNZrBKHgPwJgUvZeVCCzkIfp7SF1AReNCWsJbMwqXTORf56gQiv2r8CJvVGnCCpM
qVixdB3H+7u5UhEPdblWhnymh5I6mJiGI9wRZhjqfGI89Xtq8XhWr6JfMTjJUMbO
YGmX9bGgNVFtg6svSFdVDx9Go0WBhWKX310ShfpBViPzUwbcivuV3SH0KhD7UfWA
LKX4B6EyuMk0TZ4stwjMnTskjoEsdfaQTmyMVtVK4JEgulUF091GYQrW1T5HOmbl
p/hHDJzHpa/SDvDjlAUbkD4ULu0nE1zkrZ7HMyhQ9RyWQhVurIT9tm/CP2VgfHan
RDrotHOrOOSgmK4JuAi9xchbG/Rxoq63Qj4MYkJREA0e0jI7hvTx45JIoxku7SLW
tOP6zV6afraJuoBJotDpODwayy9diGav2vxX4y9StazWF6dh9X86V7yf1ew7piTq
rtj/NqZDqgtHsRWONSrOWot/sEdqs/oXXsEWMqPPfxlIy8A3v49BJiAM1oXwlxSw
avg46nJtAUm1kPTwhat5KET5CJk/plUMU2T/rtsQeCaZMtlODKcPX3vbQwPwbJqO
a/igpHHOlnoms3Mn0QRYfYW/E9lkADpnnLx2nSEgQH8bYeIOifc4NeXbjSpJkv5s
LwIyw4VPCo26RDlHVJ79ZM8Twtd8ulXpalcShW/BQW47xkF+IeV+jgGN9gLPJYDy
Uneaz+oZp0Onno79xdG2UVrGA66f1/aCDgzVfQ5fJa7gQ1hknvofrzLVuwT+W9cO
sg7lrueWdam9B30eF54Oth/SkppymWasapDWiSCCzX6nFs/zTv8ADl8JyHhNvTQB
B5P2e9SRdCbPZMbKIOqtnIvdkWBcRYMttO4y6u5uiGh7roQeQzr1sRnghyyUiaHP
6C4zaoXobKNktpsUXZGjT063Ld+uSjnOv8eCKzGMy87bkVkPbI+8+xL57bHJ49Ou
/wp4dQMMENGmR2J7MsWhW3L3dygW8XNHLzbrhU72nKnjCCF7NYvnb+V8BWnPCVws
8tRAIeoE0XLLuyi7SaUUQaRP4wbM7RELrq1QESFWxsxG0tDbaasU77YdOQQE7raD
zHdBQoWk1wxutW9n+LK5Bj9UvJ8K9YFjIDCWWkgy4CWxp6XAhmvnPjXoC4bqKl7Z
L/CVarXNbS2clW+OUFNl/jfBu4L6hSBcZICd6Vuh46rDw6vaT35tMFXhOIOykxZd
vbfHt6FcgzHMfCkmtgZX4+UxnXlwacgFhpFWHn6drV06MT/7Mbqc9ZFDF4bTMFba
RS8xwKOrwrJbN8OAJfN/a9MDKtMpu8yr61SxM5CXMmj/+GFLWdsaBIKNNLfnHhQ7
QTzt0vzmFn34DkW2iN6Qb3BvPpifAyOXq0cpr74tvkDhWW5PRHhukWZApy+4LX00
5NbJA12htIqSx3HurZPZdi6nTqueFePjPF5foqmeXYB7UcNQG/zl2E2ekA5dVghd
7e1xbuTy404guVRWBRneUkL1XJVZIYj1uZbAu91osZ5pp/kvUidBFFYb6uj+ZcQl
alRXW3b0cUq+Xp4E2ynIfb5S0Hcc5IqxO0HQAVOmKQBmgXBgvLl5LHAGc14smjtC
CFwzwUGx28F8AyfDwckTQzt4l2PSIqVCyrmYB/dK+rCcc/5UyqW/2ltrv5MjPVPu
GSSTaOTici3NhSeg4waxLba27Q6vK7QDcSnoSheqdjd6WNaPUZrF5MaHUymetjyt
EBTqKK6keI7YUrs30ka03ACaa5Quee6fSgAdIXs2nTSs1MdJbjrBo0H1eq4f8XtL
a14mRC7Vbqyl3gBD6PLVNdvhYL5QwRaHl++yTh2eVVRMjGoVtNxyaCu2sknH/kmt
kyPJoG89zQOosZVzyqdSh9/TE8O5X+4j7S29xZzlPc5x+qXYGsih+Hae8H0kNFCj
HMwaHmDyRPftqaIzwe8MGZrp3OtWYj18/iyxTYz+27uSWLcGWZsfs6RdnXQ+Obzf
2wCaX+4aQfSNfQIY7br0Fx2Tg70Gb1rDaly8I5hsTZ0LVP1X5WMaTj1t17I9P4iz
wJxk1QO4XzA9vQ7Ys9AxfeXwsxxI2xSIqXsTtFXrJXLBpOm74UiwX58MyDA/eOzW
2v6FQtY4TiH9jL+cG4ota56rcJkp6MWLaJ8tCM3e1SRJs4YUmVRx4eFVw5PabYB3
Z3qU1WdoHbqBLz9s7Oa7cVWMaeI/rcSg1UsOwEvMRQkIqcb5MZXZFreFvyYGnWY8
4vm+41YtvCLL1nppUs4TuKKdn96PP9OhD4p9Xd0j+DI+TWN/+C84s5eYEaK0ijmw
R2Y1GHW8gREboKK8e3fiAKjpvq4PniK3+zZj0n3uvj5WWJqR4eI+gI7md1AzvEZ/
HsAJC1DEn8xUQVR/tACaIa8aJJk1sO24sToB+EeM0bnaSsZ1rs8WDVG+3zBdvEBv
i1kl9jV3X3tt+Nmi5fcJTNGe1H+H0j2RZF6L+Geunmfiu2xI+uJLfGvg6oIBMhkG
UVe+I5sJgnIojF2jaPQ1XXzujNB4dUjK3T7lvobI7kOO2BCG8gCYtBDgTOyTRRpo
DT7StTSSx37WqR6Vky9x0BeoSpZMk628MEaP1wB5Ov6k4250gVOJRqpQzMJlmotD
I4NMoSrX06t6oZ+NREwSE6l/lnh0Wezk9uf/ybqtfjPDUFTSYvj+3iLNWOemcDrw
1fccSnF/RN07vV5vSWsQL1BfRRnS9rELMTkq3tSZxNS33rahGtul9z9mzteYxhsZ
c8N/dZ4FwABTTkcgmAkbiltSwUxao4BDkHFqBuyIAmu0+gUpfvi8c4v++4+nd+s0
Auwf4+Yk5y/Eg/vDhm94XKvQ0qTtndVYTbFFUp/ypYhyhIPgq2K8sHxp3JrjoPYU
GIUhixcIJmGZ7VRql+gUXk6XMI5YNHubnNoguzhWcbDoUcNst+nTV9KHHLW7YoyN
UEZqjfcqczzxd+PFLeJWV691lU4gcrl+ToE8OVaBs6woVpn42BtY4Qtt9TLkfo1W
pCienhYe5EDL9RCBfAwkdDoYT83yx72USZYAOp74XUxDbvhXQb4Co/xKQZQ4CSlM
8Y9Om1ZB6fA+0y0zpBCANCIMxpQGiBmQ+n0eZec9D3NYUP8t6t1+KTMQQnlASuCs
VxpqLhEDRZXu5bVI9qe6cxw+lQiLCYJykyvTyGRxR99qw3DEqRUpdpJHIgmWFGsG
oz0usaBwEgYPA76wHLAO1YMuvjvsUU3+tVokgE7lV53sJBxvLP9Jl4vhaDMC5SwG
teo7Dty6EIDJH0YuvJS4VDM5k/vbGecSO43Z/ZhMogArll2Kg63PXWGEpZzUC6pi
rT5btqwygZKLKf9bmWK135P2fqg3ojX3PvvlN6KHSExRVBI7dLv2vQmMpOo1z2to
HOYcqdx6fGF1Rm0b9BckrmZSDNyR/JaPLhLN/mhp6i2sJNGqJBLFi/gSXJmaf8MD
R3Ii09nwt+IRkKDd5KBFHA270czW/Xr/O/MEsueR7koEc0W0/XIVs0SY2zfhlkY8
J4Qgl9MPMWgf997d0nw4iOpNOil7QkPdtU38QKhsmDaUXF4wlMmtaECv2W35LYYO
d09KUOJ+7Eyq4ZZd1+5ul5TkxubeF0JI5mE9T1H2D4YuXNIQ2LhDEUgwKy+Niavr
efKBEwb4FAeWf41IZ/FsWuhFscDwMO1gzHwAc7nO3lg6YVCHwgUMu9tlTuN76Z4w
U9qVxKyqOl48pbzfEBNFwGBgVUBx/QwMIEnKuQd5FwC7FCyAXmPDejoH7HtZOeRG
9oK3rc7chP3EqfkPYwT1HHiqp6/O1OdWebErqvQp29Fe3WnqpPjir7xd7dGLidxL
D4M6dJC9PRdcM+6GuSrECEYWbKbWIXysooGdM/v1TDilLS3d/WNei2gyWkZ1tXA3
UluU8n2+1r4GhB7t0apNWK/FqvbKY/rBAeMSl4TqK2tC7HfmTDBkP+3asdIryrLm
8cI1FP7OIxPcUidPUhuIjA0BrPvCB26TVhoqzr6s1BeBrhh0aYX0KydULiGy5C/r
v0X5C/eJ83W1e34N1vKm+qEQSbBp+2kQstRY1SrS0kMKbQbAOsKkNUhOf6vU43yQ
SKJjH5QHoMnd+nLDQjKP3whEbAF24QBOFPVTtuZ3e4MklJeyXGaMezjide/+X8OW
WIfrK61E5cPnLakxfaOtcHTPP6AssrOAEHXXO6+tufomQgm1s2vnwf0KdEtqzUFv
psLHGS4qQNi4vI7N6Zy/QvMF0Viqd5SBsn1tkQWEJFu/EqWm1PGnnfhnISAej0HE
WcpmRPPDa+S9HY065Lscoe2zI9GKV7LRH9yfLh8DswWD9GsaJ69Q7PeCmdOHnFBo
zv9yY5if49s3YL6mUZSISj8YwqlJJwr0njBB7/oum4og2zLAsw4UEgdCek7tsQts
R5MHU1QeqyOPNR4pUFUh7jlb1R46SKJzgvjfe55BBlHGfcZBkwZCAp89QgZ17Tgn
JGXktiO24HRdisxNhs4Yk7bBoDKcdmVdgwQtDDXS1IP3+gDFZ0/0JSyHo8OfDuaM
xQv792jzlZu3pSQ7FTySrNOym4oLOxvYm1UoTHmWGRFZ5bAs5fjgZV9l7RzZSUBR
DZH7iTvytJDLEo+0eqizcfDHsiOUJJoelrekKOk/yVJuznq5f0aZjJwjR45g2Yag
chon3gPszg+4783uiYpf296hw5JNNr11yYVioEJf4WZnxTsHixw6YKNovoMPFDAD
iMmW5+nqMKAuoPgGk7fWKu+osSeieuKQt8Rw6Anb8GA3YPQslY0GAXfxVgm4RuNQ
5pqPk3dhbJJvuqUdW9ZF6CggU4nE1YIomjqLvFi4ptbFlcH89j5iAS86L0Y26HxZ
DnHXd5Sw+JauRFuHrajZpu8c4ZTTbStj4iHPugc+tNTHcKvsD0t6h5wvyZK9j1A/
ReXJP9MQNnuaS9aGcAEDkBwpudBV/jYrPGMDR4y/RmrvhACZ0coN9BkLX84732Yf
SAuKwSWW3c7BaEM1yJz1/+ltxstFDB8bI/R5xbt9/CCc1egt/oOV2C+l79jIlxQT
YcATQgU2kqtCptsE2IzPvRRiepMGYTvAgfJPlE/I2xF9p1+WH8YWkLJjBqURStEU
s0CxwsOaN5Wh4qC1QnUQxA4NRNQfvV/NmMN5FJyFmPD6ZmvwAlpzw/aZuHncsy+m
C9Lvt7ZlgFTYgBZQJ1FCmj3l3sIQV8yyyURAptSKGdhfhfnbJMGmVHTai7C5e9od
FwEfb5MU1BVhcQOMNJtGREX8iLpd93tqa+38REwb4iJ3v6vooHDxo2KJrYDU2MUM
ddar+45r4zAZ3lJkzH9z8gF93WG0tBsLnEQsM4faPdNRWLquzAnYr1njV1EAbH8U
1hY1iQmKRRJ8p/Rm1NGgwNf19K4w4gZldisc/UmRWbvAxlXAse4ZufGoSyuLO4e8
9J9Mh5DHlgNIRU+zguSWIclSEKryQxaqfiYh7VWTL1oPse+h3HANzaY8LRXkhQzP
/HOLs+0ZKwnay0f8Suq+sGyf0XZl9doIZGU+wk2iOR9d36TYtD1PTVVmrboibFxV
jt5f+dy+HnPANv5Li6PE6qm4IVKeE57K7zaIoVIdq/OFy6ba8I5nThG4mpOQ12QG
6xRfGWxj95ERSxzk0aFjUaz4l6F6OkqFAbyGVdyNA+MI5sVG3YZLEPet4hvK/UBB
7eX5fMxrEoENRAnnO3MJYGPTnNx/BlauWdS+eDX2YQFekRl6aElacysI/EQe/mgU
CjaB341QJJ09xsyLo87qUAplYPwJ4vtN/BMELP6w9dBCeh6gS3ne3eMeoiC97rZY
ATSP8XNXlGEmlqbTXYfxx0na4O6TG3oJ5N4PcwkNMlU7xyC5p4dUXBtPG5h9hDfZ
imtxxfVX8oJkFhvcBnlkXZBz2pQVTWbjREWAPnqv9eUGc1yBbLyPtZwUYkNO601R
u7jD5QJcfRNMQ139nt2uZye6JN/DVRk32SjRgU53Qpa67gAYapwrMrGDx7MZ5eUN
pFpJKBGjMJWrESN1rZbEuxsU3d1mt7pCLC4aV46sY42WsNhawvFCiKW2fB9ubpiZ
lpQIAC7zKBGOxa01FNhyqUDk/WgHnWIZmKEZeihaBazHReuDWS1wOpJnKXDP4wpf
O9Rdlb3t55ejUQoXqEupuoJuKdPmxIubcCIn2FGC3d31LS9tuvvliEM+bnWc58Ob
VCfP2n5uTEVU7QyRO1SsR53o+YjAOizggjh/guImKYi/wnatCBibROjTpTmOg0OG
/EyC1hWM0uKVOWRr+ErWetGh2X0z303hQAHFDKkoQGL4Gbxa7pMNj3aVdSaqntSg
woevrkWyQDOw+apI5UE+sRnJ5859fwupx0RIQV4Bu+DJEJboDk/utX4KfG6FbxA/
wssjuClrnNiYb/cMY6y3MTWZzQWBuky797qqo5WxFi7FAmU0PKilgf6dkj+2IUXm
QLQagrQAY9G+r4zNJapW9FAkMnTFaPs8VKQUyTnrJm+hIssBM8tCkUI1HJRyysZn
9OyeCuNd2qkDkuiur6BU293Ao4srdi8def6aryiixlU/8DorzCjG9hSFBM/itZtV
NJt5NGWLfdvSoVO3/6nWZIAwj3+MG9Nl5ClKICiW1B5qUTJM6xAt0scrhJXtukh2
eCJ08m6vUE4YPX/wEzhleB35sZMfEVjngjm2p78RqEFpigaFQMS9gj6I/qsPywfI
vUIDBCtEesM+IFmqeVF1icIKzD6MbuBTRzjO+gRjxn2WdywIjldc2ovg5lbK012r
o2YDlm3ICFnATs1SmIW+qxmAyba3CflpaS+bE4uhmx3smErwhBDyJyI38ikYuNW6
4SsdliXvfPAOa3MJn757lWLRQxgmpuc8N9Oi++Fi9nLe3P2X39/t643SXy4HD32w
hR2rFWJBbcpLtajpG03dTUOqNvrGmp5PBnL4vTuEs88qTmCIahDnzhdsq4WfjeH7
hMYUnjoNASfiM9C+wHwKoU1VR8rPPiaCcf1fc7uKZfeR3IIAfz/V8YYL7a+bQ2Ao
5IPMG+ttH3CtvdU5fLOqoT0GhkCguzEjvjAetN+7swEDQEcF7zFndi5wBIUDGMRC
zKus5w+O5VtNdfI1Y1lG8V0dczlqclobKTvCSDkeljF+Wzgt6LaBgr7p6oa4+RgS
Bk1oI3cfUT5TRaQrJjlqan0f4Z/dzjLrfpfu5BaqrQKfrOAvdV/86LYGhrrkoOTu
dkDMGcIfDUUhpjXPqJgteclgipGiEWvT1H5qO5oQA6FHcRydPlcSkKGNMX3giQ2w
2fQ+ee3VzLlTElefS9JmsoLQxh6KFqog3crfeAR+l/DiOrj1JzDqs4ga/OiIS4rl
LLFH8sGS9iUxDpLINhCtQzwq78vX3gzioakxSOvhcIYvoU7XDuZQEqBd0isM1PUA
nqDuqg6vK82rzu+vWQE8FrH+jbvNdPauTjVXxjCEB65Sh28OaZRAygjgvAIU3r4k
tKLjvd9kAPjPm7LNFMd/YMB0wmbzKxOAxvrHAZf2u6N4y3tg5jaL5udWLpxH6Q0O
LxSnV4oh29y6sTDpUVSH0kKNCGYr1f8T1dLAHsQkggX/F5cKybb58gtv7dAdg3oo
/shjdzWxwj2PbpVCod9gfTF9J1Uc6tCG/vcFM9N+rzXAKf1dgiVynrCSrx9BWTRA
fgbXrVf0EOF1REkfWQg+H0NqSXM2zeMdj9AVeUs/am6v9IhxapoOq/E0+BJXK6kF
OgroO9+izKiURhGBMNq+qe557EHQTbW6CwQwK5w2TkANAxa9S8yt8st/rdVsSf8Y
8lkhBSJDnxYIzcyPne3X/MfkWUMJNv3oTornlSD5rD8S6UPi244PoJh5gLEhay8C
RQ6FLcPG9WBrt2rRHD+PB4luhHj8xxxsHMUptiu5Ydj2ZS67up3FsQMUzPS35VuP
pHWfqdC9biKi0dB2WDwzCqJUFeFrppQ/qGAG3K3Cssr5Z4mtZa6KdO0bzpZv4L/u
O5z/ETWOzBzQhr6mt33hZDyYDiy09/TAwN6WRh4cANtMgl4C7BZzGRgv/ioQDMV2
wTEuW9nJJ3qcWY91CaN2+YT8IIjsHAogCGYb8IP4z5N6ffD5Od0zX1HkXAUjqSKx
FPAnFVaadfxvuYtARGzWTAK/SRW8kHtNsYMKc2f5wAzO7we3ujh1jRRDskB3+zhd
18ynupzobghWgIq4fzrvUghLqXxl6WkQUxPeA+bIjxeiY7cAfEilksCVEv6u20lh
LbHAQdBMgkhN4c6IVUlmqSLAJYqJh069FkFhk8DnPfPy4/1kBKnfX9CjGdXX7wg4
Q7KMsUf4Un+8lKL/B+B0PVZTt6/AMw1K9cYSJqFkKZVNpEAC5dLXQMxDnVe9AASo
HaulcP0kPZEOpTtvItmGVCpbXuXT4EQY0Q3oqonfqbYDWefC4uSFwgLQiJ+By281
9RXrdoKKLeIHWKIibQHoLPpkRp6LcWuCC7q78icHva5sA6YZ16KAvO7ePG/JojXh
uwKO7/o1nVA+BUk5xsLjZwFIZVfEtFBednpu1LgbknGg+20vhC0KcLLAfkYZmKg8
yDyPYxngg9UY+DQ2OsYibrFfdVo5LnrI6vFjWpXTVMBNjeGiu4lYp12sIFtH8v9b
LERdbhlmUapPR2whMVU4/2bU7Pjpucr8jg0GvnCFjkyC8dWwMTM0iExRRK6aGJIn
05ZIcYb0AVIVctZpVItbkMI7BKb510Cik/sJ/OczHKUH6IfCYssTIEc2MmphJgEn
LfZp+taxSk/eeMw5YFkfz8o7MyYXkLNy088+9WnFizg8ojaoOyx237GkazrPPotN
JQkN21VA64/HxfL9qgIvMM2MaLLl6z66NnVBfKXszCYgcexYUxSWnZygD+iU0NTT
5eN3ObksTXvb9/Q7JxV70mmGCH7prPenmWjVitt7UjuoYsYux14UW7L0nw4/CprS
Q39uLLDq444ajfvLxOkOTANvHf4JprvmsXqFM1wgFnhfK8qQmAuu6YtvNbSOllBD
MKKds+DMtn0649FNJB+vstfCaMcXqCQ1IHg/GyHsibeOszXDq4pfrD3VGO5iH4C6
c84aLDx0xDk43LmidexXa5JacmqSQ7UtEVpDH9I9Mjx2y/9B2FxgnG6mCqkgv9DD
5eKAljFNsp5pQEvBxmYFPrEMoyuS7kvj8krSLoCas7ZbMm7QQUaLJSZCH7RdyYYs
4cCyhIM1K966ob0AC3NId/+dPrzmjyFgyjEscFRb3Avl6dUQDipA9C1N3wE5reUw
P1bFhqki0eGCYPCVjC7uslLR/fXlKKG0tEkmqc3ka7/wkv7zpMCP0fES0uRp1n6Z
P2Ha8oav7Sihe2Aqqabztm4amvxx7AMsgzFdjY0bzMoo3Y/ELZARVV9yCL3fmhmo
OYaCy1dwLxpsShC4/HAW1QNYr2H4skLR+aEtyFIX8K/RPVp1PVbeyWpgirV+n+Fu
4zWa3sM9c4cGqZFaHcwJIjUnEp1CIUFJaRN0JArlnTVDmDMu3ggGtH5IxsbGYjqm
4VCAMil7vuiYEaoZYbB51DL3D967DYKaiTw4UmA6qb9aK67EP2dpIARC0jzzWtnF
5+6oTLOkEIv/ATzFLpocrBU4N1uptX5rL6wOxQ/U6MCRNcn9aWLpKS8eiEa2O9OF
9EUmOQyPH/7odSTZnqUbkzWLBy6PV5J2V7EyKeSSvOlB1fCqStTaHb/Ow2guspha
RpVyzKYdJHIg8V8om4ToL5Upc5QyoZJkf/W2PWQg3MDtk8czz2KZZ9V4PbfOM2iR
LNJ2s6s5s1EGsQi3NrdX8rpoJd2XTWS8vZSdO1P8uVMEM1VIlBf6eRhnhTTqbENm
wetYeFDtZP0PkLSO3eMDwhvAPOd7gqD+Bck8qY+hC05d2n91j76du3TGnCCmS/lu
/c1LudhhTa/dqeE2u0XTu/MukBwT5zXM3ZZIQVKhiHVaaxz4oZqZHn5lIG3v46Cv
RV+hH3wNimEisFrsWEu4UCG9FlIlHqRQhAfWAyH5woBCzWtmnE8V5+PvzNPqrsYm
vdIKDKdUeRW92uDC0m1nEnszZ7gfvZpOtvJrPBwDko7qq8ekAnjTCOL992W2s1xj
nziuZxGQu5r7slGp7lBQBUZQBO6BDLJaTz4PG+FgNjJMrlYV31XzLWzQ28WmQwkC
HMirbZWWz2qxqvr51TmLfC2Nm6L9SlXDtd3/oOfOqyLlI9EVDj9oy1fDKuFhaoTI
u7ldL9qDC+XNWNyScPnGULYMfzHge/8XNGKQSAvQRdLpOUUPIBFF8D09MFOlr5ly
2tivCB89FFLSKOU4Qxwq0+UdpzueDwg3SFXo2QBTDmPq1xoEPWr07Eh753X4aTkC
hCLVPKcQhcKEka+1LwWEkcHZH4+y4/5j0YW0xTF83aS1icLBgZGvovSpGcBIa/Y+
+1XFPf3JYVwnpyankskFKfPRhznI+ZOJnN00uEWmUtODU97N3CWX+T1gdDBOm+y+
rq35XYTIz7I1cPoQm30oXOUcf6wCQPalM28ttg2BoRIp3dP2auDXRykZcVNeqb8O
2CW5HxPBXn8eBwIiNMikjFRwsjAlB/5pFt1jL16E+tBVt9RBo/UVkbl/8K+QEKc8
HUinvMkoDi63kuNG6uYFlX+C5VC/2YEyhG2kajD0rWl53LURC72SBgsARGBzRJZo
zz6PFpMBHdQiQRVDYRZlYGHTXN6+T2djBaWHR9H9CdPtAg6WLmWvHi8Z+AmTzKlB
vKSisGYmdkpr1mZ+wWRhapdM3jexWCdZ3eeWXxGtNqvo68EWOudD8seaOXOCbVSo
rtB8zovhdzW0SrYMQM75qR6Or3f6hvzOqYBQqnafVYB/knpBXR6zMP91N+qdoxwT
rBhGYvvkwt2huKl/6mJWrGdacX1yMbe+R3r9DonROc05zrBQh9s/l+/Lx/saNvj8
g+kjlBPm1nCkhw5PJcWNi6rsYPaxClNjGgoUFAfZK1iBduBE5OwEl2IRzOTxbpdk
skucXHW71xHizflUYR5M8oeJOeIpWcLjtuaqLDJa3GyJTNCt2T6oylTiy72LmROR
v7vZwohi1JSgv8oPLSAmMk5w6oiVYc8C4ZngLjZbv/EcnWUJHZQUsEVAwGxowQDA
cIOHR/wTqid/sBeGxOQc3/o45AWf786CxACIzvdYW9dGYkeJmsrternyWPobhbpx
adwEWj8aoIZ5vHd3BEL6d+CWn33dYQFkGQ3TA+1qfWzjXF74QMXFcbPk9PVmnxmK
KArBABo05zrlWwNSvO6y/vqTKMv3iikthqczsS/bKq+ldeUTacCGMCACUby7fo1Y
DIrC/cPszNV1ajeQLKh1Zcc4RepKKoRoi0JDpmJ+O+3R5dPyX5FF5Qxa/jBG5Y8r
tKZcwq9HmUQY3dUwNcSjRjPbywefLAA54cKRHre/pLda/n41paQ+Xfibj1LTeV5U
avQ4xMP+FM9OjAOU/tGtf4xHVcjWJbU1lk2U/iwMoKwsbyskkkjLJCln98qnLAsS
2LAN0yG+tcjJ2KdusWeAftol2E7edqe4NbxYCevguwwo4l10DXy4rSsptiBRTEyq
DCEDQJiw/flL7u5kq7e86KezQwIFSxwQiOaw6VSUPyJUQf24POyxxk39veIaKQc3
sAU9fPHl0WqVti1H8EJInHp1hiqLvTFI36CrP9iUIj+x6E840KtqnGu6TrMrkav2
0aXCTdNY5ta9QcaxFF0q7N0kVgNV8gmHRsC149RyVFs4HzblawUX6RdZqqT7wwso
XFN2xNS1Tlu/L8+MgrC3tPa0Mm8rCaKJQO+clATnt9Sshs8Fx7+v/4TcRL3iHzB+
3B8r/13OE03cGOBxHpGKdt+ls97P/AzeL19eXeb7TsunFFtT5VN3vOA9tsUsB16V
Gmo45xpuj9/7tLsbhaJ/Zsj6WEnYwmLXtZBi3NE2OEM/rpbPhfQXWyIWZ5CIcC7b
3ChNgm+2+3gD2g++zzk8jTFGRIg3OqkZ/ZJCms8POfViDrlyTmvkWI0oNKu9L6dE
8rONR56NSbHp6PaUz/C/f88cgvDVinETf//VYTAWeA4yVkOx9MAdcEByBMOYHRdY
Wm6Mqmkqke3rjKm3Ky9L/guCsKf0/qK0zL3Ga6XwlYsOdaKn2uF3fiveJHRwzn/O
/fchYT+yeHOExagLZqWOfb3oOHpzrOUNeBl562Tmaxv43DiZ3NpDS1ju+eZcUT3o
rzuPyyfaHFzRwEK+rdeFyz5OzdkBFKjFP3DCJE8Lzq8o8v/TpOA6X3Kfw/fJoi0r
MepkbCgk/duZKLf8JpFXq0jee0CueDaGxjj2LKf0WYw+WmTqf0eG4oz8zgwddbbH
nwnwGbnhfoVMMLN6uLIsy3KCAk/b4+aL4rUlGI/fbsp+3h2Iv956PHr092eXLLay
7gGltulJX3+ziVmjmkKbsHebpy1DrFtgN+KA116Lfo8AoAoGHlKGRjwff0zPV07M
maMf+jyp+BJExzN+jXh7/J1Y0r/FYPpqdmBFMYbhXlk3gEJg6N2KvKyTTCIxLpFS
oXJ1PrYOvaxxZTKKMbj1bdeKVAlGRMvSgds0TDhRSuFOgAqYl2ub612+6ke6RU8b
z48Kl05/AZf9SFazKEXvZ2WdH/xrzGomAcWflVu3cuz335Lcdko8yn3DY62u7/dD
fKLOvVPPk72HCC0+NGtZSFhSVQbw37jUp7huuRsPHFEEWORa2vMSGkoaE82JkT5k
r3YBdP+qxXRmi7xylxLNQZKXgW8rdJN1bU/bj+0jD7VU2LW7EttfKOJgs3Cki8c2
fxnztchUL9RJCdYPiW9K19/T5gebgtJ3cOJj6FEa8ev0r6tZObkoF1KiLchgx4/8
0MKLDvGdFS5FMY8Ll30AtdbEXkdxsswgfwox1eeDIMwdlEyy8yfVrlMlAF3mccXj
pwU9RlhuVsV/kS8EKMVEhv6njZMo3IbqzgT/1vcJnCAfrVH+crnvajO1/yqOT51f
PRdzUepKiNB9UyeumDSUv4S8VN2osI0X3nAqzR0d7DvTiIcq4FDUoGVgXz5LpVQt
ISIMZCEJiueuJA2Vd3NbDw7XLtEC8AjbstYUnU/4744jFdDfbE7DvC8FgkAzuKiF
HMPMTbQD9IpOMhZGuJ85uTyONCY8jLWqznsLl3//DMF9QdbN5YPQLFszl25ijSOP
osig5Wlxdgvmdxn7fJyxgLuJdtO8uNO41HnDA8gIyijtDpXjncCBLXcF3KNIXne1
KF22k0SH3TEZfLgI36z1mnOo/823lX1G4IT5Rzt4HBmk2mi5TOQseSdXiWO4xVl6
r8TtBV6eDS+WO8g6C+Ow5ZaIgXhRrUHmzuFlLgoElAs7gsdikF4bPmABWp/WsasN
OyKYQojMlNSw0S9fU9Sw9dP5GjoDQ2bH0Y69FPoGc/2/ooID0odWyIKcVWylNJt1
v04Hl55WxQQTkMub4sJnyi48mgfcQRVS5WiFsx3itjEET3CMHcO7UNeIQhR/teYz
5zmT76s3hVAFLMvVRKvCd/fm7vVWnM+wxx6vh50dXTnjOi1eFZeExGrzts3h7t28
RPM40Fq7/VEKPWfksq+Shk6HYFSi3XUxlw2aC17r78luGbWN/xH78OCwrA3RHEli
3OM5yq6xNBeHA4kX0uTCJYgEQaEiwjnq7nZZxmEw66H+OqlGY46kDaB8bWDmvM7z
GTdjDJFp4FFYPOVPb1FB/VrVqoHkAJXsTKZCpI0WJeja5MuA7LfdRMoMZdJkU7cO
qG1O78klsggav7gChtPiOO5zBoWmh7YejM6oKkzQS+K+qXVPisT8G8ii6nQhxzSS
zzVkqF9OXdZE83MsMtwFn7LN3BHjYgb0qeAG8lO+mp3Ito3Uh99vb+H0CjYB2/qC
B/0LOkChaaw7FDdEvhLd6gfZnuulV7r8ez4dLE1pvHFZLIIF5ELgYBSXYyloZFPi
RlMj2wLSNRgo6CIUeBfgzOZs0gx5C1n9WjtTpGFpb1YknYSTw7aCjQOTFdt27swB
ef0RGIJo+y4t0PIKD67M8BPI3lGEEGtZbMphPbnjfUQwAL/BvhkhxlXiMQRXYK9p
AoBCkCqxW1ONhFvRKxYCXWhWOJZVKtMCad63c8akAyM+r+dfuE+F2CmIBG9yYWyO
p21XWmWUGdLwRI5y2rAX0ReBfldnmI2I30U5R3wdlsN/0RHbcxRjwqBis6M7c/uE
tvYFEbRseWFO9y6ok1NZ4G9cSwGP/NJtN/QczQgre00KShBN2zJ8n9Ju5p6ZVQQU
3EUDRS6zLQBzqioNU+CpCBwvjbLWTNW6hjVbmRff3TugyO81r/lMHe6zHuu5PA3/
WTjyW35yyQ7oipe3EO/x3Yiejo1lW77dK5WXTMdn8XPUlQMn/nStve0R2vK+vHwD
/0TCii4tm2ezVhcxGUEgw6P5P2wWs5gR1l28uvLnAZcRxArOJ1mqrejkmuhbzWfJ
cp+7X0RoRER86OLX7mwatIysdulUIrfye8gL68S1nnu3EwqlZaQpynBxtvX6yg4r
ux2G1oMMiFiKcLGgld5ohTryZ1WjuGFPPe6WZXhXrLEs0VgiE2vC9iSRY9A2Qg/H
syjco2BWr597ijXGnVY9Zt32CEgUXuZqcy365IlviQrjNRWyQF+y2Rs6rvboYDvE
dWAJgQx3WPDuQZXntLvRlsNnmX3gomKiMlM9WR+rO7/2HEX13hb7nWun9H0H3K/S
HrS27J7VXoMzBj3K4i18lbOS4UjDVP1dHNyPK60Z8CVuCTsBZ7qNhxgUb3sYZ7JS
M392yj79SXRZmq6Rbcderh6iZJLEqaGNTh531ezoeFFMczsNhamnRbIVpc1D7qfG
EylpQ4fHYKe5YQ1J+cJJj5+h7RZEXqk8F4J76tWFhp1Ar35wxpexZXa1vEctOpsF
MYdFX9wbxMPnZ1TaH6096DCKC8kauQmrQaZvTJsjLLKwTHdykgflazDLPLcN50vZ
j59wmFWqBKMNCRWqide95Yz63ABaAevqT0jCCCTrTxnTra+v5Ze5zx7UnRGoI7uO
7tz2XpNuHSyIYNlAaU6H+gdqYMXxOY65cnHJ0s1cChCtWiTSpHsHPy3QHHTRz0a3
ofM4jlQonrz5+sgd8O/l8WFQJl58rDpr+PxN7Dm/23laNFkB+4EfsfgDx4hnJ2h2
/O2a8CC5RZKQFRFroKEX3qfFMI/If5BHZsNELch7anVdu8Zjnjaw+6B2ES/g75Fh
zDAk+uryBUPF+0Te0SVXZGl/889mqlaKJrkZk+mCRYgjiyin/Ar7eyLj5zH1RGG/
mMN7CYj8LYkXi3hqiqVtGLxUMNY/EYtWuE2FhEvM2hsH7K+TcklWQ0qV44AUIJps
CvY2a+bsVwFtu7e/Z2izv2IbYnH1UpbKvwikMWEmzwvb4I2169lgmHnxM2DnrvuA
s7dszVcOWbRnCryXDB027f1urUBJ1HXPG35W9UCQUwrVLYh1GWsFcJrttSAyeB7c
7eIfF/zcpRdolnmy0uvq4KUzY+jaDDb8sBv4xFpatAPvuvtEVjkN5TJ6UItSHLvq
ABYqxbdRxO4i/5Bg3xj7T2ozhseZ3b4h6M9Vx2Xlb6ZRtSfx1pH3OUpSyIU35l2M
/kOkPmXESLzBEQt5c8nQhNebrzox5YD0Ivm7cb2V+4CbruX61+z/kTZb97oK/p1s
NYxlXyTcAuf83Xx4ALHMhYEzclONrFcuRF9hWY6IP1NdFPoxJxGqr3BV2fCXL1C1
sCEdwGnkjEFjNTsdGbfsb/rMDIwX7ptFPpOG4Dj8cGqT1EbsJCdViXyWA3pfQGUO
115UTnMlKL5J/c4NYMzPiC0YBCeaMf5pAdCA4nlnp+l4yoI2z8E0JwCVUi22JFTl
JrTycBdjWF0YrSfsirFKljSFXfeFzzJs5FIlaUZkOML1azsvf9P1vE5+lvix5SP5
5HzViEzmrYu45xKCK7CTD8wiXYw4zaeRoNIr9oJuLXgSWmW3UGdVgKcgaViNGBRN
URz5mkUO4G1Wf9rY3LHSFWoQ162OAzhMCe8IXMGCENFiK00Ti37gZOrfpcCfA6zF
1Qbfp6HyCHIDqRuPw9PMdxE3vwm37frM47y5bnL+l3wf/WucMHLWoTtpgG6EYs4j
kVS/lWIv5urJcqIpGdiae7OpIagUtPl/yOPSsRsEpR3MBxNuG1PRBMqStz+hdPLi
XXrqS7rHU7V95rEx3Awgr1SNXtlvm2uGnLCJ6QGAWiIGgdqrOKQAuLF4+d1M4ckY
La9V5OEs3ah0gwhL8sAQ6JmbyBDBcwYaOBM+4u8wy/039g54UR+MFwB1r/fosHF3
UYFKkfRKkfuPmRg0esPJM4CWYWEFCtV3Vg0WHbNYbKukgWmywuqxUqg6UAkHaYBN
WdbcpDYxCUDeFlzsqi7vf/wK1RDF46muKmMVJAhO1V+n0FUZofITG2fD0fLb6nEt
lsR/kZdQFlOU8DJarpDnpQHgRa2UbY6GkGeMHwkvVK/MHOurPl5bZrj9eigipXKJ
T2iKjFkds70qrcxbm8VcNn+OPAi/kEnFuNjhjeMv3M6qOd57sY9pxU2cRWZegZ4R
7uPlWU95mntQ8xeWcFTd96ps7kBi7sPUXQaCqUphib/OPVtGMQ3777mMf/o47NvQ
AIcZ7BzgNi9mdSleVZe9vEZ0RK+Sj/l3paW81Eb8PHJsB8tzQE/050KDdEo7mfd6
RSqC6WO/zB/aTCQXb6x4nZMJP1Dm6dH+bnNiFRV+YV7ZVBVsQZnQ3Qa4SH17ol6r
pR1WaotBtFwyysn7NH65zAidNYIUBcnjwsvW/zgFTVUOjCtiUkKuCR52Pv+AII9R
R+1oS3MBgr8bRVH8hi4ypKvqJonsVcUm/mGBijQW1xtRmnhVkuo6S1M7WOD4omh7
FOxqe43EU/soLxJsM8vfGyVMgrp8ADrbrg+52MjkeyHyah9lAZ07Poyjr36HpWr6
Tnl4OlZiU+2HqM9qbwRQV8XATtSLkmVbkObaxAVp3I53QGJNyB9zxJZLcq5UnRC/
UWMViGBVdAxZkrmONQ7LpPqSxolvCoGhwnIIgSy7FvPivvnGQqWB9BJDFQBqglfA
hOIZiHyp8e4L+qWyhZLVlk8T8oAptcJUDRKgWZPbZrCmPElhJaQS5CGmCLjzMh1D
XJmbMQx11p+BdSGmubBVYgO8ZL4ni5dWFVEIvpSAtynyWMndw/DXVluM9+EAxngw
1FHUnhXREznU4jH9ohecwPlskpW6dmiReextMkJUnrXvpQ3nYFXB7nyIWtHwOM6k
fLD5Pt3FWxczLGfNPhOTBJbH20iTjhoK0QfowKUHiXeZniYxgE3dJbWTLcrID6V9
4s+Fj+Tb+5XxFBFnEWdHh2DMoA3CQva1FOCMl+92wLaMxasGjnZEtg728+Z14adY
a0x/s7U1MbkKKEbF1yMykdNqVMX8ab9dsrUFzlJHq01LZF43G8mb31n2JNT9uC93
2JGn8zutQvhtpwNyZo4Crt5zrVSqgf9zrt41zC5hnvcLUt2kp1gSWev9gnfGb3VU
epwqUMc71ZtbA6Wl2WrRu5xZhecxTz8HdJQUZ0MWntG9f22nA1RtNJPKaJYsifKn
g5GYzODfo4bi1VVEyjDnplg9Lyy2JEpJkEJvxowRX4t3Mnq3xUo4Didl/+ghHlvU
iYy+ziDWssPtX56w9UvP4Or06LA5noGY1kCi8Kierf3mRV1QMWtUFeUo5oRlenuQ
F+wwPCgRlGy1JqqiR6fg5P3Km4dDzFSCRAmTsDGbu/DHkEhEgF8JlHqnzs++2qHp
iLM1ZE7SumBNlCGy87j5NYLfHnZR/HcMqt1n2dN9CqRjsUhr3ipYme78gb8vb07y
dCS4BQkHxV/1Y39txrcNsaW2+AxpAniWFv0hp7Vd5BlA4c+0qjlla3dUZW5YQkxv
8RTLVOn1n+BsvpiN2TygVo1iCJ3gfKsO2+2LV603qN0TeIOrxmFEK9iQD5ds837+
6/hu8zESTH0Ck6twndXghmLCkDenjgkmCqZ2rQ900CKKlrgYRG9yTjrUt98o+oq8
PuEPN6qlzry3F8/qu08ouyXAy1Q9eGOO6mbF5usHQOW2jpu5SyCwcXANKsrVNMSC
YX+iSeU6c/VL5PTh0rGfda4GZOEoG8S4vfDOb+7E5q1uBATL/pBvDIifYQ2+I+xl
Kc150Df6vKnrkWoPEd77h3u5BRHQkp1yc3L2hap8OT6UVGxQDrD1qI0pqPfAc8xF
ksWYzZaBhHOGtm5fypSIhx9Hg6fxDPBlB7+5fbtbXjyOS+rDWzIsrnaSUeY43N+I
BPEe2Ss0jvznDEVmTvxTIFBxzp13/D87RyyaG3q6vB59ZMq47970+sx0OcZTpTG8
w5TNnDmg4WYRqE28C334bG4L0zCtnL3S3mAnzqIoQWLdBCtK1Gxj17lTvtgdqMgr
rZh20qWKVdPSVO1TKjvlLruPgl061MtSTufpYcVZRReOcRCVM7mrEnoYV5mtOGnn
cCy8nOau+E3jIDFATmLE2LqJ052nHubr9wBD6khFbOR8YN9Uoo73zCnoUbJfkZ5e
2ED+O9KRNHu5kP05cRSumA9mQ3zdJshlh/YfRf6eppgKaqSOfsY1XARkk6V87idj
54dILZFnll+sc/9k4Rmi4CjNl5ukFV1zYHZwR2yNt1WowyflbIrP09qy5+Op5zSW
//HvIfSVhXw8l+sJ2aArhfH4g/A5D7Xu3eHucenGf6MapRK7mifVXm4j18u7/2u3
pjY1F+ygfzgMiAShHXOlk/afSUPWenlPJjr7xksfIoRQovRxSfUlyF+4v5HHVZnF
1DTovkjMpYiubLjdVRM+1nFNhXjJSyrQejXNwBvJ9bM9+z+nTMhRGr8fPeYDh67B
f1Xl5x3Ilbi0aoYg71FhtuXdlk/FnfuZ4N+7gFZODXWSct85r3NNBHgZIXbu7O1i
WTSxYV3K2MJojURm1+99a6fZGqVhHLJobnF5dj8Fj/oFNg8g6tpyjcpKUMnhuLJC
P0O3QOKh+NIjhebO40qnPhXT3y3Zp0muGBqhsXQa31sa9iAxffXrlYgXcjMQeKeA
ebTTPbSUUuNuBRIpneNBtzjz02FACsMBvzuFiv45sXN3+hutVOzlgZGLLVDBzAit
Qx0dnr0iI5Dp9nA/mrNWmzNB4X0JolnQUZhkblJxFT0UOjufZgJOtWqmpOfkKxFO
VClIUhuAYFCPHrMk45kCYvcImLxQ90X6h3qjQcv912Y3MpiQK9RSS5/4EboA1INE
TFdVTUEPIam6U3t6r5AZDAXNj6PBI2PJd7j2JnpHHe0ulTFBKSG46pGPXXtUd9NK
0OEuX6ygeSY7uJ8AK0flvo52KzceAvJRNBGeHUCTYODj9aJ+TyYQLlywigIyFptZ
AJ9cskBE4++NDqLuxBPcL987DP6hS4d3sh+oqoyHvbIbk0NFWOnLa3OJsz0z5SeG
bz8RssdkRcmDy98QAew0R4dyusRIt+KEGQBE1LvXDtGC0IIN91k1wiP+Zkz44nDW
ow+8xtWv1OK1qcyJ46H6QNqYOYLmOp/sSyf2/za24JboEsAXYmLRAySuIG4HRAJg
iTcbMfenn8hs0DRFdQ0ivWPx3zZJiD6wyvbLsZJ8Ri5qbQKF1KpwtUeDd7DBAKzy
11+2jZMLgZ++FgI7p4+YtiN6LdxxoT6dtLEsuWXEQdFDl5UKugwa/09MuejYXudG
rntD+MrjfIt7t/Pgy0Jz7oEfCbind/7o+Vzkep1BI2/dgrd3AErz0PgiLL2rGHCI
PvBlDa/Rp9pM/gXM4BnYY2Ope7gA9nFpoknlybACY8vs7ETNxEX0MgmYDbzjWZvZ
RofZpGpzC+9WYxLNkrMODEfHjo5y8KN2X2DDYrI0X7u95Gk8y7GM+/poEqYFkixj
MaCT15EcAm7w0zGUIRiQ9g+yWsVX/VDHqv6+PlYGpu2LdsyIGhUnxyRoTFq2gfx9
k5kqMWK7H1cUaktPgeOiZAgv4wdrvaxgZltjUZhkk9xQ4ceQacB5MNfa9A7hn1Vo
VtMeE8Cvv2SSLw2PfOGwHWj/KfaV8kwGJPsObc3BajmYYbDZw3dihDfP2qj7JJHX
KE1WC+vIRol3xfXbMHta2oO7cXylUO/AaOxcmb7Pk8EYlsIA1HigLxIu38fOGXSM
YQPonrR/5gokUkYPYvQbV1lMW7fM3N+IFHDkOJicWdSpp9gEnoWhwiEzf3bcroUa
iHI6VZMNRdrhSAKgAyvQrO8Pim9YlxL9/igy38jqWYuz3PjRhpYAgC6S2Frdt60x
QlTsf6BY0DpIYmXEsQz5RvZNvwb64thF8suDok7Qp01lLVJInS/nOpbS0mQmhsxg
aQV45LTxr6wQCAZ0vbV71bG+zKUiOrfAiU1QggyVfmwQFI9k/zj3IupCjAYOgCr3
W1+hA0iQdW/4b/QBcJBYnWVQirhkts7f84qk8LwjEz3X273dZR763nVqU3FBC0BU
dbkVAhFaL9Nn9uQaQIv41CLyjPA+DTAfpu8tUPolY90yLwLvrMcKhI6Xc8EbGYBc
Ribde02Ivl3nLHArSNOMNpEUmQhx0qgJbiOQrY3rDZRD8r43du0VMC+Q9dfEtR/8
vakVYxd6ihySEb/KgyL91QfuNsyJ27+lmcBwDjZsetT1lieZ/1PAJ4vQ0FQqliWv
wXcENbhGA0z5dVVr+xGN8wvEuUIqS5SYVGFyKb1GWTVAA4Yjzm6BCaCRUe3osGYc
/8Md7zTlZ/Mlmfz+jrmOQlJmrrnmcisu73lKCQxjAO5SX6oJS37Z9hInLjCm7ZZM
i4UZkF6p0TU6y6ux/ha14AJ2gXywic7KBJhstAasbNbj34XLGWKa35iZO3AjFKSW
V/Vo3t350TBmcB+Ph5Gdd8SE4z1N8OdLlZcuj/eSawiY7qAGhObXQDGjP/O8Cf4h
rlTWcMM8kWadU7+fX+OJom/mWVM6KYb5N1CpvAyKPp6XCz2lCy5/zF1W/aS81BwD
Y/Xbbs4MrkymPrqN6+bBUInu/hLXvebhH4XcaPXQD5pVR3/LU9JZB4bp+5IflUSq
eZYbamDxfiZh+tQewBYzXYADItu79JsTZguOcmRhWyAsvpqGNXLi/oDo4C4PoBqh
qPMyjZkQzZPKAXV8RJ3yoPRj/MnZrXbiHwcWv5Qhgy7mUkpGsolbP1D4SkMOqwv+
8mWj8S7UB9cxZxptoDTPhiKSSkDmuGRcJaeaLHVLGCh4SmulHW2XnCvCClKRSdEz
itaX3CfL1HEVzjp9d81L8hmay9Dm1VP39uVRtS8eEOhWlhuO1BsHqGHQv21pusZK
VOJ0RvpH1Jf5YjOvQYNXpGBgAotDT2EsvQGfJuVMmsdHFvsEYXzN4BkbaIIOUN81
G8w9QbXJ8vhILEbyxHPs+jb/0Xt6Y3yTZ+nbIppiwQ8rou9J4E3a/+w2hI7S0D1Z
hIYK8iCPNq1yWaYB/iCS8AI5FVzGQaJbiFgVwFGyiHkIKqArUvvic/ejPEPA2Jld
ON4V07obDU/u0Jxh7q310H9FfyV6+5bttz7txScxs3yn/grjYmCf409E8SkqshVH
aXX83hbbFc9DnH9c5V2vC1aS44qARIWAUkcq9jaXObTwAb9nCdxWnB9rBLBod9D8
Of8OoTo7gj/FosTcJglZfQlVx/ti37IaMctMiM0acJD7eF0PKChBZTcYtfwNg89B
Rzl4B2NzZtu0gr/z3/2iYLnX4bV57SM3otoLYsT/+3tp7WZvRE9evqbtxsJP7qT9
O/+oxlKm6gS6jh+dFWj87J0XVnnkUs5uvI2FAxk8VAWlZhzdcsuzkElPEI21YX83
TSG+zcBzaVrQ7bheVnI25SMXY2UdXcfYRK7zCDXtfjg6qIX/MBU+H2XewRqJIqQA
D299PxMUzwKJ8YnguPjsoCusEf9y8RwIchRUGMW/kO1UvFz6F3qoXmW2rHRgRVwU
p73i7CTKNJk6WTCU5UAukZTSnOrvSwtXifpKQpZc5Adeeg7L5Y0WGo2GZvbSmTuK
RMWGX5pr3KBn5a+RuZbyb3TFpL9z5swqiYqgGzZYt1Dx10+96jUjR3TN4E98Of5V
8vKpIcWTkKMajAvsVVBQuLqbrAdTKkX2Jlap95VCgS7kbLycpcwwstPIQByzgSTF
Zn5tPtd2xB31cRsJIi8PsBcxLQbD+pSCaguF966m97WRQa/QjuF5i8mZPOmMt++p
+qOxcPib7PgPetiLlzB+hBUI7ZavRmL0kJOJHit+9W0/oc/bDeqUszY8nQ12lKD+
oOmDqqScCRteSClOLIOEH2fFCaKbKzNlakC/nQyiYhJn2rFr/GfGR2DJkYcXPHJ+
tkJlUBGjP53blJN20yozKdpcYgKsTq3l9aqRC6IactzP2eGdcNAthe9h35HTFL1v
HR80ah8mbCgE6v1xG8XnJovLm00EWEknMHGRST2PSJSPLnmQlwA3uiuGcR5lxNIE
Gf5UcAQEV7eyx/sBu9zrf680A1xu7GyWoTHWQT57//cDGMkTqNnyIhhCzQD59oNC
CgJTnGnazfkO6LOIbFgrR5vYvcBfQ7JZnBsGid/kV2dzT9gqoSXPP2PlAHQoRElA
ieuVErWRYBsrxZZL0tnTm/NW4w9RTuGEjxbT0IMZBfTkOv4Mj/YbEb37SvXwbhWr
d3mO6+43Nmsw99XHRxfZQLuJM0rWaCTTs6FDHRNLn0P2A3udsl2EQPLA3Ni9cW+X
ewB1qUViCOsFCQP19E2r3Ktee8uBMqI2lTK5IkHQu4ZnNQHCnLx2XfvnKnUxXoZk
aQbrVs3ihnAKqNVas8Hmp1MbnDzwIXATGevJBaBrQHH0ZyzwVO0iErwDtcFXJO2/
ylX/TUWg/8HEdGdsOy9w6oMdC4ovFfojvsqDnZcCDB98CzxQBvORrKfmD3W7wrJD
ubrUNw55nAfITSZfgIPcHx/7W7Bx6WlVKnoc3kCXyd7sMH78U0Dnqh6N3WwXE0EL
VO0CRsNjncsKY8BkuP6NNia+3UA2Aov0ayQuLjPCHFUMVMQ1NwCyt673zXclXBcX
F2FWwkbAtae0nXGcoC6pc9zbK2zLlEEDiOpujpAnadqDXERgY6c/DnBc8r1hgxkT
oQ7u5bZ9HGeiQ0RH5p3uaoZ8le9f/nMYpa0SrMDJAbxMuwHLsJwnOwmAVXIz4rkT
1s1n99NjyXs/Ji/xewYZlbss/QWDu0+GMFi5SjdaCEcdPxh4o1uvdXkVTg2ZyjAH
+BAJcEba2D/jKJ8TXdQS3Y4/vHbsMK430HUu54aBqD20CDeSLNX2ZTqnqTrkQeMl
p2jS73dSCTIZlMJE3edy8F8XM+63CpzL50hsahsLyn2OeB0j4dVRqufbwO1XIKgM
NOoaRsWZyYBvY1da7jP1paSh010YMMb+iQY0MoZpEc+PA+BkBh/Iu11J4IKx5U+U
fhYmO1OWD5obk8x4E4BJ78dr3tgrTsDrNS4sNdTLjTIg8hZbD1p3o1G2D7ezlo7G
T/9lI67W192fKcfQ35RFxOZQyO9j9/SMjBf1nw9hpyLxKa+QNa/FrKnHeRoVbBek
ovZT3qM5k+6fzZScjhC1lCZZr1mTXmSX+VJFWiXjFyf/5oFuHTSkGP2ZpFqbW4X2
16dlLo+cOZPXfcX50xs6g1y/Igcxhh68XdMa+0wppFB8+w1QZHp0KKv4uCvGvBL3
Qos1HSM8ioC8b/CMJ4d98qUgZbBCOfD+K/ZZIKoiIYTi3jRoyfA0P7Kov6xt/m9v
B+oBMK7vt1nSYCDeSsKHeOI8+DRuMfG+sEFO4czw5VpgaGT5mi1M5M7ITquvHTQg
SzxHFnDU/XljoDjB1sb06EzAuz6ogZiA88+Vl6wWKvRg8jn/9Mt32mXj6dWwivf1
jnhLGpzRJlzWRBcISfRX3ORRXbqDcdD8TnDeYlUj8iEFha4Qn+YXds1p+rDhAiPj
MH2LF4FWJ9LHPFpWU8gHeXvjLLZCiBch/sELpNcYt74tooeke3mH76M+BtXDggrx
CN2lXk+0h99ls4hNheJqAyowHwknuaD+zNEoVrg5KxddTPFKuqUJF5VgfgavwpSY
cthADxrcV9xsQzEDlY0JiaICTFt6Tu9BmMZr+Igyd4Yvzm6GQ1/sQ2pbO8Any1zE
c/0TCNmoXK9QI0CEKmb9UwvHP/BHfRdD3eAcLG0/Mr9lq4ce9T25rUmQ5CODWdsk
xb+RxS0hYwrP1rHsy1L+rYNIaC6+fdn9Z4xKIzpiuLXMoytMuSMKjAcmvhM4sJ5u
o5UEMmhQW1msXMCgyrOq+8gcqhEQqiqXw7hO0kC1n4aT2tbcdb50W3jH0piPbnXK
nghM3/npT3krltommaIwfriRWyjap7u/surJDgUI9mCNqtvbCzyiu1YWVb/W0lat
98HbhAfVMZpYvid8WvNsyRlzLoLC21We9ayZj9PVGbTWzTFE5g3l5w5bbYIa6iIO
b3KV1hdl4D12NHp7Ust4dkR/769RzSIM+PUgbJi4Y7oLZuDxpfYFakgzrrBTxQ3C
3bMiyC6N3rvGs8SAUFz3MZ5F1OQuyKagVpJzQkLPr1heOkIpPCzmlJzIf0WvdUPH
tn0qXnImQufpJ5OBPO27bWTRi2Lf91xbduB2u2ef8/Ym9CK4Q33ljqlF7WgeBem4
aBJrMEQV2UCTiaw4OKiyM4wQ4TXP7Xz5vin9fhV2xQVSlDKl1w4+Nu75VgeNaQRc
I69wWEaayElcFl4JZVMBDrUU+ZLu2/IIO/u3GgLNPjWLpBbfxpn+Pzwns0hD2pNw
BUmiShGgKZbcuSs6maln5N2yJJ0gUZyKxau89WAwFU/mxYXzlbUfk8G6/N8aVF2R
tD4FOr/t+hYQCKdHGS5+lrtCTYeSJJphqoGsshh880ggh7JZIsI9TH2fFsaKmUwu
w2oy2n4lAUVjwmRlSCx/1C+avKgx3JWQZqiZHFRwwp4ugm/6UT1srYbeKOgzDnjn
IaJF2WvbWZAxhNtnVy0++umgpvNagsUoyXD4xy8LVgKbeSLUQg5VgUVemcMUSEg6
DDinVzpykhUhh9kIvnkLnELFnvVWWDS11ZZpmSXIle/Hq9GrD2YPyQoh+UVl/tBe
hREDuEwDc6HkJHjGhNrjIXdpAkSaPvmxWrnWbammKfeBfuuLKMDK7NHWUJPTG/ZJ
2aKUCOUJlgb9K7/BNyOI7SLBc1SnTVounwbuFZAr94LReX3RqvS06gaQduCU03It
fapYeE15HfRIS9fY5I89Yg/U0MhExiay9lWEHm675bvYQvdOtCEzo4ZosMJ51iA1
1mSdzSNqpLsjWkgeWbr1lGwONOCCTQ/YUqDGfD6rkUqfm5TxK+xs8WzWDtxOZVIC
pz5N9o821YE1N1XpNxfRT5T6GrLWSGLzIZwhr5yg5fnH39+11SqdDXaKtUTrjALk
raPL6IhBf/UNUHYJRR2UVfOdJJJvtaVLfV7YIEWW1VI+4423k47RQPyQoVEPYD47
6F51Ql+/L1ukt282wG2gMqvb5ycZG0mowDBNmb9hPkaGr9Ehsj4TfpsRQg88m0Wo
zbBDDHg9KwLaLWbkCJwJzcdn36h+yl7qoW1tRwULoAuig9tauIMqOYsVcXh1F3ni
v2z32UCB79bUceYA6Ne/aFXEIraPq/abwl7L8d90nhW44JMp6e6bl37KhN2QUm8A
M8LyVRJb/AUPvBPRZjX0dkry3ISJJy8hFYMboEviu9vHr7qHrGz/haziSG5IKkR3
2PIhmVJDKnj/bFOwrzb4ZS6aYhWrAPbWOAG7Fb1g22M9DKy6V0AGd7CFTcgb7uVC
Z+nXKHxaieGOv4kKxgJC2SWzwB9TasLBtp88TxzaZJaBKbkJeBgm9uLsk9CB8xHp
wXMJlCLUM5HwtenWqUn0zKClwO9mIwN40BeeHksa28KAIFYs67cWnkvHClA0Manw
Z2Y36EUedJCaAsxYwH4XHbKp+1WwNN4hKy6gLeRXn1tSDoGuJViN9LeBfUEkWrO4
dkI4Yy/YKLijJuOoZJnBricjLazn70MT+55RPj9z5rwSzY/ypv8h/bkyEC2fbeXQ
Ji4Xvh7/Dslrgx9F29VsK3XiyYD1m3V2JsOBLV/xig7uTXFyhLr9pHkMBXgHwKiF
QHIL7hdwvSj79VtbP+e5cx1pshaaoRIBbEPJDH3mnxcM604fzb+W/q/xGNuboLoy
Gqk29vBCpokf+/rKDqWH/AAZaJbWxea9NAkYNGdqr21Tm+8TmrMyy/9aPuZJXmWE
SJoavyDQ5K+TuSDXTBvr3Ryq6MsArI9kfLaSyxbGXb00id7sE+ZjbswOz8/l4t0p
VeRZNwLZHKlZkUILlpQPd1e6NukUiIBBSLaPTvjuP8t+t6p5ztmJPDK2TCX/aIxt
Bmqncu6Cnz0XMnXC/y1WKhpb3OTCJ/PuTZap0t+0gAALffkaHQ6wmKw/JhMWjtF6
y3x4A1gk87vosRcH/EVXaUeKV9w40o8FJDxIGZk3rTi7RdOtxUXaSxffg2EeATMo
XZZsbTlnQGAcKWo06QhFBhUjJAFojqTR7i7Sfrwm/woaZ7UTgJk+jYOiSgtfkyLc
0ndCYHgkNoG4+9EugIN4R2PeuLjBRqJ7IuhmxTMaANjrqt6KXw8xuc0DZPZ+KboZ
Fxc4uFAtOcdm1D6cxePFU+Qen804V0ud0r9GyFSoiamkXLscZweQ0/CmnmM79lrJ
GBDBBSZCDrepjT1cOJEdrURoGOuXtigoOQALkoxQc54mH/qdvSWJsNRLyXB0ytOZ
8f1L/9THBduLOCzOvnxx/4DhhSpcDVd57bCJRPPL0eEWLjnWFchE+P2AXPA2G7l4
GIf/se0iFdvCwBemeJfM6JQsqe1LpihQZBw4el4Ov6OPIU6KLphUoqMiZdDoeHtk
7opH7i4zQH/xaOs8sfFVrXe0O4DuT+VR2bKqCGTJhbkOaxoUmkLE5LRUZoiRHT5k
4H1cCO1Q9TWxHowcXlqz/O6zMoEVffyMRDBxvcAV0fpO6V8SahhkCzbbL5LqD26H
6LDmGthXw5Ryb7icClSUgFgxaQw2+gIHXwDub7cykRAodIXbdqd0PnTOOCwR6Ufx
bzdMKDHFcio84yt32UDoikQvOtgSfliUTxyD1lO7PJTl1QP0uqarD+QSpkB7FZMw
EYunaoI7yJCKd2SXELG+fuWagf2faXNyv/pVMbpPRpsLbweX9yaIQ9b1r0ut6Ob4
VIGiFd+O5rrtMxH/NdiX64actVyCmePR+w7IqoA/CWloXAlY27oO5oRDQ4QfERbr
vpGiwA3L/5T54hRaYpblLkB2WfSBE2bSDENw/qQ/cNI7cf8qgpJ5Agl2gQ9DV4hc
aoVeJ9vXHBuJf71R5beoFx1xSnvfZMGYialaxyfcRFTOF4IRakHlNipTCT71RgZF
tvJiITzubHNntZRgCVG1ykmjP0xy03fJGSEc1kTfqKMxfSdqVHhIARWW9fK8mRYs
+nV+UVfhzNkdR079h5mG0w21x7d6zmJa7d7ZYrl7uaTz+L5xYaLQXRgO/7TKrhyP
urq4C8MloP9y6x6LbzwWOR1fB0OSyo3KlAzQXyiA3OUh0sIRHD3qYJThBteCfAoR
aFRwh0fYjDdht9BVhciTzZLP3eBpUBvmbSMi1t9FWXNHjvT+pyoAhPqc4iPKGTpV
Fup6WAm11IRuBGGAUMrgBarqnaIckC8N6BVlrnroZOltz03OyHC/KUOD5IPDvREu
puYdef+LbrlNsVMiLksukUZ8N+w+zzZ2W01pCngiXuA6IaLfohXqctF3uFntmFu0
0uhZyNt25DLPRIjQkahKvJ80j3bopdAADlLJeef44G+MJWehJvTv9G9J48iT8Mm3
GC9hBMS+KPpaU69W18DlpQg/pJqtSMVKEPFV7Q34A3QHYXiSmE2aZEnoxf7t1PBr
3YkJ4UB5iUBP9t2PzhtQk6avcIS9NNzsmJJwJc4io5UhrVAMvsSMG2eVACX6vMUX
ElWkxbeRJQtgIQlppux8dRmQKTFZHC3b4EeGXegfL63cNCAHHdT9uqMx4huJGFGP
Vb6o+BKOWvaftszKOEjsA6b4+Qr3t8EOMgMsLVC3ptMek8wwDb90Zt4/j6A6/ChJ
wPIDjw1jwUP3HCN/XGp1zH0g0b0rIITmDfPgyLvjI/ymVOX32d1arFeBbbYijfeq
s/DMvoDJQH037fWJHny1Avj/QMVUujknyaFQyjik/dnq1Z2zI9s7rFw719R4IkIn
SgEav1KmF++ZTATBROiYfbSn6nFQI6TdGYacOdZmIWM8YEzfbwR6/2gUU1gV0mBd
UL6l0FtCrbcZL1INvK5C8XatKD0qS242i5H0Cog9Px0wCQGKDwBolGHqwD4ElZis
JiTOpNgVYTKCbhMyBxYgZdm7cSdpUpGMCvducuX3ercHB1FaG8dac51PDK2RImLp
mCpMk6vMORpub7R40HxE0jS+MLoIzNu8INvvyYG32YGfPqSrEImtQMLQ8HPNdp1D
pZ/ZtX9N9Gd1N9zKhg4C3brIcvjxBNCb+p2WsaLCdikf4KHUxtPdNz+EmteOuaON
nzsPo9f7dr3RO2Cm1yEofs16MYO2rs7mi4cEiViWYkJVPQZbqJ08tqePK5FaYnfh
s0ep9I2DFs09d9adgamYLG62FrR8n0Vmi9/WfHOCSwnYstUxIZbYo5ryzOqvAoY1
nR25JrVKS28am3jLDiTKMWlPqlpdHIoBt2r43KLdcnu0KVmRNw1TiMnKH7n3hEKU
d8hdKhlnqwEqmxl6ykVBW9xsE67s1WVGBUrSj0BW8dGzuvqp1hvd+RwBa1r0HU9B
i3fAdTxSO5N2BpqmdoCI+EXeVQ+T1JK7Mv6PfAB+CcOFlQ5Xl0oXpu3hKBhNeI3H
Hsj4vNTL336Y0MtGied1fo73fHBE18FZh/wmoIaofhZpPgdcMPKV9lIDmkfck2Yz
j0BD8KhHXzt5P78/NnjM8R98DGn3Fi9sAZMtVj8zqLfVcJr042Yqh2dEfti57SWV
imkCmKxNEevVJyPhOsrCCh1LmBwUYkh6UpVGoLbkTLCAKPdysvOPmmn39TyNMVSL
PPTs+ELPMEr7qjDEKHVzrWtQOBNTCkhcTn9eMiEPf8AXLWFyBpG/sKkCdftCQTwv
zgYQZeVpe+hHpUcdu0syFHHTeAsv6XllBT8t60BvIiPYvBs4MXW0/j3SaVDVRVax
VUSjchHTgCFKi2ZkNPOcmnYIzNArgH4D0LWNdSoUZVnrIUZ+SE7GR/cOQqCsC17p
xURHjdnhEUrKZ0zKCcMagyu9RIKA/DcH6oW6NhYIPSAwYGN4vzAVKA7HMfkCINlq
XWSSNk381epBtrooVYmQNu3kBNdyXPqTJwz/TudSrRZs7w8c1/34ZIm9E4yFuyVB
N/rk3KqidIbqScyioEFqO2NADW4rlMr25OllX2nnp04b/oXUY7PiG/fe+ZFeBt5R
c4327Dl2WEBju8BbBwKlrVxSEYcbOoWw0mWX6ajuSBnHGKpO3HypgYf0LsVIwC+f
NahH8gok2QjlGcnyYuOPBG7wjS9wFyrLKFfHfpIT+n3/O21IxqgLmXONlzEOuVK9
OLcIRR6+Lmq+l5E/5+B+u03EeQjfBRv39TtFL/qWXzqMqM/MI+ycOWkH/L+oa9qS
rrw5xNh8EPLvDw+lF8eFdnAcDVtm4z2X0sxnEkY7mt1fZQvACUQRTtT0SuiuY7T+
NKCueR03g3286U7MyWLZbtKJE6rXPajz/xMyjlM0uhKrxhYFjQeQnvE5v0XBSMsB
YBMExYN7Fc9ezRTNgeOGPh9JHJOzSJjXTEoMyXWCMXI/UTFT22YErort22TPnavP
v6+TnicoI66ewWO6AzznjVdLQmWgY4OTdCVFyfBy0WrlHtJ6aFMclRIaY9mztvDA
NYtQmSdJmevpnBqqxaUz/N52d+QVaq8RSRtMK9e7fvR7LMREAyO8BzqE5mD6Otv1
M2WomcJuT+7HNgy4YyevIRs26eZOhrgOH7VB7G6Gab0e2AFRxwfRWxFYtXNFYZna
M8mP0MISewMI+HWKJxLQi8xAuksgzyweITH+H/c1p4715qqTezZswW/yQnAcNCfq
FMy11e4rYxSAQfHT060a2yU3vPnLxJ+PwGQr+2iCmq9H2kYUy79h5yJbrDVFyRBr
18QOk26yE1MN9AueWsXzTf52ih00BgtYMSkrExBQnuDpOGfo8HAVn1qPyL2QMUJe
0J6YPdRMUqpuSv6svA27fl03G38yfHmGmZ3boLCXf4WzZBZHS4woOTPehPiwYVmA
R1d4WvXqX2cTal9JJb07Ynd9Q1DSZT3dnAZhXTA1i1HaijvOOGJZaW4gJNWXdPs2
a3lzf19ZeRkKwrNzZbLaRbVDkUVj5sMn9yU8CqagxBE10U6klWxiKZHw46NvMFAL
xAfjUEGOOFc8AIE8KBMFly2yLU7II6yJ0WiAdFBN8y9ewuu/Qn29SqlMYhwJQ8JO
4mD95n6RPvXMUOFvD27WfjyHiGbtDw7PdwK6KOXJ/IxrLomYjYWcQBNAX0xqZK8r
HELC38JrBPSvxqGUC0WCtxIA7/5eNSCuq4rJKMvfb5+UCFzO2OAlfQeSTrTg7eJ5
+YIZ5qiOWumRvJTEYNWwBxMPRxMJ29cdgSF2Z2qfoHxMT+QwwPzPkBndd8GGgfH3
EBNxV4Z0R57jU30+UsvYIM3QBXI3wb05MlwtbWHD4QBQhGc91EJ/5At3zaaCGbWf
4xF+uWLmA5tLtJCig1DZVMQ1LjAc9DoB83VjLsA4xWs7NXZTKEscByW6xhMKzoSm
0rUnjUv5fiUuMV9U+tkdhQrY4XeB4doFoPQhYcBzR70oB/LLgFDG5po/fnvrN1SM
pAoEocyGUMFn6AXkoIPA3/f83d6sUVGHvKO4A7vlL0lVKyKPJfiv/WKKHAzT+/Uu
TrbYKx2NnPQdKqt6G3UETYhpfSDBchZHxyDs7uR25Zaq2RgUdzeuY+W8CVwEQfTB
i6NHL1RaFtMPLG5Q5HrkEKb5WP5QAg+j8REqn5/BtNcKnO4DYleLcqoJmm9pLj1x
UO+EFqBW6rCT4nrPer7K6M2F7xJSERqZy4zWMeIiqXO1B94OWIDbZlLDCaJMiOP8
AfP0mzSnfPGs/zO7OYHlqyGxZtFuE7vUhZLYZ5EXCMPxRl/qZYXc6D5/ckEqIeDB
tlj8rU3d7b/zyXh27EtSw/LL+Xc9+i3y2zMo4sXSt1if3LeIhtSYjCXFjyHQqYDO
oqFvIpDm0Kd0Qr6ZQQ5UVGwUZSSmTq9++sHpaRy6XeRnH/kHbu3JuQBgs2wpqjrG
M+nMBD7EZYj+rzxlGc9J1RNHI/tcO3zKiGmXj0lroc+UaRMEXPAQP1wd2/5Y8K0l
lxuhG24yzF45tcWEr2QKp6+eJKnefmXLe7fR7nx2KqvxR4CxnzNChHitfSzLnVrk
c1zptXuC8vWAHzgAZo/6Wj0i3u+JbKvy+7T0ePbBPpBx2pCudUNeJOVVzf6Yjm3F
RlesGKcH/lqpSBPVM1YUmGFXCcYus4gfJi/ofkrhMA2mqiRJUFEUf1PWYtBiv1R6
AS3ftzl7IKxJuER1u/u1JiwNty8huzzl+x3xBfMARgPR1UEKNIbdVaBDtjMOn8Ik
zemgppBhoCUtqFeCLFE04AwZ4Spb5fqwWERr1OpjP6ump076ivSJUZFgMnfsqytj
KUAqB1MCRrLhCTaHgXyaXxImppJrFV98lXK7TOxkuRtRXENT92P8ssD5yYIfPY+R
+ChCv9IC5E4olnBH1vMmpheDE4uiBs7XrT2wvCfaIglOHeRJG8+UVv7GIMI93sWm
ER2A2YTMcSiDxBjXe94LPs+ZfEEOHsfBWExGKI78/zw3adszuG3My3228BWhIKUv
9+IVSu+x365okIDL/4FEFVduIHChG7w5DyfJ2ZgctkT59lTZExk0RTX8WxJDUIxs
M2+K4jot3nNP/OCYrGCv0gOl2m7YzPyO7jOBFlyRYqRwdvJJbMbDps0AwOJ5vetD
mvQXR4AvC1wwXHV0Muq6/OfNvVmDorYJHYTrGzT7iLj269jTvUvAmGwXrK4FOydR
+1NLY9j2B2gN3qSMJc8z5d4sqLX8q/Dwh8J990f7hgp/k1VpKcWf735KbKQxtKL9
RxbNIViCoYMyUOtbNYMb2H/AxO/k+ect7IYZUJDLC+q49Q68zGFejM+SuyVP1PFW
bs145Ezc97yBV3hYes15h11cSKMuTENatRIw0X8H78nhyClrFEVWKY+K4KrIrUCP
FgCfVUdsbWhgnhuA7+V06Q9MElZOjKgKqi7scPpCcqs+W7gKkCj+H7Ac7BsmBVNe
KQxDLl0+s2FVc0BTco1ZAajD2eJyouWZiY3Olei7H1P/7DTmnjGji4MWvqcJubDv
Ff0IIBgyqYM8HL7zNh9cJRgOZDfFY/V8D4vxgcYMNYkv9mejELX1ZrZutlP0LIG3
iVDEGIWf8roh0LvlmxnoCcvwPNyR0K05kpq/gor2BvB4TwvR2bmutHmft5ncGA+R
tumNJpeoih0h3FbTZ9F3b/OMkinJnAQSXwcnEsDkfzwJU5CtshuzGzO4UVtCyRIm
Kjj31sulaxaECO09UQHjIYjz8poZzqc8hLUQhhzhm5Y0wpMm32EPCAenIOL57aYQ
yhL3WCcsUFMm2deevw0JGjAM4wo2Lb+QPoOM/oWXj2TlpLKMjXSeHvAl27gM163B
cSvOdUM1mUAo75wpM8++hNxMf7eMMeWhrcKIJXB7cTKgnrFoCjLWzXLQDQMfDkDr
IYMdxoCp4qWkdgcc5YYenbLUGdBWAy80Y4NCOpIGAJCXpuNhUfwyFPNZEiFHUCtv
5ypg/KcIS8q1gFfR7CXS8YR4aVTKmtONYvwcMV6QT48+a7GdDYqwu0lUW8DTIpU/
ehH3yNuW97OVYt2C8NW5r0O+TeyeBW3l9akcLiZfDzn+YeW/ZvgctYvw0iU/nIrh
7xq+1FzvtvRNCHSUwNrDi2BrjGQ5cEXpVw3c3DiOT+N097ESbxa9qjGKJIjZzqve
yOUSBgSdc8wUwt+ylsoVWF/aRKU2A0ioi+e0PtNhHZ5wuFfBZW3lElRqp2L7177K
TxJvDGOE9tCCl8xe8nwf/hIW7L8e47sdRUu/VmCQRMwu+Zkz21xMhDzG41qksou/
VjWgcSRZ+Qwf2h0fJWCgQak1j7HtIIkocdu60Q1dcJbhdw4cjI82N7OKzmgkPE1b
aBJhfVz84lUPY7bik7CwO4EGTCizYmPqZe3wiAtal5nSBZlsU3p2jJWlJy5SOiEi
PNRPrmo1G1HtDid04UUEahceSDXAo1odItgeezc7D+aHkG1Im67OjoC4IiGw0hTt
U6GjMb1chsMXTJvz/dYAHw3TiS7y9QNfDSIWon1P+fOyNiWtiTmSalJsnYIO3W8W
IUt6CsYF2obZf/qMTEbEq2bJH5w/xdwoP8SlBVtSX2FQeEm52qjLGqNr5KNvPnAX
kUydHbrFm9pbYU5UOV9Pu3xdqzb3nREeaTA7Zperqjxsl6VEXxYiG52TKBPgIC9r
/eRGxKzxSG0D25V656+rGjN/olt3t89fiM1619kUdZ/MjBbimcDtuKhrA3mCfFBn
lyHfpZYdaNWTrDjRJuBLO5BGKNmt3Rswr+Q2+619B4scVgvyhMyxJfbC12oOKoOB
nQ69Z//9UhA1Q3A+jULhykiuqLXLnDRp1E7kaSUqWFJi7Xv31PE4bND3+RZiLITm
bQ+IqnyA5na6NckLOhdnblNOXPxAy7VHROHqNn9sggX/fvBD+LAqlrM+617iT5Lh
0qQsBdw7IyryI/ea3V7LeQ7UD9pSWqASXx8Rsy32B4ukajr4kV58a1U5nh8FbBjA
tBTNdXx0cithr2S5p4xTuMgfKmXP0XAbw64hAkbhk7u0DAumRulNlm0gbOJJZOk6
ufdZhWh6yZNyG2tso5tbg3IogEw9pYMUQSwIPS3TvzeYiqkifKiG6/hKLP+KKXT7
rIjIbNQH3aMhZbl6FZ5Z6DtndB2f87SDmQ/aXMgzeq3R1UYB5hdVd175z3+lXYJY
Smu+YuZzDJ3GVkgB1/QZJUqzzPjXeqOWvSWxNH9iRRyCgUo4qxVXstvecW0n0+py
9kF2WU5Kuf/dslWVFClSYJuTX+sWZ2bYBb4t1nBTTXSwYbs7vNvSf8/ty+nb+5pW
kF9P/x7ezZzuBYpY3KZZgU54q0geUoLahS+UV7nFJmUQDQagdn4ca+aHBFyXVIha
DwZkFtFgRawH6qBUD+D3P9rRlp3kAmeAOvZI3HIRjjdwSXFu8hock/v053lf24jW
KXc6RWMjbepMbwpF2cT0SGnaLFNn0lSXy4WLUVCqTwmvdrl9cc21gA1AnO6IZOV0
YRYLTybn9mNbpGEhAlEsq192BuYxphrurSwdgpLjcItBpqwVX9n0v5aQzCnwBl1V
DpE2frXmoWO6u1G5DWc3mQe64+e1sfKBWNmcHpTUC9dD4DcKL8G5iQnBX6TMgOKL
jPb+WDlORvJZmopKENDdcApXZleo9AdD788kFt5xBM/j764Gl2MnebiZ48i1df2K
jBlk6YQfD5nUDi4a6jQjMJxfEuiKfic5782ZsPxJ/IibZTX8hGYBr/zzCBlhfUlV
FQxzDvOSUGHEVkH2LQBS++tpOEhnPQgB2+cSrw3xB52bvtgAh5AaOHwM4pf10822
Lf7N2h/ziR9FREB+WI+RwWjTK4r80PD8Z+bYNiXjxnpCymC6IxDzVMv7nZq4e2p0
rPrM3jLMaxb8uPkejHsmNOdrJpFYwRn9QO8edzQOrJqNHSWXQfhQiV50RyhBHzyj
YwCCUQHPcPsbAraC+0DUzKEITv3BBrBASeAqp8UfZ8qTHt3xGVJ40qI3lPq4TE0c
OgeuLQ2lXHy1P+5JY+gLrnhH6A8bIqiaJXnrV2P7VPYltxajPM1pOpmw9zsAqY4B
9F+BE2jy63vsMjSYabuwjmjPs64hL+eUCzGn1TiBjYV+NXOFJzsKDYz7iX3vlhZz
Cn7OEShWwBmsvXhKapft9/87vC4LpeN6tizId5zKb204gCQ7sUQmpaanXi0Dt2nB
lVklOnWjmq01YIisjOhiExEAQIslEMVxsPDYGCWnXeDycFJBNTFBz3pY2uG5VhcA
tDhHCveby7bCV4K+gicindziqkxKl/nI/UJAgVRKx5fbnVnkNpolsyKpwVM3WlDc
IEcR40xSemQB3RBNDl+9gBj4IT0EXnW+tDG6JJ/OC+Fsks6Wj6IKX+Vm4HZ4UOsr
9XBjGumyvVpAezCdh9GI+nzuTk2vNZTSlA30GMss8RQhfU7ezE9p8frVsb9EaWgW
WP6PMVN8xXrXpGExZfwhMbAt5HEETC65grUyF7bsAVAaso69Mu9wBygcvy+jtN6U
dFHzbdleKqxONOmAtSWzvXsgsnSAq9N3KDOmY7UiDUEmoPJwWF4rGGy14+w6qB7r
bj+2QDJSSB2W927Y3AZSn+cRKR7F2uDNCDi1ECh+BmDAQAl4gfCcb4kXvDGtfMe2
ZZf9p+9/37y2XWsXvxg3vgpcxefwfv83KrJjmTX0/YwPjOtjUzsdLiRnZCy92Hf6
OiJ2pjoQbzMprL0g1FQT93zwvakVXgz/gzBy2RNwuzDQwGf4KrqjCC4ZqdJXmGaE
PqNQc8ODL+xSYC2n6ZrUIO+CP+lxzbnKZoW6au1BiIfXPVWLJ6Qiutf2R3gWzm5F
VS7CWO/oKCkGAOD6QyWjzEAQAv+dqWIVMOWUuacgu40zo6TXDppzeDPTEjdSF55c
XzegIFDYkLPJwY3I27BOEtx1s8dRJCI12xd7Gwb1LiqxAlVvsDWrLni/fAfofvFv
msnTTmxM48kvfChh/cCN8lj+hq75alVkzD+Gtn9r+qFE5meSWCs7YlORERH3V1pr
V/zGH2j6tx58sZZKos6NTDEp0kbT+BbnJcCJ5aCEYaq2ibRgoUkdd1uKN5LeCVLb
kLrvfBtCW6pYWFA5uVtEzSrFwWrlZE5qo+BkIUDF8bhTxyipuWg+FLONlj0poM5N
n/eADAoTKdCBIGI2YzqfDSbP6+BphosHXMY2X7nL9VXOjIMHxJGnD/k3x1GoocNW
igdQVODgLrP38NWGX2TxWseV6pqr63mhfRdS/Qw1y1/7Nm6+P8i28WI7cRdeS8jt
1uoWSNgchHb8Oba66GWwZ6IrZJ02SyKv+jGbVoTq2Lmni8lqIfC9qkueaVlXCC1o
wTeBN0Ot8d1dQcFkPbtmMysuSFlyQYDPyPQinZRIAHTmNZ79nTrMANufN5ca6xBt
l7bRgkCl1cHt3BtlfMdKscq2B3aSThOpcrXKitmLDCvZQL/u+hSE6GaUsJ9EZzRp
+m6dGOyos2c5npA1CzE/Bog6Ts0YFZmXmFtxXfLU7FSYR36d97bWuvc7mXfIZJlo
W4YPlPpVkH5COrJSMLUy/HEl2iOLscbCA76QHCVtID6pqfUwW8Z4RX9LL46k3h99
X8nOOgy7CDxzjZT/IUUdTZKRuOqG4a3Xe5SbUJGc9b0GAfYopsIwQBNoHO0aZ95o
OVOmlBnaTQ0NoPRrP4ku7uf7ARbE4nVWkgFfZrplApvxcIGSjpw/AFURhUKxCNuh
mR7ihO2/Q0oyDVPBh88bC0F3RV+vZx5FZP7ZKvlK0TCoVvw/QGlS9VQwEZ7IEH2l
Or7/BIut92ucgLdrJw7XNT82PsydqvON3XVO4UhjEjeF48Hijxo9FsKtKq80RdJy
xWQUPqqARH477ElCkwqzEDHnHf6lUDS3jflv9Ug/BePPkXKnc77MOKKDl/v1kQy8
iXmAny1+/6QBcn6fiIbzUMUpby4S9SnaeuMEQcnhw/jsNmh3tMZjCqCvT7zp7wX2
alAAGe4ip/3TW4OS2Bq1igTqsBleMZss9/5Dk4Idq1gBSnL27OH8nJhn5gQMHi1E
8871grGgZMadlqGYKVjnI7Ooh7Igu/9KQyNjB4P8+MeXRDv9z2EQmz8WzhVFF2Xm
NSTF15GMtQ35J6ylIZTCCZ37gTQDIbtZClLQVyje7cKjKXaVy/Iu0zB3XzMtT7MY
NfINBj7ANWXgM35rWhnQJRyEMK4dwD99km8N8l1cIS6isOW/bpowjd3VhTcaHM3D
kM8tHxuRIdw2iXtHK+gyIRHfjteCasMg1Bn62vRgCWlOCP/EHqR+a6D+Qq5lyYFQ
7BhE4xSWVa6vktXGlPS6bu6Sj4P/qX/SVT2Vl0UeRXVrpnI7KEHRuhlWGQC8AiLw
OFUnzF9T6gs7goAp8FtXEpn6x4e7zjwReYAvpsS9a5ZLQSLWIBzMuv/EBObKSrBv
BRMwLRgKicqY3JsQPZQe5Qz6WG6CjoIMSnt4WzpFm/M8F5ukvI4xHzuh9XjlbZCT
EIoUqP7tXBw48ebU6aLXPbHUewzxsCCK0U6fXGvNzBY7nwcHz1E0T7fJL5D5aOpn
6to1kSOm4dA4Yh165cFyEhM562CX4Z9FCCSqPz6SDIol574h3puqqQt8HC6/wbI6
8RqF64fOKYVgj9aQPllR02QnpC62A6CLIZ8Xj/SiHUtfOuK2H0si/dI6FjfVLSIr
GqPXLay1oY1AA6FOqf9n2/VnKQoMxWoLndOU2AvO4djdb5/Hb8hkvPucSX+cVvvn
7SwrV19WZf8cgcafUVf4QC7wygNxjrwZIDodNLOGog+DANGNIjunUGXcS4ZBEBvw
0aCbfHSU0fvvLmR7SecS6A36eBWMYL0bJ3TZwO4XgMB5vWMd0r+uT3LXaqzHT0mf
6phnu6Y1Pv1mFCjaLOiq0He3vQWDl+lJdFCXTghPRJMAVjZfTZeHN6w3ICAM16es
42fROxiwGjHI2nrVrlxwMEHmt0DgxQJfjjj5B2MPnvHZQ0/2O6YA6SLrIkrhdExz
MnKwNPYFka2E8McBiYzuxKC34pzgQDZS093VVcCyBGuVQuOL946bqhpZ4C1J9IRF
7Tq4X8O56zPMkzSoLpnylhWzAXnZeYVkWVPV9ZGOipvrRSmr/ZGz4mM67aWjaSx+
GuuGQ0DM2RgMGh00kxdE9MN7XUs/i/ObpLOudhbPr6F88YrFnXMYUbKBoEgM/pCE
7zQCOPP7LIZVYzNQCCKjpsR0hzZMdi5TRUgjm+0xJwdLzHZICQpuf4RhfXjSMkw2
8X9zl/rLzE8xPwQXHkWYRVaFVcY4vp5+fIpXMzspDtkRpnyiScMU3xJRqpinOOl2
Im075wBuEujiFeA0enTxC/nUQ0Ft6NgjwQp6QNLrnB2ETRrkuWUTrinR8RnlfNTc
0b0qYdSyKmzGxJ19CDd62bKN9vHoSaau5vo1ACcSYxAUoQv4KNos5o9+k7RQ7t5H
kd/yHtdWrJ1yi8yWyCCmqVj2jtuxgLI1C8nY596z0UKbNucJJQh7lZ1fMOa0Zlrw
GUI+IJ/gnAnwWeJVQo+fM2Ue6w3EtwmUB1epTTnRix5QczdcxaahBIw9eaK8kplX
45UyoMrG8tFANd6dEUkgGH0ZyMbLYk6QICXDCMlpyFYLDjuFf8NsXi9GKp2Dew6w
U8ALSuG/qFGEXq98kP37R12BjQ4RbPiNxQIuLZCZvnFxRtoVLqhr6T64pwYuRw1v
2yEGbJN7WSe0FroNj3Vh2AVwH3FacqVzWv18C1EqIrUFh6kPLZuMUyEfvMY5xAZ/
nxiyeung4H3ng6TbzhVoeHo7kwF5YAlg97LbdopmWVK6kYgIz1yMf8YUItyvQo5o
pa2ml+WBHCFgv4D3E5jrHd4UXOxBUf+2BTINBHIRKhSjD2BfhEZbFdCWrHJSH0Kj
kJCAMaiULgTItc0ah1m4BqOPlwO/4lfDA7fzzLegMXUgbShUrExV5qnziH/AQcYP
fahoChbKcK/4ezGLKouM9H2GpLREXeh9uBnuKAzycuZuJNbu2xdrvVI48YEneDuf
YbMhDP+HCmOQUTEspoicTYiRsXTRJ3WcFz6mLwG3Ue0p8lDBXSyKei6oVAvbUEYN
v3BNdJa9wVUCDtjrOJx6BNfUnhNdWDRI+h26HeaODrHopZJ3nYGaTsEZL1oWAplT
eXN/++ITwy4VVtAtduT7qsx5I0+Rn/PORyrOqggQ5JjCBU4crRnWcQTvHr4Ml+i1
CCsX5E7aA+HCDmCigpZNhAyvSN1d65Z+IzwraJKjhiCofd/y2QZJ1u3QbsTlanMD
qO/QBR84g5EQXY+vcY+VyXktb2Hxd9wYID/56U7PzWrkAL2MiGxQXYN7gx2WkpJg
fl7ji5aPURHGB9Dv8E/P+CBMf13LpaqSk8grHEYBxoSk7H436/xB3WLmTC5P3BMM
xaYPEZjxHSxdrqO0Btcv0MAc3Gf1s1D29AUz8zfu0AABhTkguXBYvJWUCBrEWG4m
puzys0kYbmQCbGbBYADAwErXshZAkiwbdxxttK0L42ADspcQQP+4xhIbuqd+KQS/
iKMsWUYZwO0mu/X4lK/Gpr7RKmusYw1QCWV4esojt6FoO+eNKpRaZt4c6Cf6DbK4
qyUsNVPFtW16qTeI62zeci97lwBQNuFZE5+nP1FNmOcIH0EL6f09+VCXLliiy9nk
WW7Ts58caxLKKxHNKH8GS39aSfGst0142/wv1AfdQNlvD7sJLz7yBuExXr/6gsDU
w7h3eSzKtxMC4ScTvu2SmmFAY2F8//HP/ki95zMm7j4+H4fvazx4x55NwBIhX7A4
rYz8ONhx+GUnGJ3A8wuD/7W7am7YP+m6F+9GYuM+2xdB8fN3s0imQy47eSYW6Xbp
kgvO38k/UPJxRykK3/EVhs8AgESKznSRMMVwk8wcwb6fW8DZMKs49jGX0lc4Z9ym
Dw9feh4/pqV70gVeB6+mBFIqOPQuzJd03tqfXvTqw4gGatAeXAu+Sxj9cU141Tma
TqXbwplirOmfeJEpmOKmMKeCoWuKF88pKB6xpZ8y34mTbYtir4/2vDadkcpFPfHE
wbNBIM5kz1GOSxmzGnGms1ouqHYwXApOZvg+8KwofqHLqF2ruXLP6N8a4kVArCq+
sEvKuaM6DaYu5BIgakgS6tPC1+qIOS4n8s5TSf7qYE/6RkpXWHhqHlL11RsW77BI
fTMv+fOlnlxgi1FKYdsHKpIEQ42avYWpZjAI02GMwP1bsPgGzcYO+8ilwLDQJvuS
qRcMnYtcu7koSr2t25fxPcKc6Vi9h+3vIQ3xTPK3qOqtV51Ni0TNlNHcsblMdhas
9mpjOd65owSoDvzdTMyGoSfFRu/IHr/OP0f/8Uamy/AUAahsnDqd1ign2kNoqnfx
Cvx6LdMdpfLvULsFxU8N6DNWt0bzT12uyP6PnwAf1Jj+RQv84KfWJSKYrTxlVIuV
YZxYa8+d+ob98IYLIgoAhafrEc2wmVJNIyJVa49jRh3qn4TMGIfDRS+DQHl9SQpb
VSKJugXOIxqbFGPL2dz/WRokZHzO8PYVmR+zJ+snSn36ye+OSIFIXFIssqm1yYvo
pSZ9ZezYfxnh3dZ77eRYNq9/WTvBj6tEOOvtQIVJPeoUT8jzA9S44mvnUssDeVVk
8Wo2KOMEfRY4LWNNTRNjHlgccLXdFYHwXDD+ggBFu/rPqL+a7sY+ZGEf/6go9iFU
ZOzbXp1DlQgpWY/GqKqX9ZfWgJbjKGaJ9voJ7A6RHyySbU09vBExd/EGH4CufCr0
HWzeQVVZIeJpm390WCQmnuBcMdfYvhUigyHctXZx+HLby+frGBfu+tZKkxKtNhgc
IyGtZ4XUUMGH91EWfkE1I4U9wWbHGgLQnbMwm9TR8JY0RJu3n1D/YY+7Mkpc0q46
qOtWYiuJ47Tvj9tYP3MJTp0PSaz55DzEhLjGLUew3HUr++QTYTAUyyRrDZ3gQHDA
DQrL6chhmD0HaHGkwB6Y6xQBGLdCn9Q2goZFU10QG1WnuUainkxdrXuABbt3hRmR
OonZCcY89Sfpm2TDPGFMroHIpaWWDqHEcwZM3O0YBajulsmbnCXRQb/XH80pSZGa
KEm3Ca0kR4l2E/MgdaIlObZfdRiCd/EKI5U6sEBK7iNymBTuiKdgbeNMX/UF1WIh
IbWKLqYxwzxJx1wNQFzfUHXxx6UxRnVdtXBntxN1Ir04eYxr2t/5DH6w7sZxUdG3
quCaoRrxJlamyDBXFnPjI/6i7z56l0t7Gw3yaJlhUvlGGXInf5yIv+JoLH3H3Dm9
XWb67KUIAD7DoNdKZugRaZfWJhRNaOExvcUoPdexPl/aJDKnT6qkZO2A3AfbXHX5
XSfB0ATpueJ7XjXQELfajpO2NmXlDWz/xhMnNn6ZOy3iM3kgeRf1bkDun/5j7HxZ
4Cma3IbDyCDi8QXBpqxNoo4sAlPWec03NeaVR5e558MbGxZHecr09bRJ4KqOmRDN
BzE0XXUKvn1vqDT5DS/COijXy35qdOcqXDS/OOheO9utDWbZz7J6r7+c1AqEf8hU
Cpr6C3LJazzhGMe73DUhmqU8N3s10nXEfjT2+oOx8Zn0NoKxhAAHYY+D6AN9EINJ
NkqZ/RrI6CwEnzCPkLz9ToZjd7ASkXd9oYxcHltU12KkEMAO36gh+SKH5g5NkkoN
hhjEWgbFJ/BfwVoHijpm4HSAe9MFJeGu/xtwDNy9aV5lTcqNV1KmaObu9xkCH330
bKaM0/LouOkqnR5GBkcHSE21Uo7vahEBewBObzLMrv1yvpWFomLalHEoAiwb/3+e
naxPddYsJ1DyU8ISeXuZvsATfhBxjryVelCd5hZjd31lQQTWrRdJx74dFgTz8yM4
rERevcAL7Rf4himNJf6bCLL++VuMLqJ4uBQYk8iSlGL5zgBrvPtFLA0zRXWSahY+
gGLAYNq07nqXWWhUitXlSIsvT4PCtDZBobVa9/N6J8lRtUPfEYiOm2RlUZO0wjoK
HcaFOq26rV2ac6ScB8b/3Yw9NGizh++3IbupHkMdkcNKANwJXZmN4Jpz0+kBPk9e
wreKFFDlw2DiwnWWDaUBpMG5UqrjWDTtJ5qhqjQ1xFviCHzhPCsuiWApKMfgdTlu
1Y7k4pD9mrOrO2LuY+vevSNdaayKQPoXqK9z70vI2yDQeWKqfMxTe4JpL2d3NdxN
xx0n7W9GOoochrklgY7Znm3oGO3KMkAY0R3RsNIO6ULsfWaRThfoQka60ttsaRSg
1sp9BitEHmMHAELJPR0ASgAxLoYrqoQ3NKAsc/90Yo6DbQBBSbsUZ/agYtGG2fBh
ZCz1gLc+dvpi2xBsdLwHlEh8iT3ihbo49aYTyGO76V4Pbefc2570Tec9F8lXNhGI
j0p+EhfEeuGPd0d8InoVacKirWN0DdjBVbCfQt75ODiP26TF7a/GNCYlgMrlkTiX
lmzsqwjYY1glVztqqPUl1/YfHNgIH02NpvzBpdUIezB9OJsaoj52Yv/AhtxxSKA1
1oJaUoxbB4IuIwNAoW48odIeFxekvcbtwozbhMsoAT0g5iz/iXR/QVaPrdi45M3N
M5LL02UjQmETPmhSkGIkA6+N6MdgK4C39H3B1jdCMm1ndzuWnpW9km2BDsu05kcW
qS7u79a/Ec2Uv4DyfVFQWIumHQj0F73HxkSs2Vv/1t4TfztPHNJF9sZ49jCXl9XK
o47E4HSaXkXK8JPrjPrFa0/kNLelv0cqD1Ernr7BiSTqnqY4cPTMpythzByWyzXc
n513+XZeWo//EA/K/++C7AkG5vpLAHTkegmK84LSWZia4BkxJ4at4X7hUJTcJ1KF
OqQOvgQroMQd5YBnf7IkebLhqyXCmJUq4r0hOco10dIdzGQSrJ5ParQYxXw4TiRZ
Bh6fgHw/xH1br51IEuH9mJZbr+20hENfRD59RRD0yP0JHoxV36l4tllfAPldNJ+f
L+9h+d7hfEUb00TVwGAx4+M7MlAmaUZxNecg5vcXViUfHhy2NXhzGUzTVr8nmNjC
V5o9L5i/nVZU4tf4+zAmBCQ85vHMOFVcqZDOJDos7QZo7NPWH/dC8cpYcbaT2Eou
It3bZVC8qGDQsN76iuy5f4zl+g9K8BJhtDDZm3leIVfi+0lnGxiX/jvweYewxj+K
SZMo+Mr8/hD3eRpyeZYdgGBQVpRTCY2RRauhJCkLwAEAYBr1XhHYnp+Mol/OaA84
z4eR/4CjGPlxZHA7duDR6WnRUeHJGvedQkQCEOvXisTwudqHlrOh/qqenwzoLjzm
5rhrDLObv9sgsKvVDlb5TjSstKICTkYvChB/XurWUghMLsTj8/FHNUJkIUh673Ev
MBmROJpwcPGGb767sn8cnyDReL7FdPjV1+85ZZ6hyCdCwq8NQ1qCmzo/A2gYUH+O
oGk0SBnCMHHmn2sOq+BuDDkowEFxca0x7cMQc1z23Z4kpTHJnQo2g+elLP5B4rK9
QUyO59ndwiHsFGiZqyQ1SUfLIPwh8beyjCbe/fnQj4AY4AnE/PcNoBr4VSsvG6yH
HkwdC7Sh/lplZJ8BYVCL/VPYlDzQqQNXAuhibshjd8bCtjT5KPBVE/6zyTGTORBX
P8UFxdZmeOEemz2Xdx4hJyklnHYSI2wj/dgqYbWItp4BBYRqLqbA0XfiwH7+unCL
A491VdVO+AnaE8eO/IBTgafUVm84Fo4Ic9kvjnF+5yRUbl56iOIopnctMSth1owc
7/E54N0WxNd1s36pMo50agXZr6uCEbWqTjb6Nk+3lH7cHo53l2eBfu3lA9RMjhaK
q7WKWkDDdBg1Kc+rbVgmXP8q/cByirFDYaxk8cM1UrkqzbCUwbIBU46kytpoUpCA
hEn2zxtzIei9pn4h3H1lSOddHwUDOFyWNrJaLZvnvrMao1U69IpWM4lyZw3lfni1
Lt3pf/XWB+PhktRrxiczMVUQa3Tg1wCGfAg1px9zLDBDa6lgJbt/fCEZ3jeQU12O
m5xweExwu6KKbcQy419H8wzR3GpL9qYo9h/nsKG0Shc0nGn+QKh693ypZtCj+/rm
6KFmeudJTpQVYPZqnSPXRfdwuGROu5Wf6sm94sKPC5TnJvZ04kut7UI4pUX9Aut+
zYwHYmfl5NFTipQT+ekQpVE4iI62kb9HbEPik0znsFxVEbuIg7fMQhh+CA3MWfGH
KDm7j+L8Fii6/P4+wmSs2Gg/mKVMpMzJDJF6OlpJMrhgrSmF3Lf6hPXNcg6FDzz2
ObDLqWfquXRhHTXSTcJlpzCJT4qMazB9AFjsQuX5uLSbjKSKTs7XpnDYiA4qnS1D
ppFEeBDa+QrzIZeWqUgU+PSifxEcALRZBSQh+W879MyVmnj8lCt2hh5JD1cR9r17
ROIWAj6Bl30jsHfhMr3gg5QYoY7spZerpeALV9TYu7jfdI1zsGGAEYW+41/qmb71
ZLau062XW4GwSxAapcajTnwkyPgHVhqGYTFw+ChKD+ZbawygEi6c7nL68qaM5Viv
y68dblOdHrMV2xnySKpQ366taQFlQAlZpTtes9m+gmBNGpHM1tu7uTCUx1ad9kmN
7yEg79lStELsqDT9drQk4Nk3BQ0Tk/dtQI14dy8VcuSCQK1YBtFlKiagvKFXcarc
tKIKdwUxOovQy/qOkJC3//inFj5fUvic/S5AJ0TvOBGg+Z2owrbAVLK4rlWrsFE4
zhQgsnY9bS+/M6+vPfjsrUZfeS+Pai2W21xnT0A5pXBUmgj+68bESp2eRE301nGl
FwJQNLXVvnCGW7wtDLjrvTAscBaLYcH56WvsQMj/XD2/392+L4WKa4nkGac3v3m5
gU7o/Pds/5GGiJC8iwi6jmzff27ptc/ahTtpEkjCHL/pFDYooSxGsawdy85pKHba
66PGzl1l0soZmqGIJ9vzAPX6USrcU4vHgq7o9Zwq4ZM8/B9/xji+GNY2kgH6qvkC
KeAt9zbyGK74jYTklA5LVSYQvHfqcVHhmRhApn+OxDGgAs00/wNZIqDPsiv90Sr7
zQcvkD4jxugMP0TE0rk/FIYwQE2CHDlkMTcJqaBh8yhcwft85JnLXVHKfkkuyw2s
ntpHevo0c58TwEkX2jUxfywlIpgYTpfYbUjdAixVHiTncDJhffBM/5YMg1Bt8Zda
fYe1LLJpiBcm2ulgIh5dBXoqS0U3Yct0qNmpiQOme2mrICwpDMlhjSOBqeuLT/XR
2F71+Hr2/d8B0Z8JhxxMJ+hdfwlUTFv0OszQ9uRvnhxPU12oMki51mDyV+9Tn7y+
b4IgojQl54boZ60ashzzGJ6Ndb7VMRu7MDh0M9MXNZ9hhC178FtVsoU2A4yWRrnM
w/G8tV+1mfxrSHHhXBogxkezvo49GCSoBuIqrmi4JLrzhiMNvTHx7XHGq9h9SnI5
ob8L5SMhW54HdZ4FlUQtMR3jhYkXLuQhAegUuw4ASfel9U2CdfZK5XMznIgodzZx
JdKJQkHBwbRf8jBd9uNNZZSBqHbQJFCtWTytwrGpO94dc1fzvvIA3gsjCo/5+0FH
1GdrrDxs45G+bgQnY6qpNADbjQcvZXWdCP7zu3TnrI2XahzbU2teOWeRps7QlKjs
gCd0hVX5ClRiopHC6Te8WhDzEhYwn4pvf73q3f+Vc7YA3PN5fNTFl5A2Y2TjCrWg
LZK7O/jF2Mw5re6TWb0rnbJ19MLSn+5xFMZ+ANLQiGYbCabVF1IJyskV51s+HQYe
jFiPgGUUhZl7BM7Zim2mhVlKstevFWR2MZDgygAOv9mZpDHxWUGo5mcyHLoMl/K7
FaZ3PgH+KoPBT3UmuBxxp+TKefSl/i4srLqlCDERhzJZNhVuhY9oHRtbj74beOhQ
rmgu/3/5W7/cLvDk1d4aA5QjBLbnxQsunNSyw/wAXn1/gV0B01+McnpWcrM0COmR
p9uty3YcTWUWLh5y0Akg/9R0v/iW2raBZyn3g8YhGg8sYoBHhG0eXTFGTdKlerE1
tLCrEEY/KvSXt7W6MB2dbTDIPonvL4gO0wqdghzzDYUbpW0TTWjEZsZQr8SIKERe
5QR2iZlGz/pC9Wn13dgHQh0OYNfXcX18HymZiqzAsoCBSBGbvPjHQTq4Fn4D5w6U
VcSWjJvBuUZXwg8n9vvlJDBbv8g7B5+lYlljk0i2L/remwrwYCQLqTj7lu1AyfCC
rdcWhr1FGctbHAvU6xFryjUSuO4E+1I33+0APo5ae265Pu5yxZDDSMBWZkOLy77u
pLbZG0JfwZYyIGjwIIH/aKRJvLYYXrVfEFev6pKq4MnrXc9e/3MR14lzPA2BNh/6
tKtiINuUjlOOc3pK2C/qdFRPWIBkuFKGbNeeuOjyuNz3HFcI6/FQjxZX2PljaLwM
npPm5lsp2fpNtJzMpucqLZBilP/rAbr6EIJl9QZSvvpaBh36GbrztREjpGrgBioc
Fch5ynZ+A4d/oyJbfqNsAdU1jmMHL6RGkpOZ4p3aK9sYT/O3MN12iltRwSv1RAfo
rNthfvTnztnWZxTNPKxOUUn2K5wCopdA1LygEKwsmonUKFUYVbkrqLUf56Uz7csI
4et+n9evA8oz9qYSqUsDYFVm2JUgC3r8I9ynoD8tZFiMTR2Y7+JTzQl1A95Zl0dv
7FgI//OopbLKQSXX/Z3sSFNgp55M1Htg0uDX4DUfGCxB7iJLrl4bud4sLucRGQ9G
DDXi60AP4zGYgav3ksmORV7EzKJZ0VTdu/ug83BTXAS4QzO6kfrIov8mNOB5fCSe
hLXoy0ewx87GpLvDWGnQD3MvA0NUibOqtDdwm+tw8LksXegNs3qbNfaXE2J38qqV
fgT9uOzb2wjwOr7aJfCcDuozJZVR2TcfCfEExVl40KOn4DaS2mWeqkCm2na887jy
s7yqxTxKGOSgy3IPWVHSJ1g2e5vriwM5N/qUkjmblwsS6J6ZuHrbGuWDJi1CXFv0
YMO+xSux5ogStRUGArnfDjh/RhnTbYeF8L9pf61pMI+lFC4ePIjb9C9V9vuJVhsr
kq6Q1TM7LpchNf3H45O1eweAaTCJILpkjEosXCw19gg98oEGk5M05togNd+bX0/x
Ji8UfsRdtmcSdOzOxvrzpEpMrnd5musAqDZDJxeM7x4mnUunthHoh2/lkXOHvVul
qOABncLsgj+R6q63H40FxbEeZsS+u9h+D+aCKd4Rs/zbgxP+d9UULqL81ExHF5lj
IR2bb9cEW+GNHJycoHfo/zerZDz7HzsNyINzpCqpriQzCW/u5LoASntTybMyTXhA
qsPAGcVHhUwrxo2G2/0DWKEX2bMTfcDt9pGjHzbPgMDHiqLMnz6ZcP5Tc/DEevnl
S/8C/LMWz0D/RlAPyuf7Om/QNcWkRgNCAkQRJAD5NZq41SYVwGpbuCK3ZjPQZVB7
hL8mmYotVQHMZfmUhpKMg/Lr2XPvSMxGDmrXLHzZfQx0p7mcKkmhlzPWVHmjjGwB
CDJ6bazpezJYDUtaAD33D8Q+fCmAdICauGJPME3fK6hKNQe4U8m3QnzWBgITDvBe
RYP+Lrqzeoplat0dyr8IHjLkErXfoORvNJyhl0i+3FUP5bakcNlicwcNGNRcmy2q
kiFRaSY6hpV9UIXqhpLvOnbXNip1cPEoT2DtFjNfrCCuA6u1Y6BUGH9KPLSkTjMZ
7/bqUb8yBXguQIdVKNGPLDic05q6FUGdkhphlCDKZUlVLxWfxE7LExTWf1vjvSlQ
Xaid6M+6FIpaXUgp1egrouE0mQ17Wk/8JlFTkJFo+hAFpXBVwnOlHm2vB50i0SMo
suBwuqn1XQ1NS7fNlLeup1vci50sSOFSHQ9WmcndZao0QwELz/21yeUxyq0+MCNa
XKnmPTMGId/R8AOFHyvogwlf3ZzP3TfI8Yp/47bp2m2QXZj4m1OWMAWJlCSHW3Wl
/ZqxaZrOH23yoyYF6ZqSemuxtvg5iDQXPtOV2C1dSYgUA1ZD8qDx6oCCdOUjaqdV
VZKo8QcSn/L9NyxU8MsiMFTfi0/gitG3dxTUxc5YNfEDzTZfeWNiPu+I8zDeBKXk
3Kn2rPJ90isI+MarGOJCBtK/su80+4WfsRnP5M3T/XL6sFxMS25i3YSZXX63PzOR
yjf0HstmYI2VmvXkbMT85SR+6OadIcCdfEaWUsmhOfuCMRs3gxlQYs2au5lQiFTq
ZOSKK73DMVMRVgKdFqjTr7+LRjoLcEDeEdPIfncMO7FYFDVJNukaP8GPgr8Icd/8
K3cO+412DnDiAwaiPhQTlwfiGBVtXl4m1vH0hr/CoOWOwGgA865HRMvDaSLtoFiH
Pm/WXHm1Q+mWIBOOqGyww/nK84idBP2qb5GMWIbuP4Pl4U/UKKm92oGAvReidsvo
OyZV6cJCbYvyq/nKw0MCf3i7+Ci9zL+ak0U9EIYOGLo1lnS7+NoQMTaJMRVz1str
r4nVuYtRd9tK0zdMAjR2X8cyldHpKeg+zV0tgtWpHfeaUGJb+XhiXrxus974xIvh
7D+nnOs791u0bQTmq896zHkBsQ8P0+hVQM7Oy8YRpvXSmaOzCYT7UqF2r9/G1Fwh
xYOq9NpVA83eUUv9p3ReVxEJYmJkcujD3PytMhpw2VRg3yQPdb/jbF5GxnCXzsBr
YQyL6idiRl/7y/xLTxLADM9vOjDefZaiHCFXL85DenembfE3OeOqtpCWrdevAifl
63L+6ciEDG4KBhgysEil0kJuRJ9i5pu3KhaU+q1fa428CqH6sSiaE/9p2C35tGft
7fUfXRurai7BzavEX/ekM1cQSAtISK9jDSbw4Kd+gg3JF08sWLV8RB0AHxEUw+Yy
moFd2262Oq9wFB723d4HaaW4zDFVzytIISqaT0sqs6CCW71poKjQ+LV6qoMxBO9d
ZRfcDQWW9hRwC4LcQIdO98YP9e39mFozU+B3Irr1r43qpYBOkbM4RMuzr/e8g4XE
yoh11lyIqjAK+ILXv7lSoiae/upYwa50kJnKItPlxaE8kSK7RzlmKEzHsy9wWp0v
WMUOMdXm7dhViqiETpe0mYsR73OuKd6KGtzMehKPqBbEXSEFrNfVoG7fKIm7uMg5
/cQ4edGrkjXQbL4PG6ItCOP9D/zz8+6GOTKv6TIIXCq7s8rf2grdiZeA4Ufxp2aF
KSpJwOFmFd7feihbJuezpF8ElPX3Z+Yt4KPd9Z3fTVLXE1aN5W7MPQGYF4AIQYru
U4MVGVrj96prJaCjuMulsMbMOHSXmNFU4F+UeJJNNheoQQ8en7bQfmbkoAfgyAZQ
Yes9kAjqaU6Y9u1zvuHBbO3IAPQmU+VX15ls1RNYlZ+V9FKXhqzzDgroYJK/o/GK
1D5/VhVmovqxdTNaAMl0NciNvEWeSRkpvHwEv/rpIev6I2LQD/5b+0408zb4vgk3
AMJWhi9SIcGx0AN1mMepUwyJmbjC9BjbmZCUIArNBOQRga3ontVi+3ikdtffYcLh
64Q+7rFvnbR2M5q39s/eoVyZhT0kpMbDauVqCYqIf0Jq7n3xigDpOa/b9FprX7+z
sQpSSMDLElALgfr9DjHDeqaUQcnJ2mbqDOAQ65T+sYCeGdJGJL7jRcN5JTRtIPr8
REQl9LTsUVfMIO6UonXMbcl98llacwIqHj2T7Lxmh0Wl3FxlOBg14sH4YNmBFoJT
h3GgITqmJlHOvxbpIZnnT/rQTon3FpIZJE04iv5oWP7YFk7eFyNNreee20iKRabI
4HNg8KWCFjZpkKnaSEu0I+6GIn9FZzf22l/VUpDszhSuf3zjQ762A4FrWJrEqJQ8
AiPi0cm8rbvWf0NINLjJv/OhOrIygyvNrae7EUO1i0CHlSHXLwZF6qb00JZcx+ZI
G5W7HF4bOSja00Q9zL2pD6160ihpoM/1x2zgmNNBbr8pRLRz0QXNy+xCGypNFc8g
6TaOgSRzY0cp+uzQiXSdqetO1wj9a0idzmrjEB6g+BFVttj5gewXOMV89wzkcIkp
ZvnxoYTAr4py9Z5EjeEbhOPIpPDMOi1QKWOcq92uoopTFmg3TKEw5c9iypYwrCZA
KQ37m5RWm/8eExAmYIH7wyi7kG1XhId81F6dItxMCMJIMzkCOTOtscxUHY8zDJtd
xAuPT09L99Vjeb7RjCnKQR+T4S9SNVg736F9g5Q69sWggbYWCQFfuD5mXLGaeqMB
iEHFCqqDqzk9xk+8Ap9ItsTvTnRI/0weHjkVeKRp6wnw7KIqUzwM1i8sjDn6kH4t
Dz9c7775dv5NgvDQa4Poq02Bbv8dNYwXdJYnJ3cg5gGT2zuleEIl/o7POJeswgR2
WFR3lQTLNgVGuH78l2lHipBqyp/1+yNAv8XB8uaiMwf9+9MoWC81PYiSqijwQbG0
Zd43SCvmAhwldsoJLtHc+RD911DUHW1ougAAbbi+ytKVpbSyMuhNo5GlurNahf5D
/31n/sAfABgnSUaaDxlgxeQYFlmmmsrEk+js+69y/brABPsZyjPhI5JVCuwpw4Qs
fxSIBTrmDQ218HpplLaJLD3M5XXTlev/tlHyG3ZsiJx7GYCSuBN3fpKTWZkBu43m
e8M0CeiDywojE/SqdKFWo2+hEYIexVsMa2MFF+NS9h6+XMabo6cei3rotQumcRxB
7mgjD9TDQVYkDE6IN3EOQcShzPVAXMeCV6kxPJTOejmh8zRpw0MwZj810knZml4c
CW3oVkIjZYdwFTgWBYcJylMj7O3g43G+zohMF2SS/6XNtHFJkkfkx3dSuWcf06ux
WW1ZWsqkUVeLsBSWRs2qaSM+ojOTghmnaRh47llcIjtQBP50qDrGyJS2EIGrV0BK
cAbpOQCfy48wEqthuB/vKmnyjimz36GI19lnI6s38zRkT6Hkqj0kJCyD7HoJ2M1s
g02XuMxfDIpYMZfqbg3ktnPIFzxHA8J5eHVE/Vu76W5//6kB91DONpF85aML/D+m
skIT5lFFLO0TS60sgIG2zNoVzMZ5DwDGY16od20Iqgdd2CnB7QNV/rNI3yNRyGx6
ouqLy47F0IgQosZbi2REJylNffL7Or6MnPSdZe9TBC/1Zt/KkC0j40HRH6E8k8JS
9YyJUsOUPQMSeMgjn2U5mla727dEaYIu4Yy4xRPWs3lv6Q674orm93x0dzjbJyLP
xkGjI6MLGI+sxgDpcWjcBUky0eZgykferfEmfKOYQHOIF0VsHB/iVZYrs+xJyFOv
dstvTgrvFTSfdJWnUgk/kL+K2PJXPT7dqX4WmCnJ/boNOw3SfdzlSi83++szpy1/
S5HvWiEk5Iw33Wn2aTgH60H/KF1RMmUQzOC7A4EP8QDnfyFrwhBUNoczrnUAefiP
Hz6i0pyTjf3ytK+L49L4lI9PZjFh9DUZG3h6zJTjFFUXGX0Be6AvcXPc6HJdPzDe
26qqWtq+40rdaYJy1FHveE4u3OmyZQjmUCTkTriOrFOkwDUOA02lOWN2vzalv9uY
/+VWTWnsoHMX6MPk0f1XWbd0VnTlGNu0r2BDCZoX5XJMCI/sg6n4thVzJKExyGM2
DibG/jDA2jVk0FhoW0pgHD6ITm77m5m/l70poPOkYYcD5X+Ke0P2LMAKSy7ez1M6
weZOaBGTRJVqb76tqv37yUXvkztXVKV8g8n8RzSsA9/kvPaBWf70AxSxF6etukCO
WYq97dkkLS3TPXxqNOB3c4oRmuS/PsscQUd0bpwvvcEbLP5a6DmU4370tjNLIJgS
FI3KvJiuclHLrAAQRMnq/cnQo97S5c3SOm2aBAVpxiOIAMeJn5LUaUo//6oANgbE
E+gITkA2syJ8oYHktxq6hS5AqRQp1BvbYfsiXmJqCOpfGQ5xtqzS6LCYbXFNse7T
YrGFHNv9Cn/Kdy+M78F0FCgXoA4nLiq4sNJ8c52HQNMNknwA8NLkKkle3UsxVnPb
IwFmIiBhJ1KQKUZjRi0vCwe3IVk0TSW69NHj8Uit5kqx5inWjMaafdNkfmf7y+Wg
ccw8a7FeljZ4PAVOzwpZE+F8Ll358+euqX8048MhVkocTyv88uV4H4wayErBJYnf
hEXMOwZhrblVBS2S+LYRcXsczXGlbMVC4LsG7x6fPmF+CYOCTuJlw13NthpMlKE0
gd9QatOL4h0L+/3w5iYTi/DhIy+MoYbgWxpz3tKm6H0NWoa+QPkbEEysGLNNjyFw
Mv9iarVy7pskBVph4jsYVIYRKOGeTiUTOFx4WcKdC6Vpr5596rAVXX0DNXOWdLN0
Vpg4lMIzjF8I/9uBDFHX8PRqP73wDj2fQ174H6S55aCZ7xQAPizfi/2EoPStRDjd
FvsglK5giD8mbTet+DvpHMB3KaypFLGgVW5tWAMMeRRfWffstdC2+xTJoz1eXbpz
96LtU0lC14WFwTemHviAzM6l7L/RKRbXkN+jKlkpsq/qzX15QSbaUYWGDTu8FU17
zT6AWDERoVD6c0o/CY8oVUEnH9Rn0/t0IuIlDNevE9RypQBSCiDhg6H3aHKMLkhC
PtSysBNiGMHpmVoA289GzrP8dj07aX8bJHTOzr9Gmd+sXtIbJUupf6Ha2qNt44aC
Nuq2FYhyZmevRBn8rqUPWUNdVazbAfu4nq3YMDtFaUMEDo+w7IXmyhsWWRfDdFQ2
LQ/l4KKhMF0NIpLS8xwtPP9xjbPUE4gOeQdABZKIhLTCxvlFp3/7LcqIgGdm0A2c
hdpli57aKTftaX2cH50Ol6yvbyakcbLvyjN/U4WMrJBac9y8/80S1xnkmSmIKB0r
RczatX3YypcPa2Jc2y/T4+QBExnPV0s+cjChfz9K4XMCNhNjX+4v9uIUV0gmzUAx
HYafE+ANgbFg5QmuRTfwpjvJ+NPjgo1qX50H5nGRm1zvgZ5kXfjBTsCkuZzgKGN3
rYr2W3GDrNP8OJxwgMJm4ir3WOZ5dX+aA6RodDcRr/sGIeRFSWXPn1Lwryg7enXx
KlzuCgPDwn45TSR4YI5TfPq0cMacEK7GFW7DJwAODg0BJboa2tuEMklI2Sx7ffuU
YaS0ePIgD+opDnrTuuQ0Pn0m8ad0v80PXWPlLf3lMM+Wmx0w1ZIeRknUDrcAtZNO
IuX5LimAlGfNHPqv4W6Q0EsEaPUqmOKpCkUawqy+cgI7gl5jtEermYFL+PouO+Eo
/WRsNwj46VsjRbvf/FGpWMc2y2NHw08AG2YAhL2BbKrMfEY8BxAat8QWbrRSmlg4
JJhlN/6zMGPdGYQsmxj/qZ3o+km+BMnZWEBgVIJxeOjYOdR7H5WV/eYTnNb+mYmh
SzOla+cR/UdINnicae89V025aVJYLJGAVGBbILJiwg65Mus1IcUvWdacwWzIuec6
uSFVDbUCnvYAGcB5Eo9ltsyZ8FKbpNJy1zcb/YwV2U7U4mWij/nZ16GCXb1vdiri
FQpj7dl02qZ2f0IlQN/Z6pyOOFFdCr9FtsYTlE3iHGoWCaaduoH3GB3opcgTmIFo
a1vT8osCB3zoSlj3PZHkKPSbzsVwcYAv/lfbXM+KOGeXfhefE9BIsUpSveWabVWZ
tpBVRINeZwkZ+yizulEAkOEk63VLBPrxf+STrjj/cDU9g6TkcGrSU9RB4HR6Upsq
iPdxH3py/SlIkXxO8bHnWZqSw09Q5HLGjdgzO9iIe92+8sN9lYSKr298d7NRSB7a
PBMX6lr3Xtncr9qNFW1g5UoDpQ88ww1wA2MsaBKasDeJgKMMm0s7pvQdvvqwfR8m
YzmSJKn+DOovjBA3HyHpXPhEmmxH+6HeEZTzKK6v8x6rpX6E1jPAuxDVEgUT8XLo
5SU1dEgXefw2KgOs0LBxdQ30FZoJVIWlxn58MPxNwp8Xd6ItWlU+KKr/8thh/MFN
Jxj4K83uwUPqGIYVefW4sRpn4ZZjU/PlRQq6OXMXkGGStQEyKfXzknox8SWfUEcH
v7Lmv9hqeIbpJpg0zag6fx3XFnyS77zFAcoltG/wyDnrYQXMO/1WyUpcdeN7bVms
ANuuHpDc7V4rP26M2DgZxucfu0f3vSLE9Fx5BtCoqAjvyyNLkViuZYpaJFG9febP
+7ah/IkRnF2FyEEXSkfC+EQiyvrlszz52Wdl3WTA9Ak3XPbkRaIveJQi0/+sG/7p
U0rxDk0Cxm594tSDVWsSh/WyCXxSGtdGKjJCwSfdeYcJwBevzLQDR0HlDQiHU3of
Nnjpl1+3Hn25HYPHQhD4fF4yN360icEEpN8yYpR0Vmo/La2ezkANvZ1roJLksm9w
/6gca2TO9YoHfm0y1vrVmIa3VJlXWB7ntR6FWtMSnpopiygXKRlHNei3AnHnqwVS
HvREvsqZf96F3ICacu1o/NniicXnNx4Z8/JRdmnHlEfNtoij9qKNcfmC8yFYKEkR
XoAWugNOfUFsTL2xyz9Cqr9jjJSfgPug3DDX2qmbaLnTuDrElIGPXS2kMmdk4iZ/
t78WCTt2rwk3PpoIOg4dWWXmfnMYCREbv1UskgtsTBRPkkPYeWyu3Z5Lm5F0uTDl
LY3y9zM+YlzskSfBA19tWQfQIOfeFGdJ104wgyVQlRHJI9D83Vjhwg3pPohaLsyC
CUAifkaafngEaMT8RuEASkRpLFUFSye+jERwFmhGHq/G9I0okyPGNb5wuZhmegLb
OGbvOQVAdRINRRlRbONbS3UWqSVvVgmRU6s4689aoMzlzescFb0oQva1sswb1RMo
nkGFmiU5FPBg41dO5VXAFWXsBgvXzy724kezY5D7VwwZTRKJ6AyCD7rz4hidt/MU
iebXmudZBEyvyrOxWfNvfXGQ8J+s+66nOJSCuoXQLdafn+twmNZrD8a+4A3GOag1
7raTCTjeZXvazHDa8/vZ0Ya4XYIxBQPGBlqS4mzswLYwxH+MudgLbyBVNPZGGIQC
7986lmlMsaXh39HPB6a0F7x7Of6hrApnHafrUrGMlTvpUHIVCtWlinCtaZ1om/TA
UPOC0HdMHJ4OkiF9A/h1SLSOKuXPGery/V6YNjm3MbAXkU3nBNUT9huBg+EpytCK
o8WghTbj+dLQJ8gTeBn+EO5FMAvsJRoSCh22Vbm9qomAmbcAWCGmoQ4FXp9NOnyc
Pk+bUu2cH59+NBBMSCEotmTDcapRp/LXbhrWV0VWwaMAenILGVvUbdcVq+t/yR/U
9G9Ot3yEOKd+8yW+7Z9331LEpwDChhv1c+KGxYBrEPEOx54UXylwcOgLrya1TnFj
Kjmgt5zFS0+sOQDMi+VmHKDQuzAFI+UVUDCv8GNpHP+IrADsCVFlQ0+u7gKorU28
o8vXdKncasszWDe9QUUxLiiQS0hcwclbJ9fMGlPXA+VyIgDXebTXdOIVuxE0Pa5Z
IdPDvu+Q08bAPz/CufEt9Kb7+2MZ2uqvUGGfKaYrSjxxQpSNdFGjpFgHr2NdXuP3
UfdWvqve9Z80Ih/oRg0X3XVxGRRLASvoZAhstkfuIl+2jDbvX5C6X4niNxgODKo4
zTVRsr+xmQh9iz5IgAH3LdWzivQwlc7uZ802ur17oLmzAwpJINr24fjq/JUJSWP5
WVChu9TRu5EgaVhaZplSMrf7ui1EqHBdF2Nx14iyVWdRSFM1RJIoplfYvFON1oOE
PdcIcSQ1qQp0iMkOp1Vb/6a88+LaugvCqr0HxX+ktMZtinqMKE3TuYf6UoyecioM
j39ZKDQaX8lnlSK++XL1+nOHZuXyjLc3UcFWdxnlP+q296p7pZ6kzD3DikHkRMk/
4Sn7QsrFub6dQ3odEqHUg6lSusGbDDdZq/17443Ci9Ijp7AO/YT1OghZxOACB37L
fuY7ejqaTUqgiiLiZyqbEpf7C5kmdlnIn83eck1vxDFsAJF147cGlMo8a80FEEyr
/TKFUqMG1xHgM1jC7B5Swt4rxAj9QGlrDgluR5/c6PGqV1n6P7jAGu2Hi3geWOlX
LwTzyO1UtWOTEA6tYENV3sVsHmCl8S2sksgONb6BYZool14xx1m3NMARRsYRcd3d
Xia3zSkFtgNC4klCKlxRr6qgezcy1upScnkhhlvkICXpYmg0Y0C2Uwdnl/gxPoMz
NSlhRXfjdwnByeF3pwPTmUplDFgx17zT4kj4xR4ztcA9KCbfAsfrdtBQHtq+SLoS
C4gYxsfXdcAkjveJg5dZujEmdklW2qCuPjFn0zpPQAjRPzmFEOObaeOOgNLxwGsc
LOwfNRgMYgKdMlCiq5L5F5LP1r+vLaXoVkSeX3FZ8Db/9AN5MBt64BAaAVbjpd10
MsHKn0/GDsfZIWLhDe3Oq/fpSAOftOjn/66JC7M2p8frscpL/7qw2ks44ZlkGbba
GdjEyM11hCEWxqvJ9iqfHFn+ZEy6TLM1RdbVE0x6chWQFawnSsiFKt3M2uwcK3cP
Ba+3J5MLAAE7+f8gIGyTdnLB/JmSO5S/HJz/hWR/fdvWODeOO89gg2hJMRHSa0Xl
S7hI7Od+9fRjUd0AEtaZw357BHobxDEZRDA6b02t320SvhVjzxAyMGJKruwT0JdH
gWfaiSbRXq53gtWCrHDZZ3vSUMFkP/UAYIFKrsDGM+c2nkbX5NXTCdG94dPXd6nt
4bjjbrwtoEDXCkEGQUsbNgXOSttrvbZC6XTfksI2HPhXW8aqdbwZBk8X3brY/ryK
TU3k5hs4Xj7HHksIvkWUZTN//wn/ChGCvHFDNMmvepr3JIn8C3TLmzSNsgy1hEsQ
2dHEqqFLxaxVeNWfGv2H6MDHYm3kUjJhkWoryOstdaBKpqOPRIYth5b/e65bJ4Vd
aMrfHRtOVC/pSPdm8XI6sMWGLwLdYoWW1S7XjsTPLyJqNVarw0VRBg7zINLr1N3y
QAqDulTNrJcNoBvaj5xopdT9HMOimz/VkCpo/5Pte+d7wJCSauFAd6Z88rjWwTqQ
0iBBKtY7h71Y80r1vhqlwWxG3ocHK4wzgDwkMuEyg4AWHNh6dLpgG0Gf1stfcYCP
amAuDpfYYenerEgOqbijhU3OVxM+u6K5NZIpsobVfiwTeZCau+RAaLVeYAVArLpU
iqsh9Ixy3oQ3jHXsQ8eb8Zaj1mNBg3JGslevy5dUo3Nz05LfuJUyssQVJzqdx3VN
iqs0C1VLQuCbD9i2E1pz/jxafgeCiwqSpobmeBePC26/9dr8G0PkguF4reCI0zZO
mXIc4SSItL8evqQSbUWoPvaY+cOtnaE3bsv1AkiSmNs+TNF1hcgZRYKPSfO6IQ+5
wMkKGjygg+vaNywQX/NKtUpy+4t/xqekdqj8FsGpKOBDdFiPl4OIejK0aHD7PcQj
Frz+u3GPjjPebWf+QHmLpSgcfb7acrcgAZ8/BVHhLOSIox+WU0yAQJqxv8CZ7mV0
5UQXiHwHrkapItWjkhdlekGvQSWA2nLMo44hy8UFEIqE6RxgdXho5azsYX5MJhbY
TotJJgVWGgxuBb9bX+RkNL4uJFeAumlISmYfZq01v7GpcwYGaBm12qN5qVa6Pghk
HA6HbXCQUSuulEdwlhZw893FhOU/IlYsjASa2a691MsnZP95hQMcT6XWLAGQ1gD+
GiwoSKPDRhNjLIWbp8FzpZ9wSgrzKf3ldv8Kc2sNwYbRcNDyzhyOaSmaWzXF4Em0
F3nrz3w602wYzqSd2FlHBM5klmhuI3/4/qbOnMMoj/mH6i6ETpR8I18Y6nzkYBXe
QMfxt8MCg1sIW7IQ/cErFqOyfjqlh8SCZ/TxQuN+e3X387AACaO2s5IGdKAJ1zGc
ZwGI6wSVRoPv5x5Zrw0r53NHV5t6eY5F7PSJVGdzt3KahXIQI80brDuMBnAjINtE
J78CLyvz9oMxkXaTftwDRNIi0Cd9BrCt6RubQ8j4RgtcINAHxEuHky+m1wyl7s0k
YfEcRa0nrQm9sZbYHJqzrE9n394TemfhCishVnVMCJZa68sigG5vauZgFglQblEj
x910trECZYR29bqgAU3BTRAcS/yqTDjleqrTA0VPZfzPsWy/U+ZQ2dgYW8j8sbzi
KeV5pVCt7UCwwlDKDcYBLAPbPbBwpCY8EnkaVQ3Q1I46UHcz7T+KHJog86jXMbP/
/NH8Syc0rGI+uycgBBNC+D6YBNv5jN7FFMbK8zmvfzNk2wj4qWUbo/JcqJv8Qz74
3CVemAw770akHLQS6FsfVnZB44JZL6im0r10XFAwVsfhZLulAFE2M5aeu54mtejH
L9VtKm+BIVq6P70zY9+YRjMl729IE35ry8+Kof1k7v6ooe9nOFeqpReDKFaqe9p7
cxrYB4w8oZe/X8gmT+QFpqEFfw0OOHPEAH6GxVHhu412u8WE9T1pVENzLOE9WhYB
R1W/4L9/S0ObYlIzqiqABrFMC/J0+vfTVsm48xsjWuQa3mAhomBs6UV5OrDqyB4u
n3kkw4ht6eb5z43Gtenkv7cq4aE5/XjCRPpexHcwnuoHKWpCB7ErKgULXJRdmqpD
o161Hiea2abEukctx7C2hyunCEz91KFL5gDj1qE1couN9jCnBw5SwRVL+41AtrPa
7SR0d6KqI7kJ7pFpWeUPzw6mxiJ5U1BsFUzgUuxDS/QZ2Tkilog9Mo1cFwgAg7eh
iSEWJ2dJIc2e1SaNi9QSiysOy6/ysmPL6R9Rq0ZuXLc4zUo3KG/ss1jp0Kueex2B
6+FrUvG8XkW5xl5t3aG/vjeaMjwdgDUVelv97+gzUykJ4cggPsd6hKUBltu86Xz2
7HIgTtQshl3S5Z7YiHhG5QZwzHemtnpu+RxcZFDER7McyQJeB75B6zGgmZii2Meu
6vO0KdsaR3ObRdkMG7YYxWD5rw7Lg6YEjc36I6DcUFRf065rFtzA40pTAAf9GJ7k
gEGr8G+igPSPBphtUfmWWVkCcGzsdky9jkDlOA9dDa2d8iJLDTzk67wiHPNZ6NhH
IhhxZMzkeyoyizUzxpVyiOjm/X3nJCRAQKEgdb5MhORe8A2gp/dvi/BizcY4a57N
ok/7ptiLitfRznG2A8vVB1T9PAzjxqfwGBtMQsiNmTHL/N3f0YaP/McEFauhE8ZI
zp6Ip9+MhwTZXKnEtyci61EKhDF04LofbhEWGco2Il0/p/5Tmgk7tWCwe4VPu8Cn
0osHsAskwD+kq3OClvFdG2e8GoQnJYlyooT9df6ur3c4XenT7uMDIWKXXevZ18m8
oT/39h9c1+PTXTRlzYRvw2bTFhCBc7BWS9mafIbkMtANJlbpN1VU5ANK9Eos513G
vE6ob5Cd/JrF3/aajvElR6Wh1I//N2TdQJfzYDsPvR7d2v4cfT/2Sp1kSzNvrS3K
I5NcV1sc7M9zonkSZy+d4aVNRVN9CQCZnjco8ln1NKg/eZpzzQr+pBGNC2MHcncJ
S+g5gz7Sc1opkc85MYsHKp1rR7cITCmolkYp+w6KcyCXPw+G2SpE7IgxNjot8h8T
eEt80qNGtoJA7+TVdC6AUKFlu8IgZa4mXZX+UxqrTUq7f9d1FBh67UVlOv5f85mg
/+SnGw8/n20I32E3dggWooSg7Lc0HO7iuKHeq3h8ousbRDVz6dZojIyD/AqIbPHN
WSPm7F3BCVc0HHF4/rQD2dvvfVLZ7z10NeZiCivopvX8yyuGDQRw8vuHzQ2Jp5Uf
rUtw+GBNPB8+3ZO32GeDsZFrTiGiyyoaSQsdZT2r5jaf5Ir9pp2mBlafMhlaZVQ6
WdMzVbrqectETi59Xs41dE4iCaBL1DuAl04ughLp1XC+4ykM2TvsHGmc4hCF3SUe
Z7rS83/1+Nzzb5rq7EorQZAHLc/PfrhcjBLT233d+tvGIVoxk8QO4r9rvhJbRkMU
TDrY1LepXYDYIdyMJVaSh3nBpA76JtbeiVesb8Hm1VM5HRZyl/ctueRjg+GTnV5W
52GiTvUzUvYPHGRZHJSszwnCuILYyCwCl0t1hI8fZbWsO4mmGMYyfwHUsc9/Vbe1
ulx+z1sz18jeAIjvk4u6maFeWhY4QbmL4eqDGbRuQtIQaK33u0TuB0kpxpXOOEDP
ITsJiVPKgdP7Y+P/z5sfOsQTDsndym1QcoADvPLOB+7oPHq2UwHNqoVmA+lLqJIr
jUleDrrF6sKYYzX+voGuVH9BMR7ovGknjZECsEerj5NlNse2ZLYYhMn6EDdLjobm
zoWfXSUjCo/Q5wemHQvjg8/QjvkKrUuHRV/1+0PTsg1DyICP8fAB5mjNfj5ChvDE
krCVaiJ3QD6CuuVmwSoURx+TYegiiONLIeombUuuQM+UnjNuNFNr8KATINIYJXvb
gbBBsvHY2fuoXzZjjA9QHDqNUgenxu/Oeh6K6A7I9y/q8JpP0gKnw6cUsAG7bP2f
qEEFF2sfbkQNifRlb3ETwND0svMJRS4FVA99KRYHGUAhA8ZN43SBCs4cPHRUh/JJ
89z8tIjzWy7TP7qXCim5fmn4k4GGSwwWfiV3Lso3BhVD2OzV3x5g36IyQRMwCvDx
D0/WPFznuu8NJ+75Xebahl8/qP9u1oy4UoLMUXI0SK8PJUQFFV5HGnnDXjowE1dJ
dCKucp2eNqERCQX5g7rocY8PbfA+EFt8Fcl9ad6EfjVF+lw9UmKZaSdtD69HEKT6
YbZFtmzWqTMZJcUMlLqHUFvNJ7Vmh8xJn1tsq9fLnib5urBof39GpuAs5f7dGsu9
sENsobbpxbQ6yISW4ZXNBipK6lZar7oZiHIfPfSIZT099q9gmKSZvr7d4zjwBL7v
3tmRt1JPY79vv689oZ68urP+Vw7r7g1iN86huu03he0jgTQjsXPwsUH5HKofAGCx
xLkBJMm82wEE2gYp2otD0AUAD+2JaUZppaK0Y+G/4rg5XV01LQLP5NU/1bBvonmL
BZ6A4PQCywYAUuctCcOJwnMS/IT9GuPN/U8lXUFGWVoCEbY0JE7Qe7Slxco+RzlE
LaaugGkoU3GmeQB+xV8VHpW8vcuRuknUOTsNht+6csj19eL+hi1s8JUCQr6qBTv8
4iNU6fefUVii3GOo0NNTcB7KVf+IG0r26V111Tft9L50rcVmDnzEOjEN4YNpysX8
BbsF+84PXKvadkMuCAE22E8AFjEdrrYwsITYcADZ6wKvUWGXWnBMAxZLW2YAJsyu
JvY5cCnKrBXDhV70SrLl7SFCSbDsZp5bJchkELuF0ft2ixKZmJ3rZJQ8eA4oiXCi
+pnP9kTKxC3oDZ3jeRZ9Toz6tfgczjuVsaJcec+pTGqjLnPBUoYzgRqhckfIrJeZ
dQ0wmBJLN83eAWGkkzOkujtpVzwRRmfKVESbeemA2g2btcG/x6MBJcOP+o3vPmYm
54Zd9eXBvcTYIs36/FQgz9ld2T2Wi06L0V05EuzA65wU09TGm0rfuXFcYuUJpDUR
r72tVKZn/jpi5k/9kEKRBYK/mUquFnSULw27PnpLNLLFR0JGGojIhYM4nUvwv7bz
anXH293f9jrbd6ZMJqCYMs3FaGCQu3z/aK9MFv5yM04wI7t75jfbgWsmRXTg42mr
NkdEU1GdRSVy5HA/bJUzKi3oysmXZ/X1wJAs4DIG0gMNZYHdR9k073KRlkFlvgMU
ogFmfHaR5ZbVNJiFvBEInBUoWdOMcjFPt72/cFxY3L+ArUEQBKWRqFlJweW7GIs4
rJnMpmyw7+Em6kN2Vc2C/3fGzSGOAhBCQgKMK9q0AD/K0DU7AtVhwAKpaPfNn9V9
lyJHrw00XxpTCc5OFSW7t3sCwV7GWihybSM9QRBP4dF+LQT7G5fHR5v5j8ViGwNR
6Aw+q3E8yPg0KGFvjQXxBeDg/5tlWKh5hqwCuYLWgD0vcn+ZrLhVGFIp+f2uouSW
+BV2qXlKAWzck4F3xowM3ftN/bDiCEjIPLlhJXd0F4e+zavpwkwRzg8MevlFyOWX
t0WAG5sXwxOURvwUJab02x6/w6KiGjXHX7mImxY32gkOONzv3Hmyv+0bU2vGg5nK
8fWZD8DbD8O8MCjOPOLmKSRxSfj7V/j6NF3kTf8Ab3QwSskBXHAbE1wVSra9ZNf/
kKWQSrvFhKoqseete91ZgiNWJ3Z7wVSBlElyXIKkYtITUov4pLO8lJdi/U0otxW4
Cf7AxAj3L6m0bx+SH28MFkTR9WRorRyu4kQft7zUDp4Ia3UOewKbne80cuUE4Bth
2eU3unnXhurlaOJ/dCHkYq5PonVlivO+qREqyhNas2J1mGkGwQ+EfF1EyHdeNvx6
6rTAMmubVLsUKa8N00OxY+y2ypXdKYJ+kf2lAe8DkXbnXq/borUq70W9He/t0vl0
DoExop1T72+tTkZKPmS9igSafb3HEKMMyy5Wih9zhISRbITyE/0MZ6vaIs97lwG5
RqG5R5hp/Ci+xRbqVlemxVmkJ+NXtBGxsj8upSixVd59gu/SrtvpbNPD2tFbnoYK
IGAoAWI6cLYCSXR2Z1fjo0JYVCG8rE7NlOqAMVs321MueL0y7nbgy/eRivR3TMV6
UGOFwZunLxjfM3yfrso/Lm2M5uFS8PIIvbmF64JHVMwlzaIFRMO2gw1HxuPbe/ou
BB7G6Hd2iWZ2ZLGX2wT8VefNyGqO813K7EVT0aLiOdfj/o5GZ2HNDwQ47akLO7hm
dnep52gPD2oOdE7Wd6SRpY60KwnJRct2Z+ArTM9Qgpo0lOK8qvCVogAeEwCwjc0F
leDvTufYkg5cX6kQ4ai8VPjdCDTcv/xfb8eldTQ1aboNYbkv6pwUdGDdGXLV70Mh
tiGIVsPS8Ob3epOm7cTde1c3DlVC+zr4Rb5b5zNjy09oU0jMM6V8zWrkN7gtEQmJ
b5mO+Acpz6uSN+KAGUe40JisN68xFiQue91Q8PTa0PUOWSBtIipzGXvM78SVZr7o
B4cwwcY4xDaXG2ZwYD4HF1jU/OLPLeScjQ9BTelABRhFLCoyiupCrtYv5n70AnEU
A1geL8WtQKVhdlwTM3Gc7DLVPNAGn2JLKYJKRzLz5tErTgSv5yhhSXzijwuM+jQG
cNMZtA5TQFZ+uZ4mhOS6U1dOsg5ev5P+pt1EvQ5kECBnnX71b4br2c3E16zbzq/d
r2BdlI7aU7ILTMOsP2eekN6poyLpUzcZjLgLk9syL5hFBLgury2KXfUmR1T7tEbp
DppBlIPAtTrCh/YTHdytb2vVe4zBvrrtWVH5GxalSE4X4QWIKXNbFRoVVrYN0qba
Frt0PyfXUU4+s+X7tnzeg98u/D+1ybWonGAbDN96OowwGJn+u5fQ9ga+FRinj1dR
TMw4D3AvIIqWwSxPFx/NyHgtuTb2WalrammxrZ0O3gZ2MVaAHIk7xGx6ZN7Y0WJz
QhZxFwGnbdJb0wlgVS63H/eoKuyvI67REQSdPF/RS3Q41LL/jsiloGhMH0CWYaD/
qa3Ad/DBe4z4DenCo3j/l+vaSVPucuLrOm1vSC9UFbQQ3dVrjXBsXOTXhaTTFQ9X
+p9jjLu+TioiGa9WvockUxRDNRIM5PcK9ZM1NeKaK7ueHMXRdwqohvkv61fjuKQy
tPxknE7Q/ASeyAT5awlgK/9F8PJnEJW0Up4+W/TpwzKwM0EEl4W8dsMRrXWJoiQh
vO6HGb4PJUWWitfGUISagIraA5wIyBdP51M8k8EG9Qh9wEydbuBAeGz5AlxmuPa/
un4XDt5QIis+av2TNRfXzj5cCcihi3uZ2ANN5NUU/F944sugNHsySJSuYaBQcQk8
imbVMS9I+DtqrXoQGAjQ6Gjli+uOgGI38Fw2sAYTwUHDvPoOVQFeEJRLBjzxvKbG
wxHeD7cAycior8Mm5Cg7XN4aw573XN1xdN8n+wEl0wAtlyS5aAjcTz1yJLyRmiO/
X8hGOZqpuIYtSSmyNYX73pTZruLzmh7jYSOM+AI9AIiFCva8kEcmVCCL3mOjS0Pa
fDxyiYL3C99S39LWz9mtSb8TXiScB2Mijm3wxKm76HRlY/q4QsEd5WAEpMQQBV+w
kIKjDubejpKtAGp+Uy6FWfn8BMces+S+GlGPDA4IV8ocg6foSb1vuvxU38SoHv0K
26qbuHHX/jg0DCG2FrY5J81zkfI9MoCmiNbEjY5I0YpEDM/wSXHEO7dMDDuapmz1
xLjOw3IQTrIz3VGxxtUVc7NpZExru/d34xlWqcxQ5PaMgHrFcq9BoMNIRXooN7Rw
fABisZl4zhb0MCgFzQueX484sHsZFo3CQNXPOXA8+FQzzXjtldJTEzQPhv11IXSI
TPrhNIqe+wQp4eCXhPssVCPf5rr5uKXDx19IN7JGs5cPUWbZJblFHQLfrFn5m7fu
/BWcGPjHjow6VIBwWOw66kNvS1AoawgCWa8FznRcvSKdxWBuKk4nibWgV2I/Mvkl
52xbH/Sh3h33FyUP7HG8UXf+F5fE0nUB25BKNtOXlpakqrQsl7aNZR7kADTxMkkh
ZoMcmpLxdV9GjFXukJaCkpmsNykzlC92NFf6vgAYwbPLekoxGwnWLTXdiJ6Ooli9
6AOJIGaqimjDGMA6ro3zbeWZCoxnjdHb0elb8SCtUlD5wNYZvx4+2Z/I1aMGx1FK
hBRsCE7GBy70jfEyJEyL7o7IJJsryu+XpTp4lZJe54hUV2Uo0QD1voWaEfWTAdP9
/LBcyFFxM7xk9Hk0LtzK06Pcqs7wFZGW6ReIjXmQnwWsEeWkQw/yCF11QHQwjtRS
mOkfYsLbh7zoy9vj+r1U0afwS05p/n177wyVzCvbPM2CY5sp4X6dGG8UafdDGVyg
BDvLrC/6JeBYzE3B2q1dF2IhBr74GUweRYSJNamtqVhYzRfSa46Sn1QYB8j727uF
SHkAeWmzdovGGkiWvGgVlyzLvwCzQHHC8feqEAytSgJ9KcsDoxqMS2Yvo711ETVz
V/JWb2+T14iYf1J6D54W5OmfNiw18jhBOpjAXuASbcDemzpjRQMX5YtriaWJTBZB
k/9+je3Q0wF+Zdylu1jx8IAcuR1nCXAbGktzoFPCZdxLGGXJLfmFVYf0avOpQIPP
3tZeRAmUyu6ZNSKjxGW/Cif/+XwHLG4f+lBEd8LSCWCVoGFTfQG5aaG2GaW9AcZ9
c7oJN+PR9c1iQ99/2ZseL6giQvE88+unOkB9+V/SuzicFXdi6uAPKGTgKt2bW9ge
rbaSrv9oT527GOWmVXQV+KCbTfsxJ8q0GIMRdZpMb9FfF+W80YPjm8KM89vOnZ3y
cd5VM0DI2pY/8wHdC3TOo+BiivWxfYiC3Cv9gra/3T9xZDS8QsKcRudXr+egRRAI
YMEsApGOzgbziYL3Fk7J8iDnxsWSPdIVHbChedAI2qWO/YVnPQlkgUAxFtZ2nPTK
sW7kMcwv1jmru7gPCqrLw1vk6byIhWl+1xppn9A08N54deqm109c8IMpLbzwL4TX
25orcRViQbptAJI/kBlI8CpPblbcMKEcm6NkjfrGZpOEzaKfMhAqClMPeVmvnq5l
Tld/Jvqawi4oXJ3c6Up4ln9O+L4uok2DQAKjggd5zlatzQNZrTB5ahPVhb4qdgfL
BRU+6Q2NDsWUaS5JfGZ4ClnwwRuagJRFWbgfl/8Lk/LOVE/bgtJHvN3Yprqu1vo3
mXR4dcdAKwNTyUQYlL85NERUeHUc3hJDCy2D1AG4k8QiPQKqfWpqolD8nkYr6vjy
eMErcERsqWYZ2hIzYSR9HZYzlh+ZD6DbTWzhQRZfCMRtj46qjW9uk7lgYLSYB9vz
UGvAup5q1O+gq5PSj9IpKhzx/6HhFXa+Cfr+eIAwQRI4Dt7pAYXgsKZxuoAQCOeG
X6TgazsSDCml5nv/QnNR3BJb27n8/tDpI5eOp6Mte0NlPCprD86OBD7WwQlFFz48
ivyKBxC1quqhzxj5t2nPBpmZTJm3hzp2TKt5B7W8TlE6rYyE5HdaP7w5KdZgl1sU
TIW6IHkqcT+4ci99Vp0YZI49Y2kt3QkNMzxylppXXwEwn+KQrRGnAn6B0tDNsbAU
5cUUf+gVuN2IL48YRp81rVzqr8F7CPZWHx858nReyzwh4Lsgy1zNrlNlQwPZQkk0
7LXijyA3Wgxv6gApFLdEMMjfdR7cjpRkq6XjwotELJlwpei6P2hwIOAJFxVV3jMx
CtnaCZJFKZTzA2n348lvXThtIioFccUnfACeUWzCpO1t3KQOR92zP7NYQJZYkgbP
GUKLFh3CZceZ5XDWX81Zl0HCWhy3J+Dq4V/PLIaMcy3Oa4hkZyZzHnqPdztM9b5m
dy8djxAZd1fN50vuPnikus9qde/cyERj7F0zZUPrZNB38etsRphgIXJB1dhqGHim
1lYAQXcUXPOBhjJ+UXoMc4CpD3KtB2LrGVWg4/OiGAReHJBHZsUeBRWfHwwwucGM
1w9lLt08yxWBrDUPwFRSOj165HvsfxEY4nrzaHK18/+bxGWlZH3XN+d/Vti3dXVs
X3q6otDpxZ5h3ADv9BjldMgcMzhhZHBEfWtD/irlscoskM2JXSafVby8MJ6aFKMw
KU1y3AesTz2KUX+DYl/LnQjJjXtdToqVCFm0qFqeHjsaumC3FCoX10uYBMYO0vD3
BzyFEHbalT3sl1IHkVk2/0VQ+comx+1h+9b50Revb0mlasTjR9yJxJJOidlUAgoG
puc5x8h9bN+LohT7koQZw4NdjFjgfH6bu35KEmXP7x1jca4OIQcp8blWwRmKkfSA
Rmv0eTIuHb/AQbPh3K8eEglPexkWMaYqPvHWY+6+1y7nVTVkLWde8Ibyp11c7uCk
Wgu/znHY1cPQffbMr3GOyhPJ7O8iGzbWwDslbkKmQHI5vPz/Eiz+NOQyBF/s9TC3
OVvJ3u+4FcBnbl/zlVF+AO8Djm+S3VStwFHJdNlPyZWVJ5wqj9qrqKigPWaYU3e8
Z2cagdYxRnG0BG0nP60urgJFmaZxJPyPxcQ95wZQ2udSYde6Gz1Z/Er3cqHW8RO5
iSMnQeBDBSZbp2eFex03oGdrVbKRmNKeaKdaIs0idnuUkGdYjvLQaM7SygDMIaZb
h8cwh0T4niH4LJJHz2Hf7XLMy0JnDnQj5vVy/45/lamv3yenDXePKIGG5cnvTa6U
FJHyRB4y9j/SEhIAW9W1zwINtB0nJNzeeAAxwAC+3lQFom67KDRbN1M8VmOEmZPa
OLNbfeH1viLI+CMP/ZYyOqZEaKgy3/oo7RRYOytjrgg2Mq7CBaNH+ulp0dnH46eJ
H8/J5pYeIuR3Fo720J1ZBqwfnJ9DnDiaHJTzkHF6RqrPFVqjkt5RUGuOiflaXlO9
4HR5+tFcN7GE9HLyDo62EIAoLm0/bBQQVEzy5cnSVQeEEcgoua/HH6/5evMSoI6z
z4cv5FQqlNior4Ii/Jk+dEd/yXane4N8WnQb2ofzorXGRj5RtPxS7Rrdia8Keoes
NOE9fySafe9zV+VGH0B6BP2Xs1NOhA6SfALlUhJwNgoj31Pj4jZbn3M++X0mdMbB
+7Do5DfIp/3W7fcxP0WlC46idb8AzLb8YZthLL/gHrwG2pC0974g7PrZDLXauCl9
GBuSwRPdjPvoCVt2G6WXKwb//A9EKOr6yTlZI9u+2NJ6bs3Cs8ELY/mt/X4nBX58
JdywEYYGQ0Gc2d+KGNhBztL0dgsraFHJrC0hhLrgt+2AHEVfuI3uTRQz8xYirJ/H
XvjhRLlHlYTaTkSbT51tAgzSUdVLVQXYHNIywwdB80Hoq4jA46qEKZ47RIYb+BjU
nlc7Ym59CxEoh0XDHRtD2ueqbwMc1AMdyoIAL/DURQ5FPuUBa+O3Gjiag9g3dDyf
HcU5RW2fuuA1HoUZXzF2W3qXNg7CoWIz1EPwm7QBLu2Xc1pstN89+8iaHGmRS0Ef
ykE998MPnEXpCSwXZN+Anpe2iBlJ4Eo1DLq82wREkpPdNHI5Dlt21951QHczwyUb
BTotbtf1g0pu71YW1gsxvFkWWP7CvQJKMLkG4b4kHKxhMBQdkDJVViumx2jyXJw6
+7XdWx4R4RkoHTPUDja6/AY7FahGfxHWUvDYfFwjz/qSCOe2UiOEpRoVuFXwfdyt
tApms4Ry10KoVsWFKzH7tAzC6D9S/aQDCJlnn/voyUwxVWYdQFwcPT1qXHunahN9
9PPUYBwVnu+0KFLG3gs9453g8bUuQ6C3suwZXnBmKU3MXX7XTHDu4zpSgKuUZG2b
HgjgsBYABELnUzkFZMRpMOsMHS3nnTyvOVcDHTYkBGDgOpJXFp9gW9v0RG+9PWth
PI9LJjkQGWSZj1+wfKT1J7Yvjvgu5IBPDCpnnWLZNr60dDvV7CezErM2tM229DO+
0p8pg/SeTE1UeDQOIxpm+MxXEaxmpHPWkBpvEfksCTpfG1DdyoGwBgVsvBEoN6Bk
BvbYaqUlmrehqlbJgTljSbbVgHUpxp8SNAtx7zMyWKYXbbpqRKzyk5pBCrZyUgut
cSmxjlWDlSB9aPnoWCKVTAS5/h1YxP0sNdUgCQB6OX6hsy7pTcdXIXqh8i4zTKfh
yqgF/C1v8rH3l/UtaC2Q8U4vxgVjZqQoR1IMwXe1kVuj6rwAg/apL1Qb51AnfQPo
OMwVp1kkV45yiEmyheCuI66SuZDkw+lUx2VLv1H4EuA7pi9Mix3U/emR8wNstQke
YZITvZDo9KMzhQyEnnRv9JioEmvhArVG7z1wHc6cML4XiQdpaUAJXfOco3BZYim8
yUoBtoIOxzAqpYXxZQpt+EGUbidW7thWO1qcXh9EUz0oqGrz3T6j1N47FHwhYgJO
ahZvmeXDFKgIMdgrjIjgpgd6DQcnalA2p3L3rqQu3tHB9YPukXaWlY10yNXLUenN
9ZKGyKMacxm9xC5o6U19p4mJv3jl/iw6jqBaraI2fYuClVkJPj0QxONpgZM01ik+
GaFRHyk94zvHFH4HgugZ3Refey7VgFABAc6Ogjj4NOvfRV2heTif9Ha5hnOC3+pN
/1+lNVDGvEApGFsxqoZSf5HIsU8cfhcpStlbaE4tT6YKnJql+4S6aLnEwKTqRfeH
/ReGGJP5fLDDcddfcP9fUHI8O+vfStPFmsOjR0UWqbDTLl913xCpC5pEkBA8Vdcg
KPUiUlRR+DwPWVGCBx0Uz2mhU0rcGp4ViX2L9AGIgf+uCws5PA4gKRpJa2Tn0QY3
TwxucCRcWTkQr3iiM5linDbAq0AEUY2v4vf83h0mg7nHkyBbpD1w4npV4xbKA9O/
JBM5iAwnGoKxIlW4WFZlmWMo2gBt9qKnPrqV7SSb+UCyNtAQd/Baly5K37+oIBVE
VnbtCp3BBBTGwnHsEqkK13oLu2qspgYm+98Wm7xjNeqfTNulqjYqCWFf7wg0kLf8
LdVe7D88m06rZkoIXXabKK6MdWgib9ASayszGZquHOtGXORyBuawhcv3WWU6ib8l
W5XMCTr2IaaniTvOGI/hUWmw2ylDFzbySStk2eSGtRnmGaVXgxCuQVHadB1uFVBB
H86fAt3U8n8Z4iNESs4yrMxdCTNNUyDEhr4JbfATI+njXcKvD6Zhn3JVfxHH+9op
CYeygDAMMWrY3FBKTOF5mR+njMEO6xZWjpTUCUwP0H5QdTWi/+gAqoUaUJ/jF6GG
5wLn9SQci8RPOFYuM+2IrSsD81Zh4kPJtfVQCzrfaT+hPDOvZjv5wnnvlW3c70tu
aTOXMJct8QjtqzJVLaslpY0HgSwOg4+TyqXJZHEdcsg1kHXUAFTaMH0Cg74spSl2
8To1TknEBuNGiCNO1GG02M6CYxLoDDgZwsjDghNJWNeyIUTYDFj/Mav8qp5EYSlg
n6uw2iGuDhffjel7mwjUPZAz+6zXMf+QnmSgudDFFCWMYeDHti2dFyso3AIFy9Kl
OcsmQEM79SrXLAEzlef3fsHjOHxhECSg+uWXm7RrTfv1R/w0QzIUOkSFOT//sedm
NVrSJFklmgqowdO8XbsWoH5KoOKeehyRetCh5WKh6UsTE5Ex8vqJfHZ01VrsrHmI
eOMOJPfa+FYXUejck0pAAKmx/FtvN3RF2aL32YVlO66UrJBQZoFhn+exxqSbrBi6
f6oYs24VUJZry2oafwyaq9adGrLKu9YVs+XO4GI9t4ntNXaz/FippX2m9I03eijS
13lsiDtNNtJqmyjQRH16TGIuy0iH+ht+xAzz7jEGr0duEq9/vmI5Co4QV85rKHpM
6hATXJ+5mVbgst3hVxaMWRC7QDoy+i6Q9UNsIRWhGV2rdSgtU/FVohq/ug5AJj+X
9mNfgWF3v61sE3WUiAYEk4HHJnLaWSGxEDqYpEpVYVe4HfvPVbN9KyhPX+iZCYIE
GPg6MsZrnZKVsUZqK3NULk7aNCspHCNz+kshSrj3PUBFlwIOk3mc91aDm59fTKJn
yXrlfzclozBinUsuLSoteRqHLWXIGAXGubEsyn+Hd2DIrDO27H7L2gUejKtSeLMw
1cB5i9tZEiHrMzNIgL1XhqwZFZ5Qq6GhyHa7Uoxo0BTUrevri3qNDyK4BGYk8K4a
AQcYj2+mrIKfe7quQlRDTEdH/OhHTHGV1jDQWSB5AexeA9ELc9vv0N3h+of1gFim
gP2rvJVfgn6WbcFYOxTUcQlU2do7iG/QJgjWQd3ZhPKy+E+4XIHJEdgtdI6wyq6m
1wcwb4wRpwHKQI1dSxwdx+BMnyLRx4xtmG/UhfG2Iqo1160XIk4Kiy0qcvQ1Vef8
qX3JBvBjUU6e7n0hLLzslAf3BZwB363MjeqZdBoO3XPG6FjhqLioZRgEPEzcFQPN
91wvGuLUBrSLAgU3GMKtHq2zN0cniqI+UifP5/mukgiswIYZmL+IJhy78xgvF8o9
lf6Yb8tQnREAcdLJIZKOUc6XK8Vmt3mA4xD1qdLurDepC9GuYaAFcl4YWvDuU12P
U0RbOfvZ/FrnPKG2ijl4XS0CdTgWBXetSI/0YrUzBisfrd5cZ4Z+Hy8/Bv+UA9YQ
1j26Lt/n7f8EIHrdMDn826TS3jK4ZM5e/VImx4+iz63DCdUriVsMX43wggAGaKgD
BKM2LlHFYkW6Gv8JNHfVOcibFcRkaSnMFCO9jS75qyMZr/0WX/i5bLWo50ybOd8v
MymRsCFXWSC0eeFohCZfUDxJvUJWRqObkpOzgteiC7PRrD//oYSGU1RuDvepOlzL
isnoD5bzDvxVAm+NCQXmOXCujlizjosh2zeYvNgx8fTAVKLVhlqNEgGN/oKQtzzw
B/iT6+DnBNxR6QY9tLELGz0H/NFgqNRKs7Lirxcnvmtk9BNpdXyGKQpZ7Kge4LV0
Mh170QV9KK8GXBz57ehUmNtIJfv84hj8d5ZFKOUpWzvmInOvCjng4cH5uFbNg2Zn
S1HvhjYU47a23WD7bxZFjKA+qQcT6hlQXdbT8WDV1zfk6DciW7ATa2ZgKqH/W4Dr
NJsubRtDQ8AsLoodqMXJkDXfDj+K9krrSLTSKNGQk7tKNUolCEdSOA84FWwI8ani
/Ev35XKbygBA8bKauHk5eT745FTLaoc60lP9lOyEQdfZZ88MnQwfZUPn2VayyvLQ
JuP/Ej7lJQwqRTRqY80QurTOqe35lsxjxLCm5XF0fiQNR4l/yeLwFq6G7Ag1Cqq9
yHxu4rT9QxxSTb8HRB79fWpQTtUt5BEixxRpRRo1E8FVTOIhkuWAqd1IDoxevdZ7
s921vd/CkZZj2C+hOs/E243Ls6OECkSeKh8su51H45jMD08VxuuCL9tbulWbQ2Rb
0vt/C+KoUoyALSoTbsuclAVY35zPWKsCsNywUlNAtNxwoAXjurUs38ytv85c6PJi
Ze48+0G7GUeYG/T7nbLkYX6YJ5weX2Q+bBrduq2Qux82WT1I8INtRAC/ydQLdXkI
cZRvMm2uGEy4QRaPThQ1KeqQ+TvkzYwa02yJra0smkttFKtHxpFwWHH4pLOjrMue
ichC6ijy1GOMZYc6+yzMmk+iqsVAm1xe4NUAaYe3lYT1IzqHNKNl/nI7vczPXEb/
+LGNBjLZ46ZiCadNBcfohXeyTeLcTEoHP/0D6Y258GmoBJm80bDtMP2Yne9ZWC2A
XsjyFIwOOT5ZEqTOjQCFf6bqYsiL3ymWTit0NWW4vttNi5iSJyYlmer5M6IFZhnF
wjtnlWt3DjBTmQH3V6sLB5qYySfoUkX5sMFAnzys5gLDSAsFANOvDn+5ksgr+zQE
G8MbcFu4Sc6LoykRjdINa36H96POSg+Igw6mlwOmglPBJGGYjD65tYxDW8fIKW7B
s65mp+k7NTiQ4mWcBEMULN6smT6/b5GO7MD+Mfg3sUo+KgwtPiOivmc0QhCchLD+
Wmcn1+uZ7fFuIRFm1AKtD1N+QB4/ztbcl1C87qjFYMkAR1mUX8AHH9msBqU0syrU
sRYEjinnYory5svexuipfpz1E/G3Yg8/Gig9qHliIXV4qpsGkolgorzW+xNWhKF4
BdM2g5PK1J+uFZmleqpEYoQOZN66QXr8PymL8jEoB+XIlhQ14pO1syujkTLwyuo4
SwKfqye+oipsuutlKBrk6H/s8loeUs6ZYLmWoeZ8QvOLVbk8C/mfUgN/1e3vHt6e
vnHbuYIpbx85V+i6axRzuyx8eF0ntPKv62M/TrJm8JYMnGEpP3MW2thXzfTtrXvI
XoJvwixrBGqZt0f09dIjQUnwHj0nRzYmruQbQqvSkSWbpPMAOHQmLDaMDo1Q/bUz
4tPQIbaVv+d4stTLp8U+9xP+ow5bUhARGyRIPqS7qg77TERYnRwrTGBBBqbboFrs
z3fISif/ArwEuMVpiFEvCdBerHiu4OH1n//LdUlj4ddBcYmNiZ1Jn5Qn8h6t8A8U
Yjif4M2MCQ6HPWh2FPqHF+FbZiFrBccHEqtNOIxhgO85AY08+oD2trReNZnAQf7B
1R84pi8Bqt/QmnUi1WHsfVyLdV8Ib39VOLDgZm/9e3Fslan0NlJH2leqczZfo6kD
sOX/+Wa+AcngoZRQOe8R926Eg8qQt9Ona+lizADU/GB4kNCg0jL0ZGMXrLYCWshb
3gyLcS3os9DzpvqYDfiYvapxhBjTBal5zphpnC1YOYkEqKSk5jmm46hZ2aoogBbP
I1qRKWvIAad7sTNlJqwi/XSLtUde8ioNDEfxTthpmc9RSdzlLM9wewu+zPhEIS/p
oglEbLlnj8jMxLUY/DPYvs6R0P7jRDXj8TSyEPSEkA1u5xZzo/TaDR3H4n0KcWVV
ldV23SQEeDnwGLAkhvDmo2lLkbeHsztimh+Y8OfitpKu5U7uNrlHcRD7HNzVHqxg
e3OJyNUdQ9qc1skqmf3ihR+ZdazOgURbYXIPGr7n5BNVXtmcTXf60IQAL4HJLdbZ
WUChe/LSxy/ILiHLUhHxY4RCb4GSELdkgcIXnisQnc5+dOvd56AjKDKqx3XJheQj
g5KRXVyiOPWJgOrwGGcByv3d5Rhs0fNVZpi/wDGRAvcQ8wOxijh753xf7hjV/Eab
EUsn6vPGBEy8IXc/U83PFxL4ApFreeWMxjB4IusC3cJbNjp2e8xc3r6RgyiWhPV+
9M8MfXtjYnYM59mou7SFg1FG6FmOEECL03J64KBIC/unq7Aib2jHtwniEeFxcHg6
2P8tK1GCruPtJ4AYcGE/HnHQLh3s4Hvftf3jSpwX5f/DVIIq7GXmryD8vyhQBFjg
sw5w9FJ70AjRXOMvArlB4we6l3DXTlh/vyYzhonpPcv3PPVWvsDwKwqZH2X6ieEQ
NE2nGbFwOi8wJmupuj8BCI10VwJZnufckBEW+8bHxCs9RSqEj8eFGxbyvMBZ2Erf
BUwD7gHnxSrTMNa/oaGWfjCznvXcNQ6l0rZCtgmYvfzX5H476RxjtRClgsLYt51Y
Fk1aMA72EF8jvqErppWldOgjJw2iRgffFSYMhrNkBdR2+b/nB0vK0WYmCqlaH5lp
PlhnLEBjniRLQtO2lQAJG8b4fOOotkUrYH983VO/iyopCLsPEz1hmF0i7vOuRWqg
iFoC+M8MMuBeMk8yopUcZZ5K/Ye2n8GuQTHB1GgDGBmLVbX2phmLOT0mDPMGVEKN
pzKQhN3fXAXynQMReah5TPuwd3QaC3j16gwVMdPK5Bji6sAsjx9Iw8xDXrKManMH
SLL6T8YnQyctYVlRwYMaEwbphQyryag0mrKJMi1lH9hlYzHTxeit9x3lJf0C74xN
Mb6f1eXENIeRAMvkRU3QeoqoFDwLuWM9ZVpE4SDKiuLiCsj0tVtRqIuD+zg5O5IC
D7nRVpoRy0/V1Rkik6QC6qZvTdxLe/I7G/kTmE3RzBE2io6S33SppaLfPjmJeQ+5
4T3PWx8HimE5PHh//Nq3Nxo2OcYFGssWM+D6YKonaZP55PYbmBiKOe/I2lVeKSsB
RNwZHR68Lgq/i2FKmiaZnGPmfZiqud5Bw1i1NXxKccnuRsCCJe1JbAEDmjCWzi8q
aM4pvB1S+PeTupyVZb1kEA+AZrOFVVtueBX5QSgWfXOVjB/GFt6Rr0CNvHWEoF7E
AZXXkFHZDfJzXyoOUIU+8tQFbMSvgfGFaSgU+HaGMQhJtwPJJfegMulX+WEAkbCq
J6baFdVgs2a/CVNcx03dvLEehy5oykGQ5LKXZLoImKlsVC70FSK6/XQf4cYPoaqZ
90vmJwby/4l2nqdattJFDyJe9Kga9tUoKWD5yC7HEdpcbttLgWvwhifeo3zEiMq3
S9nVveRZ0k1T45c6l7xCwK9DDfo65CTpWuBOIcUSZmbTjuZPFul7PyLjl3mAdnfF
Jd7lMJHe9mEMc9BZ6YF/0nTbc61qURrL6Dxc2CjE8P2YidlB4JcZu1sAVGIn8Nvh
KHVCOlsUudldrfoQkFLkYghs0HBm5c6guLHc+cKukyVIFf16DB9ROTb27ia3VkDG
pk9Qy+Vtx6H4rjKZLEb1Ds0fuIBln1tPka8KUDoS9g1sCCpBK3JQbtsVCCAiWwdg
btmbUsfmP0J63CP97a94cZS0K/2w6YRa+pbLqZcDVljiDr7EOQOtWf+oVg1Xadah
Y9mdvv94KtG/K0DVXe3/QXs1n8xCLOObDjXkGDKqn7OyySPHgAJlX0cFWryIFGzu
n0WNKB9VVkIrepWPFEdnrdbkUOwNgqXFLZ6hmDrIcU45wNZn8tSjdjNcC2UpNyZk
gDl4pTb+rX+8fPyfBxodeXVMaznHrIU7c/3D3bmpGF8hEZ2w7ws5qJRzA8bly778
lU8yK6hpxdOX+RL0E43IKeAWRc9XXlx5i18GP/GjIBOlO3isiKYAX+NQnXKI9ltC
fSeVk7YEtX5wAAbMlH/cYBwM9kzXhoVraW9+U4ho+8vf4o160Cl29uLpG1mPJ1jR
+b1A7qzcnXaZtQ8il2ACO1H+XVOTY7b9DtvSOEdDlRSuzMFmTepIW0Up7ptPyO7m
S9TXvC2CFnZVrBGSD0ujGFwV1Jk1p+05k8kbiccI1zHwlPUEhzVNOe/H5ozJN4gL
pyvq0n9fxaoC9/JXs5fW9wkMgvSWAQObgGw8erUslyp1O4egD0yI+YLaGNCI/REt
gg9eotSLaD/pdgbMJS/GREJx18wglTlDSx+knO3EplrsPDRhZMmbbf94MY647aEa
7yCON2CCoCSBp4u/6v/MKvdfOgByWQY5LtzO6rR5w7T887PvN9G+rbB7MW+bLwuS
dQdKobXG0qhpk0Wjp30l5HjUa4x6uYACfr6QLd33XOIlW2c73ywrE3Vb2EeKCsB7
Je4VPFnQQHbVrqW43F0P2cqHJ6szfMkUH1hU4SmqzCHPuTSTl7lJTsDIeAEJ2fkm
gYdVcikYhGaPjiKzG9qlgboq2X3ZBFMgl8413IkAi2BL7xe/3bwLnztHMblWw6tQ
vULBSBZpfsY0F/q5BY2lPxb5aVJnXnUpzSa2ViQID4ktW2kkehMzVpBq+Jc0UOGm
fJE6Ry3HgbDUp0jT+7oaFkV/JM6qK1nBdWc8n6HiyzC4MyX48/9AtUdObQhkW43L
DSyqUUpQp2mW0PDkJOGiApYXf8lWlTyNQncLMtuGip4y6cCaCNPgC2pXN4B5HAzC
MtXY+RvLNcOJrzmQdDYAs3QqOQ5VffrcT+EhJSudohPA72LFTKUZJ75bkILHsHUO
SLc7lwXValTw7Ee3uqzWtervslGZP10BZkdh8CPo9O6Qkld4fthl8ZNekjcApRex
TaWkWhcyKqeWJfPF+9p8wuCFpU7IEje7NHvp3AD5fQEf5yWDNl4HWHbLWFjyLi4v
vzwFE+WZxY0ubCHsdVz2++BxN2r68qLeQGvt0r0B6yOA6y/mTKawuD9p37GxFo7a
EnqU2+fr4s3cAN5xNvBw8rU28b0d/uywLNC8kzt1K13ovn1J2qrdn/CHsBzxcyRG
VhHWq8XYYNSsGuvTI2mUS0XqC6LgmDgMm5phsY/rue1j1it3rKOwOK6uT2LmiQsn
+MK2LagdTm5+OKIZMl29wmg0gcz7YiQtfCKASJdUpeZBJDGbPJD5F2gbgyRMrHI3
pMjqjm20Q+JDZ4r8/6LH70CDoztg/4/lHzYUKl+d8RHEp1EpbcbGPj8pJucO+0Zw
ZHZIIqccpn0x7Hfnt8qAWR3GrYT+GBehF2Nk+db5F/RcLOFJG8bvWBRbQY3CMRgb
CNBuNt6Pj57C6ZZ9o5N31jqXXgmGm94Wke8c/t4JRfrSD5l5cQlDAd2xdZ2wdt9D
NF0k+qLigdrwNJxhGqmpO6O53cyaVvnR5JHtkXN54g2d92Fgu67q4xVBVlj3/jir
t1b6EFLLSArfOI+vxt4OHrZ3dYTGOYcLI/a9mslxDc4PZ4IOKaGi/Md28Xevm8wG
HztNe3bR5AODAgeFaV3ceKVPCtc3XOVn8E/75AYfx4tpF4aNOqmlBHqwXUhL/jem
gLTlNtbe4W/XokeAkk06/rpV+Qxp8Yx1+ZTVXYzvENf6ODEGzDbDCyT5uXkaX/aS
4LrnQPdHlla+HY6Jdxwf9zj91/NAClhQG8PLBlyIpHyh58Fl6ejNVfk/4UdaCasm
5CVSqBxzb9l+T9fJW6FxTZTUSSYLvfeG0ZzpStdG2anPf+Dv4LpwGh+o7INKCNeg
ccIn3TjK1/1MkRcaSXzpS62mF17DrA8HyKKyVbtrFxKWHBfVrjDLRWONFBCt2M+h
YAsUPYnU7/W2xChhymfrxRotmjxwbXvhWO0yTYX/TwmW1Yv2Cmbq5UoEK15caCk4
kfSBatql/SMtJw6rH44YNm/4xocWwW/38Whxk444oeupow0kE2Q9Bl5Q1J1rqlRs
LZZd0d9oS0a6itcFWN35SjgoeVG3sOroSatIWbU1fnRdSjWshco6RF2gLwEpqxfi
1yrQQDJwym23MdNRE0YhDRNClA5ZZ65HzsNFZkUuH2tN/oEOBUIcpTovhWJdvmfQ
otGi/fXOTwhB3J0qZUqAsin4/k2QGoCiR8eRmhHECntF71InEoWlxz4LDCY36hAV
8A65T/qTh+y98AnebDI/axAuWjZZBtGS5C0sfW4zVxyXWzaP+w615OrwUSj1iUCn
ois2pyzXvoBPls15QTdZM+I/AzYwhHKe2qP/VvPjqqtMvSswVLJWaieF46tQi3S5
As6lPgCvSfATkk1jJGrOJgoZLcMQvN9u9JElYprpwQpkym0QAXcr/tT4XD/Ifg0e
eBFlJXkw7QplckZmWPAKpRnsFo8Q4NF6UlgPieK+es7lyWhfhX64vgK0yz9Q8RKu
A6Ne10ND9FPxhrUOtHAraz4MA1nn74XDKtJf3BrNaYP2GI4K6/P4EqfkdEHjLmSp
dC4YbCczUaL4lEKZjVO9VY2xsk2V9KhfnnP2JovyVxEVBC0yDWH71yPMXeYBW9eI
UUrCCuPlLrN0EVqwW3i/aOiWBHV5gW9g0jgqrFv7dYGSFBuKqdU7SreELJzyz+Af
trXftm1Hyzqu7agun5ImEczSE188JY42Xajvtm2WjZkN7ulpzGWmKs/4MnkbBsiG
wFpEqMaZsibIF9pjpdX28fz2n0by51y1jHnmtqj9dYrXvrpy5wZQi9AalXrIR13P
/DHR1IkOfi2NFx1Sw4stQafJQkAI67QNHdAcyCA4AqvqK+CyIdwciZYy/vxL+DDv
qQqqxDmLkkF/diSFRrt66jF7ieABavmmyWT0UMaxZqmPp+c+/z1So0fG69SzPyp+
QCDCMliTNNzX0ELxCqXbVMU6dlUL3NtZfXZSO4sr+IMWFAbs7s8quelUbUVbsEeW
UcqImR1UeYy3xJLrjAFJ+WprAWB/CeAR1Hflwucz2/w8RUNfick/yN+ert8nRP6Q
a5RAz/h3M3m2pjHc306c/3kwFVRmUjrUJI1bYLNKgeDMCmocwo+bxugK1lncKFmk
MBlGeOCDo2/7ChurccnABJWTMKeLtRJqQIwWmTyVPJmNg4LU1GQskfzftBWBkiEB
19g1OlA6Dn/SxUZWvI6hFrDx40+sITs7EEXnTmn8ZoR5ZYeAf0tw/jo7sk8/VBuZ
7Iv0DWueRxG0Ur/MF6mzcWd4Jj7TjQ+Mz74NOBF5PMtmKqMtFznK53esU4oD9+GM
dHB1K/wv3o6BV6bByC14qupwMNItlgEnVkBWilV0x08eONoNOcxT4SKLGFnQwJ8j
j+p6AdOFCnhqTOM6SvefvSLDQkv7OKz5MdgN3mDJrJfK0mSwKMXB2oDdtPKLmsuG
7cCBqmca8W1OPcj/qQ0BUM4Gg2zoIybv5Qa1QRleNwaX4rF37+xp0J5Ddon6PBXz
CHbzcJFF2t7m5dzQEM9W1/eYd7Bus6QrUDbwJtgXAOYrmY+jBM/HMGchmC/LOeo9
DMk3AkxNHT4i+eYAnz/m3Ew2o826J0P9qdgB0PYw2gIqhFACL3VSszDvGAhxygb1
wHPiG43422TmYyVG2iNsMZ7lMQYUOXgBpSheWRsiCD/9PcsXgj4p6sudRKfMlV9N
5RboboVmFCPtg2HhosH+Y0G811VB+dcU1ltfajKlSVPQavUJ3R+/YOWPWyZv3kL9
QG6a3ojZ7H8S0rgJ0Mbr8Y+gFcJQqeBvYbxBfFSfon8TSQI7bP9pSy9xI2KBNI4p
GGyXCVptCSlrMkIBMFtILdCIKcMc3J+tQ9Qhkf+5L8qV9sPk3XmAJttlwRoHbuUp
7W2np2s8APg4IHW+d870h4Rgrut50gSoAk1cTcGJgKKHRvPJrDKvLMsPyFceynMa
+VGNiaw3qSoO3nrmnvCzlSInzOvMRIHctsQ6GqSs8WFXokTnq6iZ0iF8uYfGQ1fW
54EQGYAj0VMaUleAqwPum67PWxwufds8ilqhTKDpvZIKrKfISLWpOpslHB8VPnLW
zrO+ADygOTD78WQxC/INpkoxCoDk8ZUCc0Mu139ynDag0zT0Tzd+sFSs/9UkZogk
Yx2KqwgL33hV7DVtiKzb+m4cLrinsU/Z/GVBD/C4d5xKKGErmcYyhaX2PMN77cO/
YFVLplrR5RxNc7mTxwNPVbdypyGkhxj5LrGPmSLqwuNVN9nNBDlnbX5orraGODoc
Dq5cMxYIBAg0kjP3RJFyfSWUgafelf/QYS4g0PgVffdxkqQQc1f8ZHHX/YQJlOSj
2E8ulkdCMit/T3pljD+wwpnJgbywR2adSKj1DnNeCC3+5YhCknU9JgxPHWQu/CG8
Z7zRCfpWZ0jVr4qlVKi1zzEAdwzbWv3mfvr0JeSdmqvjaXJSrD3YfZpNM2sgb58g
S4bxglsuni4i45WVAs+qFeasAgMFEhr2impwk+Fps1rnPCOeuR+YCmUfNe4Q2c8y
0InqnmcC5x3vCsXbr3widpqMF2EnbMkGRN6fdt7hjtkd1ycql2hFKOSLS6behhF4
eT7Gb4jyZn4ixpTz64e6IThTWa9axPNbCmoGOQIMdhwzptB0QhVOnKtuC4+ZHt2k
TjkGmqpJt4PDNGiic08rtzSy63rLSutMFeiNtVXs+KE2lYEu0ix4uQGjhtGxzYg7
b6/N/xy+VBoOGNxDrUMlzpJDHXioybpHFt8WjBUktguxICWN5odJOrlLbSdVK5od
vh1TJF0raMSoeIKVNtcmM3cMiweweL1gCD39EBZC3uhEzqeNsuRfXGOT4upN4U3Q
pb6vA9xZxFO4uNvzxm6tJ2N94L5x4O6jOVu5RKdLaIlZnM96pNkvY+kyA1Y+A/Rl
SW+eF9XTkCHkZYaL406Ja01US7BOcSqjrwC3Iz4Zf7de1WesULnPwl3sf/AmjZlm
+fCv7zi9KhXw/Th/wxeImIqTDm+7RpSGjsMpfTruKBDPrDhkRoIC0uLwDrqaNTrv
6RobR6PvERX1h9SYyiW4EfkTulFhiR42x8pNDBtRXMRxtaCqaL6tfRfgm+krBQrE
7YJ6le/WL3bqB5NE8Uqci9U1ggIMVGocAkZXhS1ZMpbymItj/qtuHAFd/7FpLGmq
19quAiYNslAuvKqMfj8clSsiFMxSc09PbDlKu1ysGAjjVX5olD6+E8MnLKfAME88
64e7+pFOgzw9Zr3GWxkfAZoG0eM5PfG/OUEuZTbREEfiY8o8FObbrs9pMtDPCK9G
SlHJGzCi3a74V5CBh7MqfMvzFH+Pr8E9MkyxPETcrty4DHlrUbT0jWFkMmOV+76t
49ja3S1KjD7oShtjjVY+d0ZK4T7XS4awfowGeia2AxULdi8Oh05OdHlINJZFxz/i
qhUU7EnBVTpXXnekecoCiaVt9bfscyLwOqIdupQh4gLh2TOSzwB8e9gYQtGwZiiz
hgwKYqVMd568eKUSFAS+beXFrYiI33FRyUdp0wQyPFaJKd+0iwN1mU2FoN7unP1I
I40cLkKQ4kIaIp2bcbrpmpb1lvnKDTdQFJg5heOO/b6wUuSSXHRKyj2c9nk/lCK5
URBpfy5nzzGQw4ZfhXgLLO++/YwxmJDzz8mLBXRZnwkqpJrGTCcplO/JQIQB2Lln
9mUpsSzQEvzsC/5t0jkWxhqZj9u+DHVgRwd63GV1F0Ri5aChA4Tjnf4zne161EeR
PE6BmmdkHdKCfWE9cLUQV3cMPHvH5uEHVc5HDPVFPn15sbi7syiiwke7r1IcTmJz
ijiGl3rXXxqL6my/cdEWnjS3nrvc0QilnNuLLWVPL0Qqw6M7IvfnENsBAjQPUSPv
YoYEntHqheNrmNdFXO5uUxElvrNyw5LEm+EjMB5IicAIEZAG0gS7tSSe0CZ6pPAv
Z/lbcPdC+ZJ5HzVVOxmXx0tn2vgYnWh0YXb2dRVl2HfcFyvHzx4oiJHi1FxBEB4C
3TqukWQ1Ry5Tv2G+PtS2nB06h0F1HmLuHofLHMQHeBEJv4mPAxMisvFU/PVbHEss
dDXXfM2Sj8BUXjQRAxAdP/wz/38k3RjFtw87wZ0fVmg8+sojgXNXIJM4QXr/9bhU
ctmdvpG5VGkYSOpk+Jw/ld3kKCn8AGGR3pT5CHuGpyaXpWIAgCgbwyI4Do1okJWo
hj7CnXlbDTTLnM9rt/rOarKXE+1uhCt3RLLy/TpL9MOmLnu7hiPz3SQtY5jk+OYi
YxeuZKF4wm7s9aZsJ4JjkYvnI6Yr3+pt7hzMczbzOWIvyBjVNEn6ornZswsJKAb0
YBq8JnKB0e3GDx68yDSWt/AUp/FIgttN6o/DqWFefuZFM40jTJxDfZKjY5j28EyK
pfnO9Ab8xrZbv3qc2evhRn1WCF54cFMSHPr5xX6yd5bfWisX4PBlzntB8NGplQg3
msNEI/qjRMKVmHOM/8CykmG1ZA5aziZ/LE4Xp99TV2c3QN30qsitcRi9VqIxWVVp
uomW6rNCZGTTo7NqvZyAawWEXMl9/2Fdrof6AsJFgnkerEvvx/HXjxxUpuSIa2f4
qIQ62ynR9xTs+A5+kNG9tMb3ahF9+U5pvTJ8lkjY+5WQcGmIx4mq8BpO7wy3YruB
q2mEmTAM17oSgXtUXoCNuU55RBwLsZ2f4EE1zdQbYCtXawlLC+s4Zdar0FeqbQ98
FVqJFwsCdGVWQDxYKExmtmfHmMqNRYaWEi3oAsy+2bUjwcV710C/o32lepDz8vpf
s8sIdV4xMiKHb76iDfL0CWLtW18gJEL3UOoGQfylgMXSGTQ7uL1xrLrpYe6oi1vu
8UAuDoHp+dvV6jsslBEhWbVmoN2eoPxlSHVXWK4muXQmiU8IuMzjTV+r3YaJamqV
NsDQkLQ54ZgcuUG0wTdLEkGwu5hn3AN+lA6I7U1ykkbSJyHhG8Xyu23oWilFcfZX
wS8hx1TEQtt2cuaglaQqQUYEFfTmlFWjE3RQ5Y1YmHksWz2W04BqKBuHkfPLt3dk
roORGvh8QjGsCiXigPLc8j1KGN9Iw0Xj6Pme9oxCe0fJGDDPI7COjUwhUnUMWpFp
wXYnQLA09TJ/kCJTOKQP8GhW0bTFDpeYAjXtPI+SU9wCqL8N1waVuESSLRPM1GNu
nr3UG+lIzBUhBhXglTZ3rKp27gMh+N4qEwkjlOASiPbSvUG2oql4F20tpEzHT58p
mjpAN3wHwjZeQKDNfBVtfEwdVVBrkWJRWJ+eWMpArOAPPJ7uC//XDJjtBZd+r0OE
/hlNv7yGluoQLhyuIIHN9g3W4lVaCI6X0UrtZXblYKavhFBMLZ2JegV9Iv3nAD9E
1u/inprSIxjrKCk3y76sQQAWWT/AyIRGFWJG9FlOge7YjmIQHkuVEf8hwvRaLF2X
flR896G9BiE3U+IdNMiwIm7FufLSoTh5FMhm99fKZHvymOgtnK4FjP4tTNi+uLpq
wXds2vMJdeyVu25/1tOsAgAK3hZx3S/kr35b09hzJG4na3gLR7mrfUkgpRrmNQeF
zYMGwOfXrybT3wjEzKUmQGDV+nv4AvHyluBGdvu2SNRUBB8W7uRZpxfUyotNnUz5
8ls39y21OaZUo0HBhfJ3CLdHSYQiA1DL/6jwpYIWcSbtzLDoOY669WnB61wgq3TG
saSpWyAybpmODkmSh1G/whgaMxPNM4pVCry7brjdbC45hXmqhM7pz81wU7mEA8TD
E0XNBMUAgrT1jmuIzbSDCq2vB1bGAIBOAvT7s/+0csbSufJOHUP4NtlvHRXaRC/G
IaUQQDNlJyCXqBxuQeffdfw8XGZU23H6UoFmu2/khcTO2VjtmJ+Y11mDDkwINWTA
vdkFGFeImpS/kAyooFx3z04aWp/peZ+xZz+pZjexW3OAylnpRDwfMHopnOf2gwqA
6rP6VT7FHSc+2WL1ElCdH90P66cdOrXqbBYMhsDcofNQoLAjA/lrlJGhl+2el9mM
RTPPZA7ilhV0COwe7mszDPvuuCpVuGxsq5rUBegHgt4LFZCj8MCynhv7Jw5i4mEP
RWlZwdoB+mxoNnwYpVP26Ck8Lz8TQdnUmWoC/SbZZChmUKOUEoLjye9F3SElyQwc
FD0L95Uz2KB7sLZq/UAZwBm5CltZfTiGadOhqekkIYcdwJuE3JXYm8JPXBlHMpnT
wB11YLrJKxMmAhr+q1O3K53LinmSiKi0r0JsF2DHEwn7LPSrL3fPXnAX2A/lX0rP
CzZmZCvk5h4FLbsus4S6YEMu8hA757UdMGfM9TXaeTXGDJ+buoIYQmCg4ovOa/iX
+XwNS71aAj0UMivvXDMlEh4oQX7+8+69I1I0ctRQokz5ye/6pSa+yrRYl8dYeWkP
e59qHp+zGCidYkupNJbD6SdKeB9uZrdon1ROSeI3xV9l/U1PPzQVuXcpZz3RGO+p
53diYt1grT2etb2aGNc9xO8pp6Wk7k8GF4QlAAFMODFdCgsNMbbL17/sadohDkur
2xYGQ/BoPOYDlXjxxNO6DHtzmPnctlhYgJuV0xUB7j9aweKjTVRhuDbHir5QGMTs
XQ38+h32pE9DOcFPvnZb2+pZrboKPOnjkqDRvdohxwDP2PaNuspTn3YVwyDOXrKP
xxUsZtGktt/iR1UTgsujbquBL+258xigGnlOct6iKn1PuArIJC+IABfA6Gw+W5wc
9O+5cdInt9D/PntpIbGO5KWEK8RGPU0J91JUYPqB+yX2QRySGF6JwTABYWH/QJN8
rHaKSxbhfnlf99WLEHrR+Gwm1oHonmbzQMZHI1XzNIkoAdm6aIhcV+gZtbArob/J
eUB/pCdMkhI4D7nQlsHVehmghw140ITyvB82UsrMaTFbfuV7xctBs+zYvizm4hNh
26HXOG8RCCWwg0OfVvs/zcwiv7q2Z907xsV27dA/gw7XT5D66SKf4+fK8Axs1GEX
zplHebck2DaKKSvYG2EdhZ60oZhM0HBYmxnC2LUM4IKnKofy+wojirmbHyiV8c03
dN8cPssktmPWLPiEqy/rumbBLC2jrB3fbI67dwqlMff+gVe6W9EUpB54W1WCG1rv
2bXa9QFI+fOsq8CsQpp5UMc6DBkdwT+Lu3KyXJfEQml2tSwIgG0Mb6mA6KwdAnWu
IQkQ1yakkr0mx1der+Bz2/SdQVAVnOBDQGY4SicptQAf4PDN7FO4n2VLXDqnCWQ1
p1YW0YP1vD3FJlpPkvNOy+rsbxAXZOmiRIvlutxPqKmDiAorArRi0jaFcZ9W2IcA
mdKRgOx2WIVDenq5EjhslXAjtsjdmIFe3PGpCIRHu87lpa0LJC4a7szyHnEGBjo9
xPFbgQM3iIdvddWCPzbnmsk0LC8XUnBqSe4O6wIduAxq44n3bteB/6QRB+Ot2UuZ
9rSSgKLyBTdKtPaG3mdeOynFOL03k1hiQ+R+WBZXgonDINlflNgBtfT0a8SSJ4sj
oXk59AiAGDQhGBExKs6D65whxj2IjeMqdNNSpXKEekIx7o2V4Lk0CiF28GcitDHQ
w7eILmBULcRtatwgjGJJmlDKT9ClOJh+O2KJ+YaAPoF5yCT8w4vaGMN8s/Srxc5U
Gu+h1A9VI9VOqTv0YR7CsNbfbwwwF3jy+azCD/urPVNJeHHZw1BobCMG2xGr5NXa
Dp+lYQuQBhoQ0WAnAZv9OM4LOFtUA+l+NcS0WJA6au4IIojnbFKFLpNWb7EC7aYw
Bb+Xltmh6SXwJqFFJycWbAKZov6MoG8gxY68MS1/Oa4jMiKjjiRqbGAunbJgOcle
PIyozON8KhTdewdBEgBHvfMM7mMpcKrtDlvGyHmpMNScNv3agBrTpxv/FxzZ7Ggx
il6VIn83/ZnbP1UFIjcECMcEiqBJUjuKB8XyeiyylOvKVsLGa9kE5WCtInVG1jvs
6SCeRSsTBepyM3qbPg9CMxRzqI6lnTkYkbXT/JjpftV51MKCjWyjeROBR62prfr9
OW7nxo6GVYcGF0Aud91UXzWzAkMGmuBMclFmV3eIrxJmJKLBELy852/77A8yMSmA
6P6z6cA6q+flfpikUklAtbNcSngkexbGZv1l8WlLtEciIUXgnBYkbZWlaqt+WEU8
IJuCJn8Tp37EtH9D4AoGrP8QqcD4nctPmLYdReQw7JWPeDAcHKqh4Gu2FUSsSV0k
9ZTy7w+bQ6A4vUCyYIxQN1XFCGsXuujlYyWAXWxh8fAmvsavvxl6JkRDaLWJgQ8l
JQonISUmG02uMVMQLFa+BEx1DPiX9x7//um2W472VjYGIUAgsQ83WT96SZ6tUhKp
/nqF2zpGecZHWUhBq0JagVuTJKjRyYjVqWEGZs4HgWm+5geCNpSuuityKOkZT9MA
BXZkgopB+F0gUeW5KJxokVBJf45kgRz7LjMJvw6UJRnAV4LDiWeKivKYY1MdXcqA
ZTWb0FAADyCjKcsPfNvwMJJA5QSMFWNInl/G0VcXul3/JgRZSf26XjdElUxN3Vb7
JfS6A3pUPKEPmdBCEmfMM4pcWsM1EYdw//d4SGB9pOpmd8G4sDkg7Uj8brjYgFXd
OejfA2SiT1wDAfNnhJAk7QGw8gcdyZaA5OCKgqgsuZ2my/mryeD/0XzMQsMUbxrB
4IcpbkQzRDhp1FRJ2RmPvux9CVuiwwOFtdEBn5PlSxPZRkYFm0+eN1BUEXxaKYAY
SWur2le8s8yiNlBOuk3jKuPC2QAi1lwZZFusaDAT/BT83cSSXtkuCgw4BrmpJaX3
MTJIEouXr/jCWwe8Yq22zjzC4pgfJxZoI35fUtdQN2wU05X+X0SihMP7RCCgomyZ
litQx09XxuEgSOl2EpXaPFUHzpoiiyzV6iYNT92zKM9P8KmASvILBZ1MiLkkf2uK
TczegMM+iHcwA2ECCD+QqlGTeUsJ6qPWMBClpid7wBWD0cpcutaNMoc2T6DrTUyi
mDfcMw2TGKz6DuSNbH+SHi+d6wGSPcW0hfGIUZnsiJQHZdcfTDZmVmOwgHyiu7qY
O/lfMwSE39uv/p/9zNyuk3LrLnBesvWNjmyhYjp2zdtBnM75ZvvD9MLavDhD4RFR
/EixYk2boC4GC+K/izyEENZuVeJphuei1HQ0zH27KBr/WSrmn1Wh8fT0bVdeFSxr
nSIFrL8p25hQwwnZ9mnSnLYQJUpm3mGyC6jRGh+j+9xFav+nlKi8jOKAFD/Ro171
lQ6sKdcUoo9DDA7qdhMlvGDIeA6Hc9c2Q9+/XikpkQHNrdBtqbvzuAPp4EzbAunr
/cp+5hADQqJQIYqKoSGPJ0jc6Iu6GTjqH1YZfVtOaRcoNiJgEojF89upENlm/5IY
jHVfOCD72UmhKFDyHe2ZJzT8HFbUQow8Ub/uMoe1KMV9jnvwcp2NU9cH23GblZyC
qW3hrRAyNI8IeJ+8yBNUFJXzXUC822SrYVT3OKuSXt2N5KFT0ghZgQU2/XPZkrRe
PEjYd6L556EuEuU9TfP26j/Ax7+kdRwkI5X1chMOmmOo9Yz/diXBotL8Y0PpMs9j
hqJ+B8UhYU7Q2X+xb8LBeAWFiVzcieWJ5Hl4FEE8xrMiomuv2EzpsUTBp7qBOY2J
vrX53iyQMjifLiY4d51+jYPyXPUTMd0PlT1IlJKz/iSyJO3JgcJwxUE5/vULXrxc
7sAoe4YBfXKO/IhhcpE3lgwqyOE4+yNn/EGU6xHm91PS9cOjBR7YzNjKRTzNR/8m
8j/3b1U+g4N9UndW4a9OLxjafcabykfHhNyzPV3GewSJ68MvVAWtbOxVcJYRHKr1
cQCKDnIXIkSSMS7zRDMsPTW6Hh/0dx8JA51Bsj9tOWFC4Q5pchMx0yedmfvZcw+l
25CV4xWEG8pKQ+L85HkiRrGdzZ0KbSTAD7IRzg5f0wNZzOtB1UkAXzK1yaEo8V/t
yctHQfpvPVuiszGyFrnN+WRYeaJewrXIg4Bf+zlrW/Fsq8DzkYzmdhWDLxrrLtc4
Sze7Vtwh18U6zh+Kagwx+TGgLwg4eB3p3jveyZDPMrxh/wS+oOwcJ9lhyUIzcI59
TqnwqKgxX3Q1vSHkLGuo++XvAIjB8Utx3VBL29lrCEYt8mlWIzDJ8UUm6Y55gC55
OimaQtoGnKbfCJzn3GQNI3p2ixepvcfKIA+hmLqoA3aFELTrbzU4XqttL1zsDopD
7vm1jz4g+2ItpqeAUzTw5HiFSswCKtkmxFnkDVCGAIyrZWssdMHgR1bESfVJTVn4
5FWzlxzX2DfCnNhvcgNiZ2XM2XPNfLqROrplXSMt3MBFlnQ1h7ZZs/eTY4sB7kvV
ZdEwlVkKb5TXY1EjLeyLprFGtOPdY5/h8fIXHV1hiB/CwsYM6Yxa4XA+F11d/2pq
j1NL2elypCKDYmkuuIxtEhWCQsDE+rFlS9FqvlBQnnZMJ0T7Se3X4EjG0t6zqbOK
5is4Nz5QZG2a40h7XZhwMgyk+wxJ7VmnhRGbikkEKSRkz46jDC3I+8/IV6yIF5N3
WYHCsU1oFvvNHGH2tqLVnPaRYjaXFkSAfOsns2XxdjFcNWlvPcnPXQVxDaH7CqJL
KCdVsMzeVvop5cn6P1KTq0v4nV0Ij0L9BO5PXpVTUj8uzJhzmGR4u4nMyVfgMrCS
k7A4bNiRcNYidLbvWgfBHOjv2oU5AswPh6XGs0WdwEupKfnvr6pLEXyWm8z55HQF
A/nvRGF+oHzFBBcVQQmcAHth4cyoNE5fXNVk1O7CQYioytnw9JBW1PpySZBHrShd
Hhawzuj9V80LqcryIY0b9Ukk8es+L2eP8YZWWwsJ1VQnn+zwkphW1pt9uHYkcRnX
JavQYA1u8U4A44x/UAOkWmLUWRam+3pCHNWgaPAH0L2xA5NrARe0Hl8WPOpV7NF2
P67LR+N5eR6hXQGXN3/AXJg+QskCMX42HJTPaFfhWc8qQHX7H5zIj9dhXnhToXXb
pyqGRsJxQjbGxEvWaANXnoBq46JGOVU6jqWVHq1mQ456W563bahKxV1tlIdcG9B6
4soJ0L93R8aVVurZ6Ny4BElljfL9YBUkaBwvZnvmMkjk09HSb1Jc1Sdi9Vae/GSV
Buw+VqFKjLl4Ku7vJYhWRckmpqTpFXQ1PQqc/Ul7daHmFsxLtRt4v1SgGrnm/8Qh
qYH2EyWVpkNfpDOubTz1YRhm5La9yOKMAounnBS5c12QOQZvGAigksk/UsdrVG0C
n4sxus6w+Jmp5QqVMxwLNTWwmxpeqN1gtXHfJWHUlGTrN1bw1otULmmlD/TlduIg
T1IqcKtmA0307+B5NbS+qjWY5C6Xhi0ixow62SMI/WY/nccmVD+ciP52uT+XdBCl
D4Dyzjsk+6lqoTxn+7XMv4m7qMK346Tmzud+roEriaQNHxOHKko/4M/XzEwuDEy+
9n0OFt2HU4ODlF+Vup+SvajEhjxq52WZzi1VkV9UZIH4Es1QrXet853zGmit1Icj
QYykKwTnf9tkaohMeFSmOSNQ0QJyTpDIbNLPTweawMax/PaXUlnEWjcHm6T4UF1L
r/3faomQsNcW5n1bzSmYFAisZfhvGK4/S6KGBNTBbEDD6JWyZRdE7xQ0ZqaPTKj6
b3xOagd2zGMtiCmuOzniU28e0+IExMXmz8CADHChCxwON6CXuDM1EXrmUFz3tov+
FvPmGaFywTJdL5dU+R2iAejBGN9+P6VvPWPxvBrTTdXufXlSkXwTl9foIjngVMw/
1xHrMIhXzXK9wnDGk5zobkGpsehIddHnUeUJ3tSa/6wmB9hrEseCBUk8a+4UFiLw
AwX0Fy6bmLMskp7UV5O2MmBrieU+JwwYbiyQ/Wz61YplOuGUVYwkYUwbVFvP0YtJ
kyAyQ2NMtWUwv1LXg2/JNZ2J3X/O+4vx448N2A5o0MR6oxlOp5zxQg8YQW2f8A9M
VUCH1PZSzXhuGTfJVtHxN9gpAJCG8ZY7fx0hbQHr2+qYPrfu1iFdr8jizmv+2xT9
kqGTSdDlykoBne9d6rXtMrPMv7BtfzS+2j7p5u0LNNR7Bg9Ct9LGC+MCnfJBZThN
IQjBq4F1MkXKVxYfHzd6/PmalpXHPxHv+HQOOsPda+hAIOvuFJpbFL2sLXHVUazI
HpIS/R78nLhEG/6tfVdl1i5tt96OQ752afbIUMlu+dhTfdLUL+jsLM1dW5SHL3TM
cDhSgr0NRgpoak7KXfz7JQOqnpXVVkiXQhd6TdUmc7m/dgKN5APijjji8lMtrBk9
/thcUMTnO/+FN2JkbPAdPTkPKcCA7ko+lx4p6/3WezOE8p0KUQG4gT2yL8r2buWm
+RcvcyL8DwxO8DUo4F2jK7EOr99EMotSvtATk614SGreeOHoXkea33Co8XCiLm50
aUlNFY15n+TsC6IAgFXb6mI/l+GR3OwHqlobdJjs+ZZixjp0+Zrhh8gmBbwdGPl3
cHWNaxg5LL7zpK+9M60B+rSculf+kwdHGrsitQHr1sVcWKuu1GBBlwqU9O1gt7qF
scS5T2godWOIHFiFJqto0WugkKC1JEhcm+Fy94DMlsKIkD6rTEwqEydwsLL1hGwc
ee2baKwk8ubrHN3FmXu5zQHupaBqaNMPkMkzuRvK8GBelKUoMq6RpMnmEQOhB2mv
mES7LVW5u+FfVGVO+DLo1l/JQ6RDNp/I1XQZdw6adHB1zH7omYmxVtZ1mTGTh6xP
z6hCiV3NuFTqcebK2rumMiyuYlVIFDWvf5a5bh7TdEBfRTJCSARxTwCfAVFRIy4K
62kil3/hHpzTpexOnjyNgQDpbaxJXk7T3fvQx8ZjDcgiE9RHEVWzD5ZL0x3iDn7N
1Il3Ruj4be13wqMy6Zxi7v/WWYrEoOmDnh6dMg7YPjkCB6jx8o0fcNkE2H+btSvL
vFTjlHcxwzDHkSoz6yg8g5QgXZMOYxixba8kEDpYAbi2ijCChhmceHZfWYO3tdEg
lXJuKDAut0rUi3o1pA7f40L4CCfHYKBVzZ4KH51sPuoXtKg9WjFy9aQAV0jowbGE
4lxHCWn9FwBVtwWIf9WvkG9wyUs++A2Safn8iBHzH+dUQz2OIhESHIkG884yEWvH
OcuaW3aAh6uPQk1pZBCUdldrMWkYbHWyrg4IY74hDl8t8K5UQEoCIpEKm6x/ScME
ID9hHoPuhobJZP6jTCfeWunMYfYx2gIkpuiT2RlTp70hvpBuV+FwQ16eScYl48Dn
7pte+oIIG+zn7mS7aP+D1b7EPCP/foJHV584fPy+vb95s06rmsCzAdAizYNtto21
SONnvcZbfIZRWy8tlFnTvqxhb+luekvUFW+293PI5hveiyBXAQCNGcOC4UpyXkjR
PAsmgmRg/nmV59Ft5Ha/b6VOqhPBrsmyV0KVFXDgGUCCZWwmhsS7KiA1NybVWr2b
pGxRhD4cy/cNsXN/CEvMxJe1zN6Y5FSblxMFRRKM7dmTtkiL166oMGO7DAbiaei/
nVKe1YRBnzsO5w9rGaDul7/zBFZpeCUc+Xvo2FzRVg/DLd6ywusn/3uoWM5ahmBq
tQsdKSYeMVQPBNdsRnRU189EiV4rq0ymzkmEh1RgYLUqX9TRT1XUfECkEP45R1Qi
X2dp8nwD8es9y+nr3mUyw9D+SntgMbqnIqREKnrUqSmj91DLy9ZYb6jFJ8PLPS8B
VYnniZc6bBZ3gKdVb6+wHthrIlfh9RkEsExbEIymVpddL+VXcWMDTsqKYHapOuxB
YzxK5zjfeQsAGn3F7kg6oHxoauBEzlLNouFZgvAraEZxVIxBveyAYds3q+7KR7dG
eIgCoQAkxqy8IhwSzXmAEE8x0N/9arA8di8Qm8e2UC4dfB5pHyHD6YiUH9jEKzYw
rfE5a+iMeVxZzk/acJQQ8Xt1/EiEfDQhWRQI8sNYwJzJBCkxvwM6lejWPzGVWdBy
swO60hzYAZHXRwOqH5pp0FKyaj6+5zb1iIyzxdp+4M2buM23ECMXVkdvh5ZR+xfl
79hx/+9kOK+s0MG0fSrF42PWNumpE5cw8XQqJLNw4WJvpDKiS/J8ZD+9BeiNUN7K
02Vi044RdkRE65uj18Jfu4ReIo3I0CnlA7bE1N7kfOgBYYygim0ZIj8hl6IG1dIB
y4uJbDvYu9GTJsK8OEH02IEZL51v5+GxzV29OMC2h7kmE6J4cqb8L3ah6AsL6hHd
wyoDKlsP1Q5x6RSEZy7q/depO235Mar2lec98HaO/o4jQSWY+nP+4nemRmKom2w5
AHTziGB4mFi+fLbESHWDY7iUbKXxCt2AWs8GPSGy3yfY01aSsjU9B5IwDxyzhuUf
qiJeuUhaFFSab/Ad1BkWxWc8snne3T8vTrMTMCwWXsaHPU6x5htieAdHbnqzwsDQ
KDhitZhAL2p7HvPEdNVdOa2tx3Z/OYvCStnPbgj7MpDYaSICnVaqOSaMdXRxuPG4
KAFeR6uApd7cgnUWNo6XRooSr/mZGg/q27mU10wEblSSB7zpWKq5i9+11qTMkzXd
NW095Q6eAOTX4+uuTBmhP9GaluYUphK+kgGViUt+/xTJA/++LdHfHbHifDUUnS5O
BdkpebvtweCjvgxPRqxz9rLr2UHMyBGJsDqw5UoJERZhLpDmJZreLypSuqaTeuv2
vd/cfv3evcxfJMxI/ZiG/5a2LY+tzKYh1pfmvIAJXOO/menL7j2gq34+8q1PghHa
z148/gG2IpBB7SZ7IvPJqYPQxZcfNV9956hPxPDdCzMoDX4EqB7YB5CfEAneTOih
gRZBMvr9QiUhFY6SmPIT4h98sxMTfa78Xs6cgIXUedPhsAzyBBrGXKCRlFDaB8AF
gHysJQI+ujffBk6xGnGV1GpItTm+sNyUjtx2F9Sf5lZSA9xMH5cl3vB1fUHcnfC4
KZ96rXTdVKw0TVaKJ+x3yRFOdd1SXGUmHi8lv1WB5DptI3IDiZkrY055/zcxkQ8k
rgEV57ZcSsboU9oj9Rzwca1iniEt1no/9yGDeUgZY36tzuyNenpr4m7HWUNKzfAU
3QxfW4xI/+h7f27H0zmBYrfr6+dxepvSXJdu3xgbB5tEOY2rTa44qxQOo0CanURe
aB6vkm56aqogiDoNV2Ta17v64CxUU4KlKtrwEzsPIRTqenpKV7i8cPRfkONj3OfO
3oDDgqr2rgspcHjAEJ8XEEjFuy8zeEyVLB7OmIiR9C5PRz4lajSaZozFdNECdW0a
3fPglenaeOwzS+d81SoHUCfdGGTL1fsOlNwsnBNHrBNfVS576owqFrjdf9RAnNV4
lRXwa6Ft/NuXbJgCrqF9kpcP+WSEb1uIuRXItLAbivNK6vxenpxUaeMMrPkWa1c7
yKzPWb50PMcpjkpzwU9z+Ucjx11WpQx4bmJQwgH2SAas9WvDSTtp0Cl0FKNLcNaX
zh7Lz7pNAIPqS1bbg/z9+QvascaELweJEi2Cz+tX4vtUJgwYz02qoqsico7IqkMO
B7C7lAV7JBjvMCXhDudszFe4LEifWWm9x9e1EgYUI58Y9c2Asp+JO7XCvHd8myRP
R5NbrCL6cmZMnY2fhu6NUrk3N+JpJu6WWQqcFnuzFdcDDF5s2Bh5Ujwh/7H1ehaO
LnHVCDX1JN3n/TSyRVDh1jyJAoip4QBD2RVzoXbySzeVVAifO/ZrTHxpc5FWVgNl
iUe+4ZGzxBeT7vBwGhGhW/vYITXNlVgyV+OInrFeoNhIggb65z+De1mY+WVClDKM
Vt/ug3sd75R1l85saM/njQKy1RK3NNr05MnodSANPyocMNGaCMCyVTQ/mn0X6VGk
zSD/Gu+Mj6X3kJIWOWnyXDLj797ewTs2fYeCzAHSqBHEeAcX94l3vjqcxFHtaZ43
LLBzQac5oT4gEmM9S7KEjOC13tnWSHZc3P8UmQTr/9L7Q53YRbxkf4YzKYYoV27M
QOAXz9jCOZ1VGysijVjZgUjA4uCOUKC5flMXvvZgTr7nvBW8GRL4Krx+m81yDM6R
71u+IxheGJ3m2pWtvuKGbVL6oAGJV/+/2psdq65L/NGlaPAvmPnSREmyj8MyI5yx
S3xi8XOBXsi+zCLetHZyA6JQmpgZ/I3/8O861y3gFXp60xPhc8JDuE9d5+wmDO+g
BihJZUWtchUpv0JmXzvR8hM3N8BPVphr8dcTEakc7x5TOGXvHPZSXl2S4JqyHgNu
EHMjDgQ2C0zGg+4v4hzMHeAOQf7zMurQsBE6o3W4HXmaLBFWwxz+pwZ/IaKGxMpR
JFKQUEOicP1fRiNjF79l96cpC/hATmEY/dhwNKNi/MMrfCzI3tHT0CIM2gDcTC3q
U0O1eKDEEMzyX2rog4rSNTsyWVA8cKr6hpn3TJf9FXTqq3gPtdJq0YFussm73MyF
DbUqPtwMaqJEJmgEe1sqsRGORvqlfOtrGmX/qt2mnJKFD8Ta1Gg12yp23iiB/E/Z
JFzrYBLQWYdxc1tQpQBWKUXAiXpC9P/S1pUgrc1wdd6Thx733uBFbxUXKdXI7TxP
gsp6M0cvi0jyXyUZBgYDtP9OBCuB6dc3ZTk2mQv5sWdSAinlY2Z7lKniniZRvzFo
TA5hPF6mr9ZmHKRTcEnz47D6pL7U+SH0trhCRWfugoGxYxrvUDmFoLPz/bMwhOVp
B+xgTLyQpg02PnXP2pTIbHcEiq9NmyU1u1aqOw8Hks6I4JcoBFLXsUdQPUjl/YYw
26Dduvq5ftC7rtPtPs/BQse8lrhA4tNA4j56KQQCasRLu79+HkgsgQibFhW4tZda
YJP5gu/EKCfXwHWcqMA06d9idcAsmyvVow9y1ICynBOJ0dyPCQ/q/ajBOZEgahOJ
eS5CMT3rN2TX2Z8P2T+iwo/4mhHUoOy6enPYK5i+wY0bmjrL6KMXOwxiGu5MsPI+
lOPacvVQ65qK/ljsusji2nu5C0e1LdEYyKZFnOSO5gjhCszIMqGSeamNqwB5XTIR
Vr9eSSDVAC4uhnFY/QjwJQqHQHNzNWLlPmaXU3uIELeTX2sRAdrgSv74B2RWwOhU
aJQglEswgC86cM1Qcjv4gJhQhAL1sMA7A1HmHdJPqSssdlJMwZJR/+25H10yesxM
OeujbYmlcKfi1+AtQ88oMF3foW6rUyv/eJttoDJpkuj51w6Kj8nENnu1ibMUTnEo
Uw46jsBP90OoDLv1OWbn8diQfoAee4V7V1FNm1l1jqWSoXZLsuMI3hIJKFUo1iFm
/V8wpwj4JS8dUvbK4AQhHNm3CdkkyhTbkNy/24yhfjxvVwn5IAoQeIeHPFO6v2oo
dDm+dtuPqUB6x/K+amqlFRgiaUW6LoxuTm7sxZ0mKLC0SKF67C1ZZmIcaniyIa4x
HdxGg80M7YTqAdPLgO35ceNE8IT05eJIYp+LawgGwlyaY0ZKWQY8v6oZMzl8e2OO
RYGXiB6wqL8p59qlA4mevNPZtCq/4d5nbhoWbBPXGt6KMdFI1L+2i1G5wFiEfizm
LlvOm6NuvxDTlwYc1uXxE6zr/J4QPUr1DozhJ9y3oTL+H6Ispv6mjg0Rw+ysAeQ7
Hjt7BXDjnHqQjCvTgVXbxpCLxzxlx9frFHLXdqb03qodHGJuajuMY+R03BsDCObt
yIoE11tB0G9ZPMKY3L0xy81gylNWRF6xQLnItYmWbE9hnf/8cnC+x8sCHlZAZgnS
A/yDZ0kPEBcPNvHBznki4jJUCH44TqU5V/Mr6S2G7hqwtt4OP/nqhEp2UFmA47aT
xtDWx+ooq5LtU1MbNCZCtzVhnQ97D2GJqfp8aqEj7PljGhvDuITy+jqFdUcnCdTe
vW3E+wtJ9zKuvKHvYwx6Y1oDUsMu/tLO8Mx1gXEXg2xHfpgB9avSTFowt7035gYa
Z8HT1EVhREKelyRK2x1q3lCEk3RjexIIzBCQXuRKyAzVXnl5Y8pfImbicZ/2XS/X
ahArgwK2DWZgJFjDkQovHbW4krIinkgxoXWhU8pN5J8Aoc2+U/SGsefF4ZXqdtJT
h3lb3rUa9PV+uiyp2d/yu1wJ9XSRPcOI2G4pAhy3GFKJwbMc/Juxs2pwCD1FzELk
l18UOdER7MuEfAFHXsYylOFmvu2U/yfo0najd/JMSi6SLxrXuq2zXsmDeHNvCnRb
R5bgpQvxmIflQMgpJjzQCXlhh1fw3OhY11/NPTk6QvWHPg0iEnMEAZxUcjQHAlPc
0sOKsrpXUhKWdIlLL4QJWrSkA5Z9OnXYPPz32RHKaX7UeEJn25X9dGRReDmIZFCS
0nI7HrDE3KXGEPAyB1l4lxHGd6iBk82eqzjhHtKrvY/Me/NBgZgoQqP96lHE2GTg
5viTW5A8CmIFOKnXZN6OST/bXRrNOeX0euuX4c9fm4cOceQDmoIKaV8Qdk4O+/nN
IuDevmPmLTVoNGNboWXy6lFVDExh+8LCGhLsIoXwOInAJNQXZ003/ZHKBmt907Ek
YuEmgL8I9VQe3InJ5b5lKv+7fMrpcuo/7eg0gG5b5sYvJb/hPbapna+pnePDEgsG
+YodYZzeFM/02olTiW1CafF0vB5wefmA0vAfm5DYFhpvRzqAa42ec0EqwpEUIem4
O35s6n2r532p2vrUc7TN5yyr5hEKPa9Z+xkgB5KOM1Pa4A5pyj+G+spVYnESe6Y1
/uwPtf/meF89baAssfumXUnQa8heZWgLHNWjAdE+W6Tb79GcL0n+bN186DAWzMha
ByVFns/R7jrScg2JBiPGvSV9oFxLc8gtoScAKu9oVydkiVeBQFNZZcskjcqfXheT
52bgmIvUNHRw7eJg9ONSJYecth6Hs0Q3WY3pamE7LyB6EfZ1ezVZ32r5m5mLam2S
Z/n1LfLPIwk3TIQQFctubQtm+LMjQ8KQOgSBMdBvf6ppCzy0MctWiS7iUjNhv7Pm
WjCQGywKKuPYgVxlZ5igdSltN+mNJjbcJb5AU7xQD3QIWb3oiycYzGe28s3HO8IR
iTXKjznJ6s6MhbdTW4AmZzAhFIcsQxzOzSDgr190fHNYGTiy+3eYAW4TAJwj+Fey
l0NYLfJZ8HGAfMp8dSXna+pWduMQkAHXql2obQCXXN6UKApAGvu9Ctx66aMImVxw
zFhGpgstvnVPUP9haA88ebv/YvG62GdqKRNt3ZfuZ/d881YXTvtsWJISf9Nn6D2y
vVXdOV261Cdo8TTnIh9enzWZ46uPQ2VHs2gKBJsOpeMtezwfQ8aNMmftQ/IHOOyd
g+/ayyksgtExrjZFv0iT2CmfiiotaujPcaR+/FL4LQCqpSXxaBK6Ge+aiC7UG/eu
LT/DMnVKHWhEBgItPDuZ/JXMcmGC4s9qKXF6VmNretbvc5M0428yA63sYSP8QZlG
eGCZ0kenh/j6NsmFcsMDBguABhpWUzc92n3WPOCX/tm3KdBPqb1mxnxfjHOsM+zq
bq4eSNAaP6GqhksfVpWsorsFIho9uVHuwRtfZQ/9q86x8Nu/Na9QK8Q3VF4OkAij
iohzAdSxaBLpn4ELfZxcRaXXU19Jj/KA5oMsW6MXX+3Hn/u1rEug0miuu00DwW7e
fGVEFN5X1zaNLkhcy+/MFwdOmdd71rzWw0uxfbK9R4bqEGPL5s+pQeXs+yhSKF8j
ROljFkdj2N5NuNDS+1dkhqLllBDzOgtStIJZYiBs8I9hOzyApxRoqHeZ65uBThf8
3e+YLD8aCnQ1G05Bgbsuf7DKPU5yvoMNOXCdFnF4QTDWbXpW5Lsq8adlXQcP3IsU
oweUsgTiRayE9BBujohAhix0Aoz/S6axbycFZf+ulowP2i3D4Y0pa96cE79+uB+t
Wai2tWlnauGuRryjjpyOxWF1ki01NIbzC8pZq8xOdXcUhfWaWatc1kkngBpoY3oS
fy2/LmUx5rYmeXk9ob23FaSff4JWWIGpJ384J9XQMtg61N8ceD7CocCgwrkpzD8J
WhFGrB5BM6Ceg7xGbTc42x7fwrDBvSMnA9+b2BKcF5Fiptg+BN+C9NOIW2DQNCM6
YBAG77yOku1e0yIe4R6pjg5kYRTmaHrr/VcP/q+H2+tX16N8GgfpYGaNDly6/EAA
vqtOiq73ELmwrp32EBWTqsD5ZxYuc3uzmBcsPhjQOm/o9+9jeM4ytppHj//ym1Ir
hLVviQ1eGRRfi2tqnuxzMB4nBFZOp0KNMZ0EJAhq2DIFlcIGidi+K8j6UYxWzxSj
YlFuxF0gTlFVrJEb+og3obOf6K4emgq58avfHc9z0iCC/OHIos2ONFEsyrLwXw2K
oa/XLmTVBuzeP9sWzTNSg7hdMNc+hmFBG6nhackBhZhAdwDJcgdGtNcyVP4fSMZb
M/zAa/DgJ8gkZTmVNTw2aESNKNEEDQQM2bxWy4tesT5S3itlsV3tsVlTToRjn7IY
RqeCY6r1KAZekQ16XSz9beYB8hDFhHvLtFtTQpI/QjVuCKFxY1B1oiuxkm4/iPHj
SA6NKsUTG9B07LCkVFouLw0gPj0aHlMjHgVhje7hOlhcRIBCgQaVwNepAcinc/Yg
gkq9ZymXpk6d+9k51om3J/jmvd3ru8oedERa+SN44+dcLLv8QEy+4iApHjbBJ3rT
tT7c7k92szflDYj7SdyK6sqC5d0KUsdfJzUvZzgKqvWBtsNs5XCkgO1de0vREq4S
cEOpwADlUMR9KpaCmfLYd27ePeohHadYVQm0y9Z7Kuq9cZhB4DNbDa8NxrDUlEbN
+VBHpAw72oK1cgkB+sg9UigUyFD12psGXePMIX4y3PETkolu0H9zp2B45D9ybF5V
RS7dJJKiy7rGH7XTS6Be4dNqMzwqhkwLkHV+C7iH8G4fiBGwmrrAntdYE2cJTuZK
07nTITUysfLebG+lHugVYSAvQwlkSoAphEsQhAdVUHO+jR8CnT4ljX8XxcH3Hm4R
KqxFymZPkLw8HlOBPqyDortUdkajRs0Rdi+bmVDUUflaEXDJzKB3lL8PWg9+mu2A
yLdDGfXgSpjcrlhOrRz4l/kBWtJB/3hhXTTRTizceyLLi0kSpIGHQO2usJx3FUkR
epR87HSgWSk0o4XA8scWBrlu+iWhJHmNlJgAY8q/rIDLipHdiK+G12ywAIqDidzN
HYLNaRemuP5J0uAwWO8TbTJ6Rk48XcqCFDlbwvmYA/50oi1GFvoHuoUH5g+dALQE
SpO4BR7IfoXQPgxEnqX27euymsLTLSm7/MgZYKOtX0c/ujaMuJw6PwbyYYmRlQ8g
AdPrN0wBXIwuUQAC/1jeJM12+gfa7gTa658Bn+bOZVXNqSr/M/NXUmsY4hf0CMNC
S0qVl9fVycLgvTlb5J6AToLWJxziaGN2Til5wyc/da8tSZtQjnWGc0AiP1Pcudp9
+mKHocc5SbUjUfGocRHMflxBcRqMiUUiqKTagjxlqPnSGfrIyLcpqsCcnz3FMWn0
8+FiPSyp9uYEBNDVudwuQhq4ilJrsWTDacOHxkm+sXS0oGUu/9NextoeLc6wwV8/
ENt0qqnwIiJVji8b436HFENIbnE5oKVavgCYZW1C/RYAexFDnr/nQU8jb3W2lFRy
jtjeeRBLCZRE0tUsB+rTTWV/4by9OjyUP/1O2RarffQoFHoz09PlLi6x0lenwpBy
Cy6vk/LbSemBM6qIWfplUAMQdtX/W8iziIaNLVXvWM4IxURMuFImENS5wVfoZqeY
LWz90o+JmFw9q42NgcRMxoaQjhLssymfgr0X7kfeyHF0sXLszmFSmSG+vcX/Qqyy
uykdnfvOxkREHGZqInzi98iEvjL9XoMSr0XmUoGa8GPj27pG0aVtFH2NYBx6XIvD
l+EYgkydFmvNp/m6g+8ObQAXVlazBMk6PpU5Qvd75nj9MvMiPKSdUFQyWfzmlOmz
88HIIqe6iC468H9mSZYpyWVhar2QFCrlkSOes2qsl9/DGgVj+bP5WUu4Upg7vbpj
RuUv9gVD5xzRMlyf0+Ua5VkB/Jo/tvsuTGUihLJ2FN+VfFZvSNTenGWeLpbSY7Tq
mL2kcqBwGswSyQ2ozS3GjdolL06whJ0fJ2Z2qeRDDMcHP/jtXu7MMnn3YuIYyelU
/TiaGxvZkbAhZNiHdd6waE7VZptwYColtiSKuOMcBy4rVYR6VNEmDu3mmp3/YJbd
U+YBAqwCvmoBQAEUwGosULpD38hpcZEFGHwqluXw9SgnlOaJO/9gSvACTEzvMHrX
HZc7uj9YxrGaNWaSA6ASzLPvC4OULe8M3XwrElwXBd6UVlENj0wbXP+3yMM9AISO
Avh5kEWJ/hp2mKkPxFpTTjsVTYPZqAp02FWtDAGXWKd0lO5MrEhdtjqReQrssPaR
51J4oKiOLO6ERtu5k6GqjGw7naC0xeaHulkCW60ULIKpfISt3QcFUomUHDpu1Uzu
/xEGeBcBUtD9Y04SZQG00mpRJCFM9bFB4bRZQhgwUvRo7n3y2wmddrxLZ7j0hAOc
uJqvg7QodAU2MNUBQhvVAV/26OnQkIkulQxKi1aEIr6wvlCCfwLAqnguPhN1Oo7b
2tZKbMkME5bNTUo9vnIqb9xyfsqCbEcDDS8r639LR2pq8mPd+BAuth/+wI5klG6e
qY8bPFqy6ONuAZ/kKWHeXn3mpYe5MDjGgVRB6uF9bUhRQOeZeCHZ0SAoSnDl8Jpi
+v2pNv19G7eKUnBOY5UHwxXFto28Ls61sAJRF+OWvDrrecwiRLdpaH5r8ZN52Y1N
74CcVR6m+/chhAjt7u+DXelhiWMxmLisDHaN7k143ce/9zdChigp8MUq/4gC2443
ixED+2YZnuymLMqeGAJ3TqleLc0VXsnTCaBSY5wyVg3yJK/0tXpHyFZaEhXGvYhD
blEZ9MtfzPW25YEZ1a3ZRZrbj4ZFNjjjvKyn0nFpR8WwZhJlkso2KTDLAXfAF/2H
awbwkwUcnt5mgPO+/FDpgOESkCgVmIe0vnZYuIsRgI0g8DADTKrj63ueHt/qRug5
APrZM3FAfoUj+FSagCo0AmgrkZr/1DAprQrz2/YcSVvitkO9AQNCjRurMaJtcnDV
aisvOO7lJO2TARzFVlM75tsybVtr9bjWMLO1Am7LbdIglZGrLFD/gSPvVZ0glxaf
tAY7m8X1DnTUg/iCr1+7q+QORkSHQFUwgapFH71w6os8eet4JmBnI74AU8BtrDSX
LJpmnD/iyUAFdp6J+WLopxYT8obgAE887KlFWUgYS6M6uckkcv1wrrVIOOSJqlpZ
SBZK6RmCf3EeRE/KFJjSSIIfXLO3cdFvMpIjh8yzUgFaP16o0G3+Fq+sgfdYvW2j
CPPGLQFyO8nnPEuDGVXThfN1ZtDWyfkmIRKm9TMr16jXEyn+RfNCicrNpQdEwyEa
dk0r2eVA2X3aXaodSDy4m6FPgcLtlS7wK1J++HrNeD2q2jVbGMbeP6PyQ9PMbQuv
QQuiBuaTryPzz897sHuSl5ys8bv3nOVdg9Kl4Ww1TavrRZWq69jir6rlABJfzu87
SBPy9ogv2JA+T4MD3/Rivdatlq5U7JCCAJD907rg5WXkHgHJf0a8o3ZvMnEVTDHW
rS0RYAzK3EL8hWQvVwl1OoCaKRq2U6biHXWf7q5Vs7isO0gyBIPGiR2Rw0rRaY7L
Fo4AMKq1JjsezRLCo3SwQJuKc3sJpVSVZ7o2SAW/sEtU8GJiIDNeDXbpJgi9c5aE
7rM4e0lbxx6UEp7pIdmJsxHxCPb/NUR7KR6eyoFt7t1Lt3C4pUDRVYCbzpt7te9U
wzJp6hURPyjIPTCo05BZd7mboOcsn4ebEmKUpKmn5VHSGwiEOHX1NhBVzeojf4OX
n8+E3vaCeluKdEiOtXammc1TxU6VXBgtFpiBd0ao1vxFPIdVOO0UbINkKNwewbIF
Aw0CA2JFboKwBIYxeJco+n683tKdYLElAaRzOzPMIS3JcL/ZdPlcZ5JIG7f1VrvA
WUiJK+BXOmzrc6up7qfsIfSJFjjRVzByAYf9yx+EL4VSCVvoO8b++SDNSRH0ayTP
luZHSgtjX9BPs0mQK9+5JZmTHgXDTAzBo0uzMPPyNIvvlAxx6UeuUqrU0XQeJvjJ
n9jkblYm1E4ALHDHcaKPe3rL+Y8obAuw+MCVytP6577iJlrEzOnVYlHALgYirLDi
aBYycAs1jMQfVXukNHOThosUMMj4azXnL/DYH/CiYTySl/g0XZRfhN+1ivkQ7SaJ
KMceKDgjSmz/Ic7FBwWos9dusLzXkTTuOpG9g8pRwI690Mgi5v8uICES/Zk8j8+A
Ry3wtP7qBznvqhAZ6yUOQBPM3kLUabUfoGkaE/8vJuBG3DGBOtKBKSe8uKd08CH6
b4o8U8Xf9j4QQAJGvprqA1bEgkdqtw4PVgXlMCrD9Jg8aKAuVZuD6ezdX22NhGru
nFOrzpQ2mPutPTaTmdckoIXaD8MFiL/v2ENUoTMHl9L+Qco0iwHmwry0eTMBRp4q
YElY0zkAvnlgrlgwH7GK2uh3s5th0jR2nsOIRslBtJnSwNKfWo6RyKY9KXC1o9KC
7sJmZXJ1HRfNATBIx6rubEanK2X5SOZzCu4UxWxsKSuJ5nlCY+K4Ep1dCKHTMQ3P
VaNOzHIxIDKro03re9USKiM14Dq4BVC4yE9mAhISdfPpuWeAGK0hpYoOB/sa2/lD
NYZYaMqYok0artdkFs4d/bgjFp3vi2buMhU8KY11vBy7q5kgSwkoZ01x2oN34zyB
bxXbYf2iIabAivt3dv9gu2q5SjaTfYoCeWAZv2F2jpUNKi5A/PlCcAxb6UMAMCJy
FexfNGxoOcDtwflP/kdjn1oMwMvpC+GMf0jDGOGlnmIZ4xj6JfwrTjA8UJxID3in
h3WwUZTkjgZzFmV4Wh+jQKNUZhcMHUBn7f3PteEHIsoqdtC1GusVosC4W8omWCuw
XsFYqxpcwwl5hjENxDw+nd2lrALo3eL47QNleTN1MgAbpfBCEzvegPugW5mxyNoS
B8KgtS6x0vBB4dLPfIxju25uyxl2DV7ClZ7R9yWNAGPGsi1JguiG9WBTsXvOL3gn
PNXoPee3fZLgEAcq6R6zqMi9j2iDKxjNrw1GJpIryXY+iu+kS3FnJvU5rwyQOedS
k8IvmNlUvcjIsrQfNVzqPGGkF97I1wXqOc9EccAH7TDOLwvIiisxDU6XAllt8KMz
+c+4nzjSH7davCNPnTWi/BHc01hBtEMKkvqpMGatxPwXHi9H880zG1p07QItuw9e
dCWkLsjBX/Efa92xHYsx2SPyzPyYtkzyCnMHQjUCJlwGyRttcHUnlKL4sLDYr8wE
O1QDD3xTAKvvis5wDxkDvf8Rkclf/98PdlS3t3xGB2oTD0t7HzxOrXI7Q+Z9bpG6
Q+uX6eX5MVzktk/g3RzuzZdMFTEYTBjzjQmJVR4bZc9m0m9U9MYCb//eVkh8P8uE
2syOaHjkE8au8ml62oCNpBuT1j5QcjDd7WTXV8dwuUVIqDGMv+Y0XLEJIdj9ZxxN
bOEwgRoCVsnRVq9MnLZP5CChZRFs+vqhN+ro9hFi+Ck0D/0HMo8GlQYyjBR/KTK1
zZNATq71IOwcnw0/UGOU/WZQ+kQWzUApLN+qLh34exT+J3IM0ZJGDpHYwy8A9GUs
Gkq93CeRxFAqRrnoX1FHH3b2K45l7J/1vmixVKGPozfQ9Z63wynfg3M6ZK+tA6HA
kt0orOzBo+VyLkB6cEi+754gw5dTrJvBpiC9xtu8yfS6qKfSoy2YJukD2jbPlTT0
czredW7bmq3L9W9RooXDKqHL5wFymPW95f1uiMrNmiuAtKSqb/SWIfHorjG5B1o3
sfLvbdZtrfEGsIDzE0nwj2pZ9aBbSCjPOhJg2qTE5UwmVJ8090QO7xibYnaaydlP
FTCTtahUOLc/M9gXRnFONmP1N/YFcNGdpm6NvT0fqgdiMvH0DfKEbqC8WFWRRh3Y
CnEdv+dLVtfJfK5zsGyRcNxVT4GkFkzkoVgV9W8gKAAPa3nieScD8XTlT4ZPiYXq
Yaz0nIkCGuuHHbBej1FfyD9FCqEJnxVkTas5Fdja8F1nf3D1UThk23LEWob2qn2y
OdYlTTtCmbJY8hmAkH0Et0njjknWyidXRb235HYMMDdUaIaFuDKiCkZUOljEwjQe
By9SEyNJ6AHwg8P2Jv9VT7ve0U5vpmFP6ZIcaBNZ6OcxfsTqzdaMabY5uOE/A/a1
X+2ab3619J0fSYkeCnPOB+9WGMtENWaixyO85wCcEkPES0uM2b++oEwIr0aKi+uC
fa7uLCgd67b7NOAQk6TqSXWjpzv3debwrygxw9j245m1znapiPHbUjKEGVj9w5VK
miHW7crbh8lyGpUG+eHlzvvwpXjnUOl86uTP9+GaIzx7tYNbyWMxKWdBTMCwk6k3
G2XVei6X9ah5xAT6cayErxRghgkcWXP13Fx6MxOAfIFoLEYg+Q1RcZt43VlbA2z2
qUegKddIyD+bTXq2cMpSKB5V11rj0+sezDPly5rWzVVLFlvjGsrfCNNl2hJ7I4P0
tyb0zHSQiKSTR+Nv/omFB1wFVhNy1mUdwUaUUaovO8AtMU37f8yhKRScywquVjk8
dOhtcikJtBbCDI8O9FZIWzZJQtDn82TvUP1dxqAHxSRPKSZanJOoh0ynoIDqAjEE
+ZSpzsjBdQYCXap2N9QOE4qlJuppuN832MbiFFhUM9qciecqfNJhrEcXiw0FfToq
3cGo5TBUH//pbUnKWg+hRWHCoR4HAlWbpU7IJnM2KOpDe2OhU/Uz8BR6P4jacnHN
WqYo/Wpc4irp9kSkBxuXmcrjyxT5oBzaub164JWkTrRIQh/Oabv5ArxkE86J/im8
SAE3ZrKfPT6qpaf6VfbwupOVaRD7F/uo23P3LjXduT/W7XnOrNbBweX0/+SOxIv7
KojrQv41riXDmgIUuM4Erv3aPHUH9wXvVmhG+L1EH0DQfo3AhBDpenQy/JKEFfZI
PTBFB4F1kILIGNjs6eKoCWXT1eXu7iFxaBTfzZKi3pv/XcVEMDx3E+hvJGHs3BvX
/VkFZtzqiigyIMD8ZLjpn0xlvO8fPc3nCcKKN4ciDijZTou6iaL2xXGozmjRLwgw
Ep8iC6wSu5p0i0EBUw+GJucqJqQLu1mDZ0MVt32gAqQdcYbRBIWCi14oSB0HpyeZ
ce85hbKhcSBispe5JaH+yy4aLhavS7qiXo+fZP3RvHpONAUVJuizqewUivhgz9Mk
5YOoG3+1Mo/16qDJHuMcMJ2zzy348yvUIqf047xikjBD5GVHsxtMh/asxRUgeyj2
jfHOVMS9dQxXtMq16J8GdQ+i60UYgJW7v51fL59haWZ/5QLk0QHS6ucCc512Rxlp
1cTg2pay9gkepa1lSS08hA9/AYCXmH5vFcBGcW2/SO4MT/uQOGQcnWnT6ZbM+9se
E9tgIWyV3CtoP04fyqJ1j7RC0nPq1L9q3ZylWyHAPtv1SeOkXJWOsQFPmd4wwp8u
CZ3hPv+N4hyieIgVXhT2LSr807+oI5lpkpbScIudAqn87BoibZXmR85DFatHoHzm
f3InYMpTf5cEUVhyhXhjdWYYczTL2X2gZ+mLDjU4bDfcofXOPEJMOmtqcmqWjFJp
WN525mxGqtsL7N5oKQJf4fNhIGgNQHhEZ0By6w3IuiDuFa6JuxiIq3Xt/zp9fYGs
d8bqp9iiF+m03Lzuzg8Mq9XZxeszuOTZkImV72xzfVKDcbdwdQPqnGr/0Q+Vy+OV
TeiMcgU5qmZISAFKoKzgn1XX3K4xIBrVPfd35Np2T4G+IfEHRgvQsZClh5leEfYq
TwHl06UPW7tzxbCiM21Z9ziX5fTAkYjcBliKo2XGG3UfYmBIvlGMJuKe3+Dio3H0
h+8mB9H8CAD113eeFZ2FH1EOulvMsC8gMqF2PN2APhOvYs6uvh4EWb6oOprwUn/t
jJ6Xqa5bzm7SXqxdqf1qXAWr0Ifbq+sAFdFjAyX8ormJ3BeXITzQayjwKy4lrG4l
Trh0HRB9K5N27KRKJ9TimQfBFRN+NZxT6VSd9ihBmAuxlkeXavzRE3fbHwafMoYZ
VxM0wrYdLEYKo+WzDs9Rriaw8Op3hQ5iTadurb/beOtmamjPuQO1e0T/3CoSY3ND
gmVaMCSdHRbrzeqg8CZ0RZXylXz/WQHq5rUL/QclYLKWywNtLNSHqgTbnO8TWo5L
SdACph871qq4dwRjPACMKda6P2sPt0i8z86DGICzUuX3OMAS4aLi7CJG17YVEnr6
NS71Ln6Zca/yiseE3z5dRI2BUWBWHuvaI8KRlbLrtD+2d74+8qGdQdtF7fwJyqEE
j69rEMcCokSKDyykSSCWzmw0qUL1MlSzrS4PzDYziaQ0OildJHQHcdTDHQmOqBhL
lCvF9LeEk8ho7DDH4GvIlvVk+SWI0DkjfJgPjy0feBYsR711Gm24AxKi486DDII5
s8DT68l4LXOuOTZoX9R/xFUAV/RRzGL1J1+1Oyx4y3ctnRNdaAcH3IIAeyoUOyjD
8SBU+wLfbSkfJPkMPGQRWYOOxeRdooee6gfjIuTPlvxDFob1Rn8kbbT/zpihsonB
pdcxCq995/Uj/8q/e701kUszs4DFgrjdBnINcSjIZZT1sv0oRycBQ7FcSyYuUao7
uyo63s/AZ3LKBg25JLm0LCNqyP0bSlqH/T75LdjCO7gZOqaPvmQ5FBvOPEgJyned
AfbAND+mU3OnqmDr/BZlJrYA31h/nEoTeATOhZ8UY2M2zMD3ENEBdc94X2FnhlTN
Kg0PjSoRsrlGSRNinbWq8D+q0JbhH0dfAaRfQtgKNkg0e2Z5DN8x8Ldd4wRp7aaw
eWxIKMyCayKvo0vHSgfty7YtyvWGo4HFstFkhlfAZ4Skt6siIImPZLytah+e8WSY
jHA9tTuyVzs2zyqfTJU3qYge+Nj03JpxfUV8ymoG/DfT88kTgmiUCK4V0qjqgQMy
KmHD7lX+h36kUceeicZIHujCyFWeqCavSAUxz78xZoHYKN/tL1rIC/ESrBr5q0PC
DXo78GzGIdG/GEXrGxHA802eevhQON6Rt/eyUGrGeNXeBUwd+rUX8aqa1wk5xAEJ
thyC14Uy5Dk7eeNf2DEKL1r9UTx2mwz3Om1VQc1DvrsZIbtb3cSle4ELZsqOr+Fj
vYQHJaJ6ZMtXdMmQVxxP2DBi3g2iTBtGI/4nV9YLVerhZhZKVo0RRyZsr2z9dytP
WO17/0qWfIXs2ltkw+qVxj5ZrsVmJ33BYJ+AIOUGCobYVn5dpk1ga9AYVgsS4y7x
+25UYp1eSPyr1reEcRCy9zn/H/ViEP9Di7qKeX4TeqqiN0jTU9mzcuix55ETPfXH
RfRM7dudZAzB0Xjkwjlw/F5/TrSVu3mJNjKAA17FPxoAPpA044qWJRsIP5gAqDmw
Ypm+SOTT6SvwKXC9Gh7qMPpQKuoOLnWf3JczqJRslDav2kMsXZVyXQoxQ6oID+fO
umsuzzH0MhOnYdRx+Eh8M7ZsXKDE01SpE5UeYYJgBnzWMO2SjzKiJqrG4yl16m+a
AYqwIgycnr2+k8OwLi6XEk9/tdHTxmA7Ef0VmB9YXsnrPbyLgR0AkvrgGAac/jZh
ivllu2ieIOWX+KBKnZNvca6fumsE1evlBOZBby6HiRoy4UxuRKvmksF0wSut2h9D
KOfRsIKVBKzMtgWDvHt47qGohWDcvFAK4UDgmgSycKO0xRRrIMZpwmZj6HQucUo+
ymwDNAoRqce4494Nj8Q8TV5GJH5Bv2810/ZHX0SXrQZI+TrXYauW98TT3nEp9ikj
amE+c1hm+7IAtdvqb3HXeuIjFQ5cBrH0IxhcDJqa1zOFkAIQ3S7B8irg/gzfOAyy
QTWoMNwW+LgoK1zvOjiiZ0H5sw1wSdrvVml5upMAR8K+LPSOTNum4JA7v1kZrAkp
YKgo26lkIYw/kf3GLZ2qOWJ2TJuTg/P0LzZKNP3JNSNli7P9t63Ct2NZrSzlYJZ8
GNt6+ryhScqU7od8tdGLtm12OiZPfH84d7vQfW3rE/llCHJG33DpsMX+jHNofcLT
CKvpZoY8EDmzRo8mN+n8BcU0OiMzhTV2x05CQ6ImGVSLX1VRgrYpMrb8Klu2mB+O
B4vzQDAKnERNvm5yN6OIwQB8sEuDDJb7PlBmUaF8QZW0BcBLRPf6royv0l+uUtGN
ckveHIzZPA5LGOxqMEgPn892dngSHFdXUs4HLfTEOdZ6AAtz1I0jDcz1Kk9mPpfO
Em5TDsPI193LSsF98xUw9dARXJXoNxsbm/zlH1CfrqZk9EQXc3fgEQzIbFzRtOop
RViw19RWguWZhDogvDzsrmzyuACvk3iZYZDSsYpM0fwApHZKHRlbowk5Kzp8RO2b
IgGkYXEmhK+j41aWE9ygLA+LEF5Lop+zt81+7CSgkmUIyKD3Gb919oO3QjewlUr6
Vsl6/9OHnT06/HPWIDwE8Y5bfNiyojU1Ces4Q+bcDGGtC/DQTC7PEwItuXXaNqd/
NHvpaDH1htq3grcI0SNkgnMGNF5SLkrj+JhwJKZOIaVkotQYomrjzBtszV1kUDwc
U8rTySPFwsqZUVkBPlGfCE2VKtPVsePyfvGNZvsDoXA1JkijWCGv8g9SxQgXD/hq
XbuleZJk8ImvgxaC8iSAyczz8V+Y6yaq+hb2jlWrXuveS8Hp7Ef/o2a9EXMOK6kw
cDW/q98ymx5CZTXpl3KBbnGeqUfQoNWy4H7Of/058eIP5a8qf2SpKFlop7Sgv96y
LEPmCTzg2zvrmFz8wBky1yOQjAxHJ8mxdLqRXDX7wQO610dMQLIGIJMa/5FP8z8O
Cn6zqt5Bj3tbhT5oSXEOWkHJH16bs15wJJjLP/1jijx3KE1PEbdqS0adQ1tcbu+M
xFZoFfi1cfyAl6fH5kBlWLK1E8+/hcnlOLCKrn56rAqWzCLMBLXOwiTG5V6V2GrN
lO2dWNDNHE9YkmAAIyn8PUEdy1laOLimLEgm13KnbBU7nhIRIHDcIsMWRBnuW/Oo
CCSV3di2wkAotc4jdGvFlDxgnYl6WnZBIDw8inHefvqiurGW60OtWnIkkq8W5omo
QEdEyBpIAkQ4aw5X36De+dLWA5fimGruIBJcbE4bKrScvRoQBfQq9RCFCHvn7yUT
SPmyBKKyLNExhHJHvhWqU9MtexrUKOVZAmPIKuN+uo51UFMDNEyCNmxfPJA6QaOx
tsuhRwvM4JOP6Jw1ERSCx9JlUNb6YfVzW3qNf5zUTSJ1M902tUQnuY5FKY8YLD5/
tyj8CvPAU5ZbXiGpjImvNk7iKEqF9FMpfQQmeBSBaA/SliwT4N93FVFVOxR5N6an
TuPUSnfIK5Zz/leAaFWiPyR4K0F9CtYpAhUAkIA3OFZk/D7tVx53ZZy6SK/0F4C9
2RQr37D65cL9HCHX9BkYIc9t4kLUOVGO43wUi+H//Tlubjmbxuazorrtjd9BHRoW
8BiQlFIAUf9r1G9qFNUJi7uwEChcX2Q3oxHkYaevNTyuOscd48E/T9uTVmXRAlA2
GhC/721iofmPS2lThMxcyTIv5C/IfGdkvPSuAo093aoB+wIBcODGAoVN9vnvgL5Y
3Sfo9Ouggdob4ZBDcc4CPnMYKwV/IfZpe/sleHliBLorz4zjgLNG8gYx0Wb01fze
3uwEwxSaw+FSPiGQSL5men8EOgTlDi0IP21Q6NsjlV2kVnyy9HKKjmZ0XoSnyih0
MIS47x9P8NKHnG6y2uECZ+EIcOUx2VBg/4MFFIu6VErHC3n2R8HHOlD238Xn1U6w
B7Ny4KGMSRnGsYQUhfb+V/7OloGGftaUzXgf5cEylpvH7aPjRgSxTddV8iZ4aKJP
E1jTLgWh1DqQl/x6MnEkh12dI+vbTL3GqGKYk9AIUdBxh1ziZu9aPUZvRnzkpEmv
zjsB5dxeiy9KB3/Qm3/W0CO0O5pYAZGZrurYAwCMmpxgzeKgaSUhVuzTUmWwp8tj
P3knYcbvPl/M0gcls+n6BOTHH2aKN7tHjGGaaqj4C0ns9C9rN7leUn9KOvLME5PO
l3ePfKYRZpopjbic8AJxixjSvQVObpzALPjG0fFlkiRpH9+GY3hgv8CXYD+82Uo+
bItEwfMIBq5krzfAoelnE2GnSTVZtc34mnaecpISASpMaxB4NzXxWAqpnUYhBT8U
+pLMg9wO51MMduupp3uigj7B4xUlA9g4HchC5WxZ2E3iRlgXdZAHxMUrW9ppmq6P
c2wb8wgM1NtNdTwZG66tLZck66rlwDg0FBklYGzWdCuKXbbflY+EZCGBSyqIlQ+5
6ht7p1wJbhazATXunagqDgTbaWGOMT4f/57TU/wX2kCtBpmaHSnaJUb/m15pZrd7
gKpt92GQOE51LxEkx3eQhQExY4YeR48ghfCmpN0YxVqkSXHggtCI02HepCTK5e/6
VQlTXHel/NRyehiKCiJ0MtPtTQ6sLL+M6nMWd2WN5XDlXkkkLtDri2Kde6KEDW9W
VDcwnoMKL7BK+W7iCMZxRcFjYcQm4FKdw+a2CfcZxFaipo8KoHtos42c28XYkPPS
uUGzex5Rg3QEFaDBanNZxAg+AyCx9ulzs30k6pNoDE8h2pkmPOPGKhRRLIC4PlSC
sQ03L4Rk1JTDAcnFTvBP2jrfoqcSr0k4OW94yuUuTjoIMY+MSn70iro1nE0Slatx
/4e7caDVXyofU9Jxjsb7o7dpf4drLsLUBihgfXBCBCf9GF6hLW4XQb5nGc1DcoUh
jjP7ARdqtWQiR7ljiVeKv+6To5o4/YrnluVZmf9iI+sZo2YETIwaWoWtGuXQY2fa
W+eVGvdmizgBrCZgAKsvoHP4fSnMnlEnLnx2UOTCXQVoQ1lJx3+i4SghOO4uWUIg
v0B/4eW/0E6+UmAUFH7eKjtPxxCv/u/uq17gNV7T1e3rauabe+UnBVO/laJz0uBt
gFlAW0y76Qk0pF5//rOCka3XRzS40EMg21qxOzNYheJk35HZ+BNEDIAwN51YM+W4
FAK6Kmsbl8fj3iajpJuFkjc56/3SPFFAps6MAYJzhtu8/z39MLYI5d8Mc5qr5pWT
GHvRfQBGFp8YoYSCGz5aAtKYaURdAV3Z0uqGLGJeStNeqr9UY91dMrYfixBXRjGW
WKNPxkNDMnV5U+CGhfkiHAvfx5aJXC1QV79cv2UkdFVqj6m6SWl6eDIGI6kWov4D
iE0cnEt4UQI0h94TzcLBVVqIGS/HxNl68PDvMwBPRqqkHKhDZojtuFetBvZhMPeV
5E/r4WqapXsqK8AaSDwCdfKk+uZEz1l0o1dP97WgtxGIits08GVfKNrz2Qol8X1y
+q6fRZOyZqhUCoDkmUuljocdZGslQ5LqzZEAEhL4K7UCo6kVV/RuCYKYSgrG8BTD
vZmyFTmO3UOM0hkmOnYOjHjGu5G/ffpWIgw3mqD6CQ5GhlFZ9idQed7otF0rZVvW
HD6OfC56x1ac2z2C9+EwnUYcpIk08wWsaAE9f+VpMFPXwmJH84Bx3mE9KUBso7kh
M0bLuHtIwH8G2ABwDyvgYg1RTfA9qfaeSRh6PEEjF9kLSllCNSkfrW5rQN/Xupty
+7A1S9U7bQFPlR9QgG0obhobTD0WLo/h6LZDef6b5jsMSkr/iWaBB6MhKC4S/CuL
GInqt7A+lmgSUmrGUSyqN/XCIXUR8VqciGjsAcH7NkJwM8SC84fcal1vTL5+SY0X
ASFEZjEcODrdmH+xG1WNadJySIt+YT7zgWDECU/kNdOBJtamAKegvKks2AZQlv+B
WWjyK5IkJN13uqSkkXrzpqQfv6QB08gkACAlP7hxYebdaKAnf7EfSL5c2kwVAJl/
72397ApVKlxxYWl1mHQ6vqznW3VwYhLGFEDpEILMqC2SdMbyXvF05TbDy5ynMvYw
fwMRR26sb9j4Vo3/3SwyZzTfl7I7WRHPI5UlYvOgsDepBCOuFc/mW3w+j4+IUEEf
ZJUxI3RrAYV51cazxyTbgVXp3kA8R/Nl57hIIpmivrbOmS7+ZhggtXuS87mw/UC2
GTlaWZdFDaOeY6DgDEocG3PF1FXG7qH0HYx0MD+eS2jZ0JDZSzKCHHPti3JGgsP6
FsojlB0NqpEJo259bvhLMUck/UWziFsEQhM+qu39/NZNzVKGdyfD5TQ+fQmsDZyg
9Q3shyVCM46n7khFBaCXMo3J+/Ni2SwdJQcu7NzrSvZTCiZC3O1YHVcjs7riOmGv
M4nQUzD55mnUNSqQYh8K170DYkD/H7qGD8Jp+WQG/2x0IwAawgjjfZI9kGStz6Ye
nwwJCmcNMWpHBif0LQOcb410ts1usFktgv1CGyXVlSeRUv1YFZdks3VQnh1N3Ofo
8DoUMX4E11/gfVzi/o17K3U/H+k1bg3E05SlZkTSScRlVbdqG4NALTfEPq1o3q1q
owvtgR++NoKave4X/S/8QAoAP8QX7oP87p/elpS0DqsCqWVjbHEXdRbcj/oVSqrB
3OHsdYoHcixvANEsnHy/iA7fTG804ncmTjefymhLepO5xS4PFlDZBDlY7TdcZG+d
98TVexI7fQ5+h0gQHDKfXKeTA05avJsgu2hm/PbruBh3NmPmUBs/+L73V21sUbY2
Ke9u/Vslrz6ZvrAAYfCC9p/VZsmRKNeg+elrpBJyGeZd632K3SqLzUC9A3pTbj3c
7h7YxYeUXGY4ZKnBnlFuMCK4thveQ+GxcHuER/tnvZBwCVaCA1pkyBqk8aIx0jfC
x0Bw8K4DcGIib3MkRNUQ2UXvLk6Q9yZv9lB5vjj3ztwgZfnNeRPDOQuqeLekgevZ
NzBHf/gl5jlhH9Wey3H1u9okQT+a9lFU77RQNdUMPMiJnBC9+7c8t5L3azNiSbHu
OclHr7NbPtDFhRm9ilW/F3Lc7htVgT3opJjavR56Oz3wF87Fd2wx6TC4MprcKPgC
GzXd9/ZjpQg4V4VuU4HLTi85k6UbWB1i/uxBzNVizjy9Dp+/tapW9W39IQq+lr0X
bQMVfWXC/99glf1y0VS/H/1GGoi35HomQOoQlCj3hODJutRsDvZUp7sUt5YsAF0H
d10DzwObge7VKwV0bC7nBl0a87bSRxYSJd4cT95bR0hsVaCTxen5P2W2ukBdOpdR
GQLBtL+ijksWyr9Qyxn6bEiTE7IO480odlVvEvrisNmcSIPoUCUx56Ywl3x/nn9r
3r58moOkgs3T5TAMhwZW98s3QCyeKgZvYJwmws0riQagGmhsX1w/M+PlxmXI7cYl
e0FiRXTUDiLE7WHkv4XVkx86JDEcieH7miwR2n5OqnwdfLOjKAUOgf88oR21H00D
r6fx7RlqlqtPUW9fNSCtUE/ctB0P/pJkkMvawU4PU24ELdV9kPcMDsH/bgZeeHhq
P0tE4KSmjxGxIyUmRG0yM6eGaRlQ6PSmZWpxC8/2ee2u4WkUvcwq8g1YKo9Qsgs+
PNbgxFrHEVlZCPTaNcP4w5ntYtjN1pAGw+vRkOEWKMHjvSxi6p+9Wen5EzKZzzvR
eOofGP7Aym9sAdyUh7S8ZQaGLhU15wC7zLzoVoKK88ZPi0UXJwBekTV099U8VYSq
5c8mrpzea9K2GcdIwpTo44rB4QxWz5UPd7weyaaMKWildcruVmF/KoHfp3GNDZ55
xSZcEmCKtBqMwxiXUwqEtYQKF33OD6ZKbNj2b1J1nsu5WP3vwA+IUlqvwKUsfN/C
3x+RaT4shrKtIQKfY/QBKUiVp/gtarGx+u7DCL/mEqVwZkBJmQTwoGXuFi6Obmxi
zmSVz76xeeLv/9C/KouanpxeZGnoAxfYWU65H7bSYEdgBMxT8dZZJRCXwy8xqjYV
OuTpZLgs3u//wE6Li8g8eRWNFEvY2S4bKAkwIlwNZ4F1bw0q8eA5vs1QgQAqan/9
7+fVSioQUo+eZtoK6b3+Jr+EEjgno1yDZWr7Kph94pB7g3WPwlfDNLI9p4hdvWaq
BD0mS3PmkKFi4G88eRHAAD6D1bzSdJIVecNS5gLYnXfAUrxXIccq8+T8oU2ZjpCh
f4sK5Oc0YOHgjrh+blpvYMwITPMFVRviJtYtFo3NvbXgMdlRDkfxCS6941/fwWs1
MIguCg+dYIjkkDbT6bFFOsf4VYAk0oRpMK/d+t1k0Wk8PseAemD4OByBfZVJT2GP
iRjU1JRDsqAONhW7v+oqcZIzjhwu4IqW6JQbM53p/JAPcIIkONnGHHfD38IZTHRa
D7agLbT3HgqMEre/5Kf6wNTtxTORKc2OfKFTokPXmZtdKNn9cxV8cqXb+oM7CHQs
0xXaQi8zxDG2eUoqVoeskrSNJBxB9dQFZfwUDi9tJk3Z9qNR6wZkEwk/SthhbZes
mLEyS8Hd1a9gCxSNkJWV2D6m3TnpoIERNf81VMDhI+VGCJ3tmA2yOSLrKU1yOZYp
IGuzthOjYo7Kk5eLD4IVlkp/PJuQEXEwZP/2tud3v+JIxBeIHSafiE4v43aBGM5p
FkO+YEMdti6a0ZCpnPhbkSV0ghTroqCNMyhH5vXDq24FB0DC/1qPMXanXE5yvG7B
qIcUq/SanE/t3yjS6o72fJ6JnS6q8n8apXiyVPHR+84OdAVDswmeZSIT12YOiDld
lmp905nWx3SwXOpJwK7S/5LaP67lxEC0zImASamDNWADozicnqSkVSbC3AFg8yOk
fql17qaTbqfLs3uTDbrK897IQyJ+cCa9qoOKOamVYvFRdSBTvjFiSdV7O918WOwI
mb7wc1LdFleWXYoZW0vW4b02q/gUlTQLtCgo/+P8A3UxxtEPNhGocI7qvPcBlKp4
Ifg4BcdK4j+Ddv3bPtk54B9dWBosKBRzV4w2Lvg34Gnm4nnh32u807omvxLb4IoJ
+iJWrBkewCIronNoBVs7F3Q9I3Ba6LJO7whoxkPT+x3+uJJtVn4KmERx8z+0kpu4
Tfp7yqYkufwGz6/Tp5G3JkDbUAEApH/0XRH4+facE2itr9QCRlQtn9tcwbcmZiZ0
dOiUHGOi1pm8Y07uI9gMxKQ/jqmsPjwjbnyuvgl/rTuHJ8uuOzwo7Lu6ZqlHLQIt
R7FXs7gMgGkuOFFL/yMTdvSZpTcJU8Inm5oVb8J6PxTnOX8tDo6cobA5AilFGG3V
KMdNc6JsjVENZ++4G2XPbO8uCDnkSZqHzJkM5wZ+WBFMNAZ94FkmNxQVvdwbYdvG
4VhCoQXa71yTmoMJq1qXZU/sBdYjjMfUi2Fai76LVy/UYbIHlk7KMmq0vJdVOvJo
27mQ3oKXwbgqDR0Q3EAzctozf0FWd3CPDZwqTislXXma1N5Kj7KWw5B2shzWeLm5
XNQAaoEiNC3XA/1BHrBIfGhr+peLddtkuFx40GHlLWAyXBWdpO+ipn4YeJu1TRYs
CuGJFJqL+QHEYjfOhdpLP2WsLGvfGYQOtSMbDtRsx1On/hF0YsMgKLCaLWyaEWV7
6MQ8y9XFWejtkBHQX1KT0I75DHNInB2qQOkqRTYHZDOCFOxIxCf+ZhqddaA2seTh
xAKF62Xs6TqziVWJoYl2W3W8/in9nYDiUGoxZbRqEXxO94KnEbmRnIHnuNQiI2X1
IOgx1YL4NApMFoaZzJAmhkzioGSFxBhVJWcVj/sD+VDNP+Ov706DfL8xuAiBJQNo
336XC9Hr39HQ7acfC3WWUQ7iKT31QK92N7fV4WaP+iKjk0/W1XvWcsMP6whAFoDq
UffXdrizJTGvQB7vFM6Q7k+pWkcToM01i++eTyIT1QY7Shyc0jGLFrLS773wF57d
/+Z9jO1A+o/q7QyOdBtIHVt8HSIGJ9sRHoReqt32E78M8Q62cdTNvfEDf5OIPt1h
Cc8sOynMkeVHqBZZ18gtMlqUPkDVvo8FD1MBJ3q5lDrUPwWfJau2E1F2VtNU//Dl
fmENTcoqzuHcPgQOVRVkaUBLE/E04GwZUSGHbwCG5gZSfQAACtZaLMr9hY2Z57Za
dIP05ivS4Vmrz2muLKW4zO5jFqhccKKSNRQ0Y8uFDTFutWtHwby4sZ84gP+LsmT/
CFv29mj7zfUgw7o9er6CyEEOajRXiWVXeTH0/Xh2lwIRITR+RgeF8EPGTn0lETiY
b+J8iofGm4bLPHQxDuJ9vqBATzXS0+RRoxyBPTPdF68mJNBwnCYLD86AmRQr9NDU
s7JewWv3q8Oze7VWw34E+VwHlQCLGOC524dQ7U+bU7q/2w6aHhN4+L+Dps5TOAA0
IZxWclFWz0YD82WjPnuQjWucNUEsaIRdV+w7VIDeOoYd+xPaUHOsX6aUAKdIwDJ8
ct/dpoAU4/V2v6iMGvtsVXay58s36NJZEdh9VGujPUfDhRSvkepFjPafn1DlgCXm
DdSuEXezmnZ+tYU8ACLoJaQ4OkkBvVGP9qoZ4SbCZpuuwn8+yXLBErOKquvu05Z7
9+FdyJZFv4yVehCRV7v+eZpxa2Aly+ma/4K499OBc99n2ViQfeCv0213pdpHbozx
WFewxgqngEVYRmEWfZ/gJkVbinHUmcSfiJRXjIvCelJ8O9zBbhfptUv6BhpuT8oJ
5Ri/71acz1N5+VscNyXflwyW+Uxk+e+EpEXoncHZwvIie7RcLT1brXf8ijnrL5qK
XwY62Pc6W4Sa8jwbufY9xCmm0M1W18YQzQ370puv4H2CkhCwy8bPKthfSfrgp+Tw
w9yOt8dXmcYmHPSjZmWtzUWSrAj+tEcUeHOMrqZpXPTe8eDSKf2NsvwUGIOKgr3h
cLG7ScK6HsrfNniuJwuek/+bgOxX8VoOQmjNpePkj9jdgWk+SC9Y0o4MbVrz8Lvw
dGLlU3fBK8M84lRw6jkANIzLLajA3bDgrl+lV4SOJ3F9F/ANRjQMBy1qiNrH9tfe
dhVu4NRC9CKGZldDxlWqTD/7XvNgFVAdJL98AzkfzqxhOVav1GMEIBe3MSBJ6dAK
pD1i7CVkDh9v0hZJ5dPq1gHCcJ2ZFtV6SnHp5b18TZ+VcpQne3f9lbMULub39QL/
6kt6+H5LbRs7PMfQfYk8TywqigiT8dYpiH5GIhmyHzdLi/M3WKoIEpwQm4+4X7Zl
fvkCITGMaDvic+duKiedq8lxx0kcDNb82TQq7Aw7gsx6y32pT/VkdVNEwqaxYwOc
M3MJCf/sZtR8wcWW1h/NXykaxeiDzyEy/K3X3fMKgUVSlZ6VALTdb6Dlxco1fvMp
inbZk9rRDsZArArRMd4a+o6XQoVMgggqzCMNGJwMlA7wCSp3CXdhCvnS+3tQzQQz
DPD4K8twKNg4RxwcdEX5tooOfnMyRFlXgulK8DEmeoq9X+W1WqlWOluEtGH9qyqg
U6U6i6WcLOncVqr2dRiVIzzdob3MxmVuWy/7tYxsAHOmYBKjXVvPFgL57uV/bEfO
aX5hTIj47iNhTmmDwhyg8qh4A+j4UBDEygZ56wbj7CDSxbQ04zQxHRmPk4dep371
+5PMC0GP34grk7210pUyvnF3qTmNyvmYX5EJZIk8+mJOf4YZ8GknRrVfUL2+eMpQ
J3cLiSGRFxWmwAZC1ZGji5YJp0dP779KY8xG+Z/9+cgBCKNA+NkGW9LnIb9EfsVO
lBA9QedfeqdcfL2p9QXlvjt65dvGfwS2VrN78xRYHjpKC7lbZ7AWBwtMmf/r9kzh
vOAE0Wy9IHBJ+jUmZ5LQF8NdM5GzoV732Nq8hOuBeRG/EoHngasc9ktgbmIjLRGA
iAmztw3pJK7GsDW5YPUNgzpT14hlBm2CRC5iAcfor+tjK+mROQGHIs9mL3d/HREw
EaCeX7ondwLSRLuaFzX5GHpQ/Zr7lcV5EiIbf9L+Biz5KCyKDvTpvo3lk0+znVpR
n5x/BVtUivIiKYU3xrpZRt+GXsqCsmyLkE+FCm2W9eiLGlsRwp7S5QQVptEoWTZ6
J/j7DXpJnvrOK7MrU6Vx2YJQm6RNWPLi1QI20FddYXmdaQgJtbeZRnXn1pPRJCdm
DjfeXUGIZLxXwcJLSMsFpk7V6asBol/ksbjFqDRuLpbQxr+VZ6cMmg+3XJKpOGc/
nl9f6nmbotCpFfnuEmE+/UgNyI75lA1olYONchMl7/FINAXVhTT2UU8dIDQNZC0Y
CKT+9et3WnqoRShiHwrnmPMy0RKV+O44pHu8StDdE/1H+ps4KwHXMMm0i38z/29O
6JXG9MerDYP1UCErtHhI0S4hxkgsFTOC395pOor069VaJMqGIO9xRObXWbg0l/fm
RxuhaXDZI0czhyX/3qE3xQTD+pVvIPaI/f/vITcldsCjmC0PVl+DtL1cEQkdAIRz
TBVJeKvGBRZaShLc7p2GYmSPDaPqiDEtkzHkXPnbrPyLQMI1/PNthz9DxghIydKb
baNg2mBCW6/tzVrbE7RFWHb0ExrcxJaQ9xEAPVq239sFFjhjSEpmvGHjEXEMD9rj
VlAvRMb8oaP1/2kxDY3qH9f9cZtJPwQGR7shsgIaWkVtuubmIGd94L8anJkxxjRJ
PUM6C7SnPuNRpqThe1m1yzlNB1QKfImKrVbWDtBn3n6ZSdmjjI/skHegcmvblhzy
w31eQrNIiOL9xYTqy+wvM+Yfv23zd3+Yh7xzwxLhXI5GW68WUoDbr5Gu0zFKkHgo
5LuaRGI1iBXUJ1WBNqteg3Q5ETZ5/6EArjH2Psl3Zh7OlZmTWBzuJ31+SgInC+8N
x6GgBGwHoneCU+KQfJk7U72SdRv7wfTz4FH6Wvoofr/hUHs8PQkMuGgDH6bp+Bao
Q8eSm5wZMkLAr34s9P8R7721NbkkwILFOl9lg/NVnJ78l3BYNpC/f/lA+o9bek4W
mMxfy4QbzVCI6IgU5ne/hd5bQ32lqXiuJz6dRZDrGCIj4gkuWs0Qf6YDrsZgxWjY
LI8fo/MkrE2rOO4VChObp6nYfF5dgQEZN77/IMjiHqK0sFy2SkCnzeIAOTTJbo64
kfix84krLOgy2yb1r65JXlSRWDxjOriVGSmR6PdLB3nYcJ0yqsG7omqmTqspgRDv
wyoj0ErSlXSeRxDSPd3xiaT0SBWqP0TPQeCFmqM6bsjM6pIFJnjKZZDIfWO8ZIqy
ozg+Fjqdm/12YHrdtlniGTkH8M8ItYNLPgMu2ft7pN9L+CYkjz4i3o40LGOemAYP
/ojuZkty7g1l4phPeo1eDbpdTsakprg8yR4I4tQ52uIRr+DxgkhXHIj+1CpjA11a
q2TRvF76lACWe371NFeQy8u85L73i4LR5WaiycnkJay9+Ckn34Nqt7Oyc+arNG4V
rJH/sTEcFtlCcDjF4FqdjXl5M4cyV5i+fxSZB4dAU1Rqv1gmsxOvOO3qOGM1x4vT
CK/Y2FIAJfWErhfEEtiUMNags2yXhjUYf09OPl+gxbX6QJy27LXKcYDV1TKKwIVc
qamk8BJfWlaae0iLNcL1wLWiWRhJy0QRRsECCkm3B4eyZ93u4os28fNHJ2QQRoie
mz4J5BTl3VFqmZTlFaH5pYotdCe9FK3Z8R6ypCOkW3kYUadljwwUFqQYjFhhbILZ
Tmw7yfFT7E779ueJ+3NERzRyUyHFwllgGhsANB1Pvz84QgT7B4EZLurbSgRDkivL
ttpQQC7kH81cuT+en2DT9wSktXW5yrlJTXXJia8dFOzu5HDTb/WaFQl75/J8X7i7
Zat92SDa9C/Y8ENk1HZIpZ6bGHae/BqEJJlPoVwllIm1xENsNv5s3aQUAI6+BMU2
KK3HVxXtveRB6nq1xXMexhuX2S3KYCZW879Cm8vvwL7yHApu7JcVj6vPRZzeTJKD
UxNzs7AqRRoYhxgl8yw9ElkfsdwDSmyuxWM53W3Dqetb25DBoV7DCSRknPiv2r1u
Qr+1U4wBSQAgv4Ulm7WGMl9WN7ta4rVHZyPAPjQoHCAMgv9A49F+z1oqNkbjWYSx
deBO5EYs7tvaCJJz0G2IY4dlBi6kGhMUhMLRCLEpLlno/xGDLe7GLKYQjQru9E17
qOpYiF6dt/0o1mh1b1urZdWp1XhLDk+85LCAJrFy9bp2OIlEVfsH/to1oEw9w/do
0xh0rmXSp3oN8aFV5Sab2Dx/8V46wIiOB4pv/LxUW1+RLLiLyTU64LnWIQImzbXK
T59NH6LwrDjoTvTSmT5vZ4sxVnDAsdNJ6AVFIdqwVRmAAeuhChOk2A7pVg6jRCnz
/xHg0hLNhgmp0P1Vssb4HeVwNxtt4j+ek6Tlby8H0dud80GAhVatQcyvD+ZTiFM3
UDVySd6DjPLjzI039Uw4m34sfe2wP8N3CTp8rZJ7/XiNSryI2DXMzsZlTtVT0GWW
qSeY+dsnj/a99YiCfUa45A7SFlhu3unoH1Il840k0RuckclL6HG3H1hLlp10Nek3
nDdecaoBu8gHaeNbMZvww7YHRu5DPtGFdbRNeyQs4LR7N8xO/du5M9UEKOz/bFC2
UIN1XFd+Fn0wsjtHFkyUMdTHLQIqPppQn5i1JmxIOIoEEQHMuy8pMTv2o8/ymr7i
0NKaIx532JzxoEvhqZ8aHUEJpKpf1b+pfqKhB4i5/g+OOMMLKOuk2QkE2YJhxLW5
MyYgjwSlFpjOQjZoSk5sqOX5UV8DnwRKehOUUurwLwQrh/WktdC2CzQWI+eqKJ/n
NbjU8+vdpgQtMLQITdoYBpX7vHLLtU/sZkzdq+7iK+pMaLigFhxXbsCKZTqecvdg
b2yD6DOjKq//jtal/ce2v5OhPash3k2p5FEVxeDxbsvLoOwo3XWjEdjqg/xwtePX
zZ9E0Gz8ExD1177jxj3N4aD/8iZB00gflaQQab0XnYfO35hXErHpliQfwDKuWE4z
d4OWGgY/8Bs6IQiBk0MT0RT98KSS+MydURwuV40XZlKZii/QIIrXJZr7A4BpuKmK
c3uOd4HiOUYcSQCvkEjJ2fdq82NFbpdBn01eABdqMjXBa91n9acvuB9pr2EzxIJN
puvUL+a8xgxikWa2GVAe2r11F/6lewdUeWP9ZagQ8PNHOd7s7soecVpW6GYbPEZP
ZCwN9ZzZfIkF+f/E9BVDl8kyiFGeVbNWM0i+eX2U7oq5zOnp/qDNMILidq6Fjjq4
HKpVGF4fWpYnvEVgBFMMjtkZ4HqejvwtU/AX43NT7Ra57EV1FE9JF4rI+rztCB+V
GfL3fmUW3v1oA/b/kBF8untV6G3N6P1YX0qjd0bgD+t06hyK8mDdltKCGLb+RboR
+uFUk6tuSTiEDWrnC0e3rMq7vjxVBXPPRhIZVhQMYw9+fUKfxLorHtbEih5cqeNd
Ra5bRlZi2A57/sKrfugn7eeYpb+FdBNJQ+B1kJtCXMLjF2Qd8zWnL/qdnyHoCdC2
MRCp8V/eh8tfBCxErslFPUoplH7rOn8uomKrhMLxfcePvSHAtzrv2edJ8qbWIO7J
nHPA46vJpHmAU93v7W/G67b4JeS5I9ykxaaXYn0kyni+iqVtYDEQ2FUraLDozFQR
nlnjiTSo8li+LuJLxWKH0rs23JJ1pgh4x0tTCOCan0ci1pdgcdUyzI7XcDyWq/Pu
4YzLjwcT8cKaeNE2leP72fOo6sPz4aSXo6gdhcuo54aWrWMkou8PoxiaiREtmXxt
d0deYoSBmv0f5jLDhcbB7caFIJaKpNNwDf7ivQZcTXnARuzqiJ326BThZLBvOytF
hN4jbSeRNd7Im18XRpuCndGL17Y06GK66LAd32qriHpgLP9xX/oM4P3b4CLGL9Yq
rSk0HFL1hsx3DiW2LxZCOx1acmebBsSOavbSlZd3e+Ng8SzGnLGvGUogpeq69i7t
5bR6Cm6uRdZ15y0FQwQBGh9xPximWfzH0852y6bqh2tTJm8h2oTwHNltkxuHgsCV
tAR4Nui9fsZTYbhlrs/yCL/oYZg8YdzrmqR1M6AeaSMT4Y5T8ot//NYirg0R9ynj
i5CayD+zED6+avUEl50Bb81HYSqb6ZsUL1SD1YH0Bw7z2jWFIqxkSMxtbwUDvWeY
pXJWREq2XAFHmtuoasRhlCZMRcGihv6wSHJoGZ1O5rc+7+U800S3y4Fex7pHR1Jm
0XxYDLcPobIxt1acf9TiQbARDGkS8lhC1R7nO8Gl8mM0LKh2+zNyn7F/aV0aE+E+
+cOuzJ2g5oqWx4a0s3zp/27GybVPYOzz2e1iooq1PfMqE6LhFCPSE4CV86bg6BF/
h8GGGZi//wvPjIMAGWWNpTRhYNkMrCv9isXpNdHiyRZKRVPf5+RcGz9WoE0Hr5Ti
lYIgjRXquabnXMG7tdzzts5GdQY3IguJoY8vOE/+AV40rnff8qPujOrhMAiGoTlt
ukU+1imh1jtbhgMmdZoN5tEfMqGs79ERbf0fJwrhLSbpMCg1RYZPmLV4jma+mWFM
3gItUr6Fcjb9uMAqXV1p3JlPPOU/nxOOFMC58NI35CY6OzkBqKG+vMVka0zdSsLW
+oQMrpxAphZzHN1iO1oEyZ1SOgfyxa9YN1yyTAKneddxFhxc+WO/iCgpqoNz4Wcz
468l30FaV3BED0O9mp403DDj+qd86Mt1aK3tI7f3I2jSzbl85cozJltgAym9ZdtR
8LItlesLcJ4PCIOqjqs+1KrPKhGnV1h8NgDwS/xVioLt7yJsGSum0JKxoBVDPkLk
twkEJVTXvF0HOrNkCPOfqwNuJ433f+p/Kc9hzvkg4IcU+ZkgOOn7rUbiqrpaD+Uw
TXrunWnRq40mAgiLtNsEktoWwXfo5+tQccIqppdFI74R528WYp02E2tuYIBEvqKo
+CGz6CcZthqSgEu2RtNMdk6vU9lPLyD4gTsZv9xeBaOXSmZ9HGjZEzJ9D6huLsxV
77yHqQVMkxCjcfzsYYM0E6sl8d/nFCx8xyM1jmAYFJaC1Pi2QbFaaKHmloZwoJB5
bYekDOhA96Pr1vEERf5sTm/uCnFLzV+C6zUHdhJ0ItmsS3/33n8NYbVBPmjXJ1MT
Zp7ZgKGNFXEOapKmesr2IqY4mOIGYM7PzTgiCERQ2nB/NKx2isO5/xkYo40V01Lt
QZ911NUzEOLjvfTNHMHRcqD6vwkumWQ1fsaPBFOqwPh2VC0OJvEl0CNXV7u3B/67
IiIKrOy6Iy6ppHcIM7Dy120mSMANH1ziIxmiwjuhu53NKWBnh4E7r4sBssn8mc45
FUm6lF3rcDUwmqjlYDdKZ9qa4JdnF8BRAhqL/F6Za1wurdB9AlvWPhVz+zKnR3hX
0fchTEwhaZef++yNPMVr79iTVNgZ3SBUYoFCJYl4DxbpN7R54B9oghemwilkGr2/
Qjm1aJUCY/TIF0tWWTtNR3cpLjGo9kgk0bxWOgusbmqHhCg8JAdG/CmFwN0UKzUp
R8Tw1LJutjS1tRltiz6FD9HBjZ2TSZLKtNnu1TYt6JmCApF28qWN/+0rV5MieKIU
FsfFZVxU8S9Y3mF8X5wM2afm04jEFI6T2Bi9cQw2qBWWBCyyX4dGeRwWqOq8Ecxb
GZQujw7aQzH4/9AYUpjCUPSb9VMAEFfJ9msw354SLpd2k+JFAx59a1PBPMDT2+q0
fPn4wzxSRLLbXP101mooaBWbBoH14csnuwxPdq6qJdeMicGOUz2jKd7Sz0XY6dPc
WP13r4MwfZ7sIJMeqAbVz1XvAP21UglFhndUv34hDo7PPVza6iTy4tdGWUdZgEcF
Fp6b8JzO3Fz2dwdt91duVaCmWK3Dq3x0WqkQiN0E4dYsrFKcW3rAt1n0eTWf52fV
pxbeVDXeId7Wuk0DK2Ort9YIUi0aBtpboZcEVXRAN/vpu9VMvNWtN4orBRIeSGyW
oXDMPcmvUUhnFAFoNBVJ4qy7GVetuv3cue6jO5egR4e27njxhRXrpc/s10oZY/5X
JrBPmA2EV5z9ZrmBcbtFQm7y+CfzI8j9t+OLn2a6zU3/29FcRjzJEWMgE2YIb5AX
HayJ6ickIURRmh6jGaq8ytIl2PoMJClq1RWwCt2+9oX9dWk67ZN4sjJiwo+gls6J
JndkXH6KPCWgQxw2Qm/A/O3tKAGX5+O131Rp1RyzXp0ktmqBjx8n9SqCIZ10zUuG
yaYd/2TbQcaxZuDPCe6KJbSDGC9+50hZ/ETUSizBa4l9ES4gKUuBkplTonGbvdft
CqkV8Oy5BwcCq6EDwB/8XBltymK5b1C+y7mp5+Wa3xXx65zpDdYihsew34RgsLuA
ZHhOYh1bo0s47Ot6TGiOrxrQWK+xwWC5AMdmZ/c6qmJnjXLDkoD3H1XAaJWd+lQW
oUhp2x5nM8UNhFICFTVafiqvDW2evgFzBHMoGo7Wpqu7msRYnbEIUVUZdvQCAnmX
HXijv7v64tqr9QE2NG9Rg8+07M+Nfi9YLiaILpriZaEoDWtbAaD/pHVwyywrnliv
3MtZEVf6FF9sBURr18QEhzDCwAh+uWwX2pXYNU3B7gQ6hMcGK20P7LRSXRe0y1lP
gfnUZTPsQy+6EmvrD4QY5etFX5bh/tuOfqyXvfAtD8P8xgxBB6wsZvwb3yodDPJr
kuzWcH60GWufVndsHKeCDPmKskBK0+G6NJ5fEwWk6ZVF22QjsGaIbxZahVor4ztA
AjQUnYABY+yaYFKiUOk126B+iWLzvtZN88ZiG/tfolOZ32ULUDRsYZMXVJIRkLuD
zLWT9jqhdpYjNVEXF6YkbGSvfxulA/tnOVfR7CjKGwceVEL07eUOwNBw8DWqxj3Y
cI+3WGEvP3Lqs4wGX8NGDaFDfs4Lu05WJoprj/kDPIf5E7z/rIx9BEamdgxZp7TD
wPUET7D2zw3nPmLdOdSZ8QDJ+knGrS6pTqyemhQdIgn28ZlPBFkTjAW0HGWQN0v8
2znNynYiBFmP5yJfgPfsFO7RoZVtNahB/CajW18uiFRwe0RNR8pXlv2i5cnv/B2r
24evZGchLm4cmQyJfWVv2vgBlIcheKASwfagp0w56tpGsp15Y4oDJjtTI1vzTZDa
+PgtYqvlvRsp0hgWo0JGro8GvWhGk+pzCa1Q1d1xu6d5hd0j9k9BzjaOk9pBcIeM
MhIp1q+Hu1purqka5F/HbA/r4XvW8z383B66SR7zG2/sHqHOqAbchWarMuh5WK+D
7OvMNGF6VnoIzOybHoZiu85z13ZbehjiofPApakJ5GN6yMDuD0+NCt+IqMoWyvy4
CBgbF4IY54c9xeNdYF28VU80F1div8vPcOWSmhjuwlB3Akn27nSmOgOWBaIVRA6m
7niWcHZE9irF8W3Mby8EndmIwPJOvq8F+qq7gcE6ngUNiBSHNf8Kft/Nwm/1XAmY
Ay586GKomIrXTHWCRoZoWrWThKElVegq4n+gOBvPGKD7z80dEdwY0OxXkzBMiSr+
Igg63yhlcnIwKixTK7iTSaS5Af7d0B0C8vNs3WnZB3oX2FapZhOWWlahU4k1rpwk
nb9MRk2DWo6wXyPp3YAgToIwv2EEMf5dmwods8Br1jmQQ2yAesLVJn2dKEFoGGbr
JfUETiRUy/vAz3KX4egUH1GpxXM+zrjW1FkJqd8blxzwMosJLvcFvNc75EhpuNox
UqAo+dtXxi9TtVuU6KKaLJDzdpKoMfncMWI89d6R13GV/JPXDpyt9pGXb0A8X/io
I9BLEJEJdvMQv9lOdZGilwss1MWvKyz1M1VnsUybccmurWQV/kobqoCl53WeC4L6
a0K6RPVXT91BHUnNudLrJAqWlKn8HJIz2IaTP+6oMI4fIkAZBdCA6IyujHDyTOSH
lzh8ACXQ+nUYS/XzIFP01w06gtZlSOLA+3gL847pOSgQxDMtLL9xPS7g7eQ8oOym
FILWtPGo2ddfHtVDO6SfyN0atljtO47AiyEJUpdD7ka0GLLbonY9IGdGkWo07BK8
/v2O24VTXanVPYUl82aDqr7aHvgy4Ww6aDV7vlVsFJ2jZjpundz9X8N8d9EVhWKJ
rC3fCym3qHhJYgwEIBTTFf/EgageETkQDgElpHQNE3VI2hS8tF+oFykFWt8xPCYE
lllMJd/YN41jgp0qDNe0Gb4IUhiW1yvoT9POnZzrTsaCUq3cNyUqibN5qWnlJ0eB
7sYr+11stJH8Fy706koyBPY+CeADXB/VD5t+Wrd55+ioYL5b50PZbivF2ibLgHrT
m1CqZkESw/b8/jkex/s2PnL823jgAy17XIpR0JcltbQ8Num5+BtjUEoQCm8x3xF4
10QLL4Um5dxLM4mrutZ7RcNIw++X1rpOsNXaojMRPjlVoYpZP2vgjNO0E8zRgZXi
A3XveIXVnlNoxGEywbeCKOaReWajyruPVED8i8a5EaxXiW6ECyXVjPxZZLbaSb5H
R8MkfpwaynNx7xASVa/u/VaA6Ms51MZg4idK9sUHX9xc7T2TMJc0gbzRcZGPHHTk
J777UBKQTLkWvSXf8m/la9RzSZ+7WxBg3PK2ZCLP553f5tO0ZRgd5n4g0nUn6ThV
FYEvdyVnTM2CsxIGsrlAA5YwhLBURbCumrNem53hFEf0rNTPZdbY5ISo+qruL0XH
doNJLqhpFTSFZT+hCnodRr+Y+aShyjAiBkNzYMPqu7AN+3DMRMs/kA9ZfiB1XJoZ
+IVmvYxv7W8cDCMBuue2OlE8d9VjNCGA8t9H/AgR1Gb4Jj2j2UdXidTGmmsNtsuV
nsMHiKqWb0D8pOTAzjuPN9LDRyenQN22zhEInAwUxFdtPGiK6MsG29P99ije6gjM
e5NGlll/FEigiONKsN8J6v8EnlIvBa7L3p2GomzMdUAKaeAci+GMT0KKDkTMq6/7
suP5/YhLMF1JBRBNYFVCdB9eHKjYsptE6VZs7Ppza31FOXY3eZgmmAvFQNeFGz61
QCf8YLOlLP9F7HwquQ/047xI0T8pd7t0qa9LhRlL9yfthrna1X0VgNPK3sTeXQRq
uAB9UR2AliRjkSMX8GhUaaI7Ik6WmERBPgW3Ji5nmPlCs67aMRg98fj5hYt7Hmse
JIjTxs7nq7cE8aKgztRczDhPExd+X0xYBJ41eJiiAb1Q8p6MP+1fS1XOnNpRAr9V
JmAFApe2XV8Bc3VJYtAmDGXT1eA/Ehv78/XHBjgVfmFG8St+hiHKhIYV3EgRS9cE
GdJMOVo92xnNDQsWsfV0hQve7B8+hxO9hq1cq1abXsDmH+YJPgQBCpffBy7Y1L90
dL4R3M4pO1URvGQPrWlUxhXo4ftzA2QoAtPRS9B558kxwIDLMqPRabQPuflQ3tuR
uTcrdtTs6vYCXANwAny/YwUcBr+aO7W/rTP5UwcOu6soawgCp7EhcH627X40BScw
90GSu0SeSuth4wFEKXG+Gu/9VFScsTSuAp0c3aU0slLPwX5JpLS6ETz9enWa3nBr
TZVe58+1nFlMnE/jOjltV7LyHVwlh9IpB0XBWcVP19wC+b9/4/QxI1NZi/+7zqZB
gSzaNdUhXSHAzkdPzWNxfO90SIEtlXUHRUUkJKlqJ/NQRR+tsngDpTzZWOXAeQJy
Ub28XDZ+wNxA3BSHJShdK06h2W/rli+YgPORSYywTY+5vO+gQvymjUZjQp6b30gN
M5db0QK5Yd9p9X3cRaGROY3Ljx8lIaVfQq54ht8B66leQs9sCtU3zV8IqdBq0kpx
HmEwq0DdtfO877Ez53PzFutn3ZAn8kq0SEXwXsf62sCLI1pF3ogvMWMIDr3XyizH
OT4ocGoexQc6Z290tFJmaWCaq1OuCc74Vibb2uSZjiCcuUx52CCHNLBHNchXSXSF
b9t/0iYUmJxDJs2SincN9kpp+q17s2IRxOHoPlJEZ9wo4GtXmk7tfOf5zYeiIfUi
1mhNR43ey0+jsw/K+llciEo/+ZcxCxkiX//1o4FQvh2tWSrjus8FmCANwYoyEXbL
PYHZZ/mD/MlfL8YspanljoQ+rjNCGgSrDcZp7iBi8nP4NAjZuiv5mrkoTak7EEkE
UPfxoyOq+37ddKS8dg0R/EP/P7mVAUzPVm+FSkse29z7z118W9Ux0dK8SMizr43n
ikXKoY1F1qDD85q8jTASi5CDZuU283eNrgczwsngOwWwwZTWDUmzdc0G3764FG3n
4SuuDY18Ue37xohKtKUG+PIZ4tdRHZvZLNxwJHFm8e/Vqa1JvOFrAOclyqqVuDXW
CxQb6p8LiO9Wbbc4BHCpJDF/x7+5t+Wwpiz76ok1L5QMNmqG7Q0x/UZ9587bnqFE
zslef1bvO6CGpJxI5OkQ5hd/npx60cMlcAnQ8CoARMo0R9nYaCnC1TgfDvmKQqV9
zIt+Yl4hd647mOA3X8MBCDV3agU13pQ3eSYb18bAeKQu0q0bdERfeX27JitG75Dl
hym14fn1RY4UC4ueD4Nqlso9yDJzkAw6GjMW/96KzoGBpm49Qf/l9e5f0TwY5xq+
dLiZMdK0xbqfiQXK7miMgy4x3+uq0N0Y6gZYBEs3YwqnjbAIrvWDeto8Q7nY9UYP
MQgp4JAS8DeqeTZOLAY0voNuliibftWW9KxJCu5R584T4Fn1FwXSGQy0Wz1i8fsR
pS/m1lsvgbrj6acNqrEwJ2WyWgE1IFhRBanWUEslKGEePAbkkjs90rVHhnzVMkNL
gHSfhURRGWsSzhZVIOPJs74+YRgxRVBlWFQ75L11gPzXNS3UEzZEE+sfvk8C4ljo
0GIKlm0Wj8RWnKx80Vb3MFN84Zv4nZjFR9g+D2pnMhN6GKA7Ok1W7ow8Q+JRUje9
SGIlk/VgZlyZkwU1W+/xOPgNjnaitByxYRqgHowHJIwOYn5c7hFwm6aWOHE0JN1x
gcJcyAIX56pFJD1M+XKmQ6E3ePr+X+yF+KiHENGWvS2VInha6wk5YRsC1pTAGeyC
zc09KjUZCtz4ZdtgJXwW45r7pCaKUeDHHr9kcPhMTzP+i2EhATeWV2k3YZJdPgkJ
lByndBZo8eLnAMeA9IL6mCf9ixD864YOH9iHhuPFBG3v227+KN3Jah2h3ZTXZcCV
z7FhT9AfbCbPyqn5IL8lt9fDIFYkSWLEYdFT+L7Que1qJIQcQnnpgWWtjof21LHk
p7USg04MBGAhosiw1RI1BefoTzvIrfQnyHh8qYPaxL6rfqEM558xcvB1ZZWfTw0Y
O2kwb55YP1dOPG+WYN/yJ5vEWuAeZTVbokpjr3XTi3TSxDmgafNDx2uvCQWE5Bjv
O+aMbbb+z8oGLA8Labz8gilJKlqqMu/YeHHG0dE/rn34YTcHqYSZAUazLH0ij5kX
1FA6Noj46bwst045Et+4tObgOHlVxjWoKWLP9n1AGIQ1UXm7WjUo93V1RZpBua+O
7FJZy03xUJzWUBC2n4fqBFOhl5CL8/yoxehTpe4nroj6xDIRJSz65iuG/jOvBG0F
AAo2ZgNOIPIECXbzmIXIzWnyPvnGNyz4K7f5HLb2oYEsALc/iXlq91UvLwo6iQUD
F1/yu1mtjQO9gJxG4ABXtcMcOdtlm8BPXTdQ4EInFMC1twATgGuPKQeLmk6ZePd2
J3/wy9+J0JqYkTlhx6lBAosZH9iEP7B+d4Q8fikvPzrXSx8qBaQu461s77oIBV3/
5sgodcx+CYY4eVuG608n/0i2uZk4HEdAfj+N3owNm9M6Vc1hRytCAOG90jqvU5+b
35pX8g/3Jmv5rI/8ihiOci+CXmuHM2MBcPsu9q4afvc4U8xa7BpVrBD9Ngpedh9r
wNARpWq0ujcNVLbHFavF6Cm/pn/uFs3iNsCjU2GMeAJFjDSwztm8dQOHB7SI+JDD
zM/KS0Pzi0vz7TGG4CssLvh1YXYyQJYvI1C03ynVpHyzYJlkzPMJErgccBVqx2Zk
ce2vvB1PERNp2yT8Kslsrr1PETQ/lDvctbinAoOI6zprzuI/5//zzfWa94/LIqAz
UgjYXxG+TaEhpiXKgIguHKDTPbf39SXtbhy0cCaaSKr9KBhwGrKSaXBvgdeo344y
HqVBhUzfK05xmrgEXpqhwex5GSCqks8K0pnUORWvpg9p0ZxKrFocC1xETX+YyZr8
Z8PXphGTAC4Nj/tODbC+ycqTdp1uciincjJhLB6ORltp0bsl6oZ0LLKNxN3zDile
VSJomULrLrs1gcxqasF3OVD7qisChzCGCcvGgmH07gsKrEZnFoGwBF4pV6roHbdj
x3uRcOEeZ/NJizArAqf29eXJ+vglLTbENYlJ+gWJRi06tIz6/QrG6SHJnq1yPWTo
KLN4mCYb4PSt9xJIGGJaiPXDJMP2Ou/+gvYD0GgxaSwcoz/M6xLjoN4sl1YgzG8W
PNSq7JK9nmj1UA+tgLjgeL/FgWAumJNxlosKhYaCBAzmQfP0NoOZ9XOvVkeeivKG
0PHt8Vo2Lcu0CHnvew7YDqM2hZfyzjvMbYuzhnzm94XSsp1s0snWpMMI0cY1UTOu
YUSpc73icjM9WtWLdPRN9qK+iLtyVZENPHxcKuQYD+BmQf2+6YkBlJGd1JikVgfF
QNd6Ug+gNOWiedwxI8RV4mAYQGtWJs2gehz0Dob5KYZtWnHwjmew/GrwoUl2Obp+
sJkaGjwgqsIdIhVF8ygeHBmsTRpe9DyVp9ABpYLYVzl+AecHpFUZR2QU5LxkorhA
QqHnYwdk6KeeViKibK5ur9Jw097r06LwsMEf2ymluEYDJkIx5TjydAdHVnrTP/gG
IQwTz6/HzN3nxL0ijfPiWadzma3XTfkv9wGA3jpReg1i1VCOX9+r6UYUUwz6/zBT
Qkqt6X+CUI8298mq8zBSXCow8vNhYVpqlE2rfctYQ5TwJAAwIW+h5TyyEWb8/jxj
flAu1IbbwRfE8EoQe/UIVlOiyV9oNAhwaGYZn7utjGHnZxl5F6XcEMW9wfuzrQmJ
ickWUKbglzuyQMe5m1mfZ56Yd4A1NzOOWh2/WlNGP4Do94tClYucl6YiTxqLbTuC
hN00pjMEutlWDzy0vcpmhC+lhtqSWZAD/XcSDJFFbLCDx3q3XHAV5GYFJJJk270U
bbMJF3H5c9cx/b/Eo26B5+Y/JjdtzbF6vVkNi5qPd6YS9VRDCe9WjitaAQTCoHoY
i7X10V8bwb2AZVfCPTRsrR+/+caQ8XHmo3yeZA6O4y5FbvO1JD9CkeHw+0/H4Uu6
Yb4FOChPWtE/jkrynZrHaMQ2EsrQkP1FV/u/8OglQKNqTMEm7gpWPuWOMUsSnKP5
2sm5lh7IjCCZsfswROWG+ze3lhuDZdFbcYqHqYRWAn3sMNtfsiMnWS6a8AmhGZ5z
Tl7/yJot8/EIVucq2Zo3UzlFOQUvv1qK1JMw4M09l7buGckXMHQeWybyImUxnqMb
z1ltEHmYspLiNo4T27u7TWjnaogv99FbjOXiRRkJYtgNWVKk68si4TW04Yh99k+k
M72n/WN8qThlF1w8lxejXXaCncsCmapAOM6UwOz56A/kNGfTNGR1sCb2da+TBYeD
1/HuDbrC6AS2RhQ2LPKhm//K4aWRMiQrlkR/ujZPlkCSzd+vTLpTJrOBANdf2XkO
PDwTedlX6SBpUsi2JBj+H+PIND3EB1gCKHH8KaTh+c2uWxNsShpP1R3lb0ikntNa
2kFVzRRG4Tc4Zacay0wszbwgL++JFGO+E5+ky2oRAW1PlG3MuHMw8oyA6pfwZu6a
hDAnTteJjqBXwr4fWR75khs53GQUe5y01qyTlLOrBzwfrejdvGAMa7uJNSr5zy7B
eVVo/yWn8WGIv62i+Hq0HZu7qjdeLnq1VPjmxBNbtAqoYh3n3+zTpzrTy7vRWMvy
OUkikElFRH3jtATk7BvGKZJpWFc8EwASa6QpIqC28CkfJ1311e8vR09MiDuBr4ay
mCjfbHwMqnpPvi1aE7Z81AAsNa8u8nMcrQEzautazqL/Y/LNkEBAlaeeqkbFI2Yi
3ba4EMdEyDuWHf5c2cIt+0UL5ulxcWqrAXNTZFHvs5jKhJFIHcXCsoUMTQabyaCy
GlqFfDfPz6pRCPhnCsr7Q6dm0WenNWBoZUN6WBTdQ2dUG+h9fHGfHz/Fp04ZEfrm
MFkJuvdswjAmGiX5qCCN6M5SCmTtGNNUv4vpzsJxlEOVXwgmuYm8gjKdgjAbq8pT
GK4lpQ8s/dEXhXWI0NIoLToCEd9MWC+SBh99PFkfpqo85zePblVKco7VhEFGVeF6
X1+W6/sIcIxZuve6wk9uKEfGL+YDj1xI1MXt0rSb1VhDIlNvego8lGJ863aSIXt7
ibiurJ1P9cWAGHE7csIE5Y+UBLUiRZCHr7wLPk32jJBlv8qoKplds1HqMsBdsvDP
lRMvabbZpBykOU/PfU99SorTL2YTCC0bigNNTFuvJlryrvCLVcZYHchS/fxr7koY
fwihyME4lLICHb4LmzYhsdip03jECmfd9SiJHZ8KLw101JE0jednRsYbg5bhLWvC
BODn6dXMTN3fCTTIyOtKLhAApc3BP3vr8ePWxT5xtNpoHLh+uEVJz+HzXWFfTa9a
f7tlET5um8wQniQhqjSayHn+jCaluGqGQ927r57lC1d6wp1eqwvTFrzaBWBa0KlM
1qk93XeKR/MvFVctSyMQHyyzSPhPZ6+HiwDR4NSMs5SbqXq92YEK/cmbrT8we+Ci
tPI24qNRAphj0XXpwuj02s2C5WCMAFjKm1iKyZASorJkFejTJL/9TOB6mCkjbzHQ
GHnRhYYdCa5QEXmoHHxIVS5DhzeC3XO1KRikoyfRyprKEQVcUPA1ySJpLkcKQ16f
sGsPdQMLb/X1EOVvRNLCcxt7yXfdmBLVAX/BrLCUWu8mWmdDX6SrDNNAXBv4q2b7
VfNlblRafaySbNZjh/f+KAOpdpapDgHaD4ISFAPNaJ42+hMwvkq2JmiZa6B68h0N
VCZWBLVuuK6aSziRaLcJ4iojRAJsf1uUqIhcqAkxvadAt50qmoeOQZ5a+/M0FZGH
5JODG62KGrN+uH9THo1KUoGBgAIJV1iy7zwMyWFdIh/AiWN1fDvfESly6vvG8SkC
MNjTJa+5XppJQ6fjw/Do+3miyikiMsd3tas0dND1Sc6BooucAA2bZLzNnZefQ459
7eJQLS4Rw38r4s4Zd0vwrVFR1QTbKVkEgCvouKwFX/jUnOcid+EwGJELrLUNvnoi
52BppC1z2luowlywj6261oaaxIVIwUehOISWLPOh5TTw0lw/N5Vk/blDoR437IQk
Jiiqr7uXjbZQZVsr0uS4jddSysx7SEv9DrXhZdMauS5I4I9khOXPalrhIXq70DL3
zO74E9Ec/vQy3rDKpJTn8qE483ny/v4BqnOspx3CZzxUjd7q+ULD27+fVvPQE39m
BihLTHIICt6k9r8tYrm7UBoLREf8G+sQ9hdrj+hF1oIN7uHPW9iovmnZoZApEZRa
pdHUzOEwzsWf0XEr1RMwbxSZv8g0YMslIKFrw87BViygp0yIFMAlIwHC/crc3u5D
9s2C01lMWV2fJBXAfAxp5fDVOvMJsF9wd6hqiYU52lvfWQJlxCDSPe1kxIeoweKf
j1yLomTjO9vDxfrmp+Q5D0RAHzW2vF9O5+CEpUCsgVOw5gBPg2lj1lE9qc0qJBXv
Kx3H7nOZX0dvNHJ8m3iImfYTnijkvTsRyn4WPUVV4i+NlvqLJwklrOgI7UlVzOsL
sm2ipEsP6Ck9TE7ZdgewFJ5nPLiAdXzgF0AHPtscLKMKp+ET71jTSChKhWEzEzkf
3y6hJeA3tOhig4hGRypysZaC0vbkzFxNAbfVNThh5fWY5K5BfYk/xVuiII7YcJj9
rUpgytLxXtS8JtmliBANdTG6cFWdrzMQMgUrus/6Fj6bErWp+iBspmKiA364vimT
xdYQnqmKzeFhlV2z4MdcgvhPbXOY1aWvKtJUHe2DUH8++9hC7D6Z+KeIs4jqmuQv
9SNd62s1CVqmPLhGMpPS/AQslz56pTxpOwUdhJJCUMmEzY3lyhFon7bP8MCilX+M
/O7sqfqiEw+xaBUr78XKPY0wIUwI2ypUOX3zSCcos1oKozcaAUxVMBKrhwlAHwGe
69rUmmqcUycBAREdb9wOtzNhFgXZZ8F+RrRlxRYOMoz/DkCaahAvmoo6n2qqiuTO
2W1MZm8dGTd4vPq/DHwP3iurfBvy8i9Nus4z7htcGYvjhQYidWBxAIA47JY8yos8
XWcUHlZXYhjOk+7fysFjyCdq4crUlLx+IuzUBB8D1Ge9kFhKSIGv+UoyVr+bk7PP
rCMbGe7+oxC+tKu9pfTubK1hmmgEB+T2QQSTsykCobGDkBOyMZgGBGFIekTJ/qeR
ie3ndPHGCClW6LxxLoNRWG+jXLatuxhiiHYlhhQd94GeZZFFsA1ZCWZ2qhEfw8iH
vzTl7MbsXlAN8kSpYgctBI7l9jFXeip2sZe6C0k/7w2uHlxuGJbt72wGzA35V8RP
E1D+duS44qtWXhp9jO4yg4I0aZGdXi+PPfTEZgVvhnaF9DzgUnkXSYp7kvu03VG5
CYHfyhoSJOR9o1dDpCAoWPQlWxqj5IFH+SH/XK7tzmcchU5hAe7kDCaeMBUSUoD/
bSlmXG6JLCnoMqBDNZ6tgsTzzfMeVuFY0pfgT2Vzb3C3dwHjOUQSiasQ73Dysmur
eyuckq6zHw8jwzaY8PZByM7ijAMRG79QjSGxSxhAXj1WSMKyv956kcKa2IB3SNkf
dw1o9/By/P6mZSlEj4IkKfxLgY8DP2xFZV1/Uca+vuo8ThFWoozLYZSXcSsdcLoy
BH44ELPXs1OUw9+aRjuESyljEXoo6+NlZ2drlxZJV068B5GdQSIblHaNlgPKOimk
+Yg90EGDV1Nyxq2rAiA2m0NwlRPnkfPQzmsEra0mDNQGfN/QNM1R1aYwYtY4yxWs
tSEUN0H99A6YlyQCm/koMi/7kSOefbrX5whPrPqKrU5BaB9D8l8jBdQFSbfFmxFX
K3MHBqpcVbtiXFhE/vCkX0N0z9RFHttiLWPmB0YZT0Acmvd2F6F0/oIm56tU9Kqx
+aZ55+qa9MeulSYx0plcgsz5tP+28I3zF+abNrM8WDHuIaGnFJauq+DR9/1R8oDU
IbG1hl3yi4fggedTJu2UizhYBdBr5XupTlrAFTgge9JAD/PIH7nApgCSxQpVLswp
rRU/DnD1pD2GSRjjyE5T1yyXKSyZh8Uzo2ST0sE1+1rsLM18bIxe5Yl2f7K4u46Z
mJZWlFqZ87o1oD+pl4xHGLDI+Euq4ZqOkNZ9UODOQDZNuCmvlzliQam73V8Bw3mo
v7ImBJCs5l368E8vnwIG0Y82Bq2Hlj0LJmNU6EUNhKuijJGZ0e2Xz2GVGoJ1CDEN
IQMbEdqbAttuLHum0BP4gzU3uoIHpP8F3LK+bAlnNTdJBUhpmtFVzyJsDFRUZjsy
qzmiawhz/5XWIAn0o98c17cXWjF2bzchnECb9Wdh2g3/oZ4ZdnuieP9Qp3xTUIdv
cWXvE07xglQUk7I5F2IT13/B0oIFBUwqbfb6TtNH+bPkLGdIgPTK1WSjsxVrbzz4
wswV38Q7cDu7gCYhHj33BLK0e9fpcdw2D37ZpMNyONhNkvclwG0l0KS1TF4WGBl2
9QNkLcbJ7sxBaSaRq4xNGJFLlpYdnq1YphME/Eb9p952VQBdJ6pLXKkq/M+K6DFZ
lRm9cf+KzT6ZHZNYR+gq9f48pktaWl4rp8sErDVe78OT95zStFNRH0P1yZObatgC
jHK/V0N3YHfbP2FOBveQwhRjdTp+n7hPpOq4MCFcrLqaPlYgl+Qy/YLLpulf2FNL
hJm/iNCd/NYdUX15L+MLKu64MGW0AqDTqA3e3ZBpcQqtuTvtkMPMWXz287Kn4gy+
Gp0TKNlgKcca8w4m4UeKu06eX7sexnN8vOeIQFkO0rBMVjgaBPsI3pwvLPr9UM2p
WYC5u1meQpwORILSDK99VImpOVWMHFypXm0rR0WkQ2b2jln9xTmfWXQVqMmbsCK+
0RmgwK+Jze3gi6FzjjCCYL1aqEbLwJuvIUucm/+WS3trDKCIub4VYJeBc2QmETCY
KiN1gjlRPd+fzTqsMhtu7PmqOwUee8+x09/bMesJYeOA+uLazMTjMfW3wK+IdBov
0wcFI1URRJy/mi0CCK4WluRejW9nwNQxBdklO8EE5dHc7dmmAlsoagx3ATjYe6HY
qtShmGfHUFQn5YiMcnO/C9h7JdaDiSc1Qtb5eGTJRLo7BZNOqKXnvlxBeLL/kcbt
Zc670WjnS8pzCnaqdARbx5YaKwhKrQ51lCsyLNR5dI4oGovlX9zwMVWyB8C0aNXa
E1CBBSantf+C90J2O3aYqlBkSsIHr5vk6CyiM5+62rf5EE8/K5y99xFJjsgaO0MB
wnv1jhvTdXKf15ztyZoFm3fiieLWZPjFZaQzIOUKuqX3xIenEBy0z9EiAGzT8vsH
7qVroXFhIQ6Q2yp6ixcSPdJv8XdSeMfPqC65KjZ3xb+oHXzPqF0MqU00AKO8Qebr
Do1OuxJR2WirsFacZwpVPK0mO+GF0r1Gc5pmR1KEIw7FPkH2ynAjN9Ctrb/M/J90
PZ1vkNxjDgJvNFttRiKv5qgWdaoTRABgjR/z/+x8CvBx9QKGycOXheKCe0/Oe+/X
qRCFZUZc0nm69kx7BvcVh+KVlvAWrqedgLq7w78USkKdQOMJVS1gzi6mXBvNa2Tb
Vu2zyWWQrHaCo5k0WDRxsh+/EA4NoyhGN4+ng3aaj96dskS14Ye49NnOPdQLuzZL
EawZSxLyfIsATI82CmiK266i1whTnBhSC6VF3FMm7l0tECqlH0bxV+daeGBpn74q
0jJeff5lthc3O6IrI8i4fRtqyhMWhBWloDowSM7weqEQzAT1GBfQREP0pn9g11vi
qJsb25bIujjHStvkYHjQtBi3+Bj8+hhljf1aqFpRZY/8fGUcwhIIUuHQMEFUfatK
t2q39eMLg/07TjLNBU/jgG/9LEhcSC8zu2Kw7nFisS1kRP/y5u3w9PeLj6sVenFn
96wHWKHfXuNeiz6R7HVlwLP5cHMVi3ZemmNDuONm5ScopscGsBIfbb3FvnpRA2Sv
GqN15GHr0rrL5mQjV8tltIETFH5H4wuUtyBmT/kmu50Mnz+g7tbbQQyI/as84zmY
K6kpLDlUAgE6fNUNc+F+Ac86iLbkPJIXYzdB8OOWeDuc/4NhPC4roDs+TglTO/N2
pcvcMAzjJrIzWl31oID4lW+D40lHBn4gK0mqMnIRdWdPaD6oRiJ7Lpj6gchNqToQ
qDcsB/FW9IsYQ7SM09q7gXMD2kzi8HbBWj93hL/GbKpq0WfvwyQ16CnDTAm82Ld2
OUHqjURVDFTSmSV+ukcml5X6N16a9smckWYjrhGDwN9ZPcwwh2TMJxdcXVGnXaeY
HvqhfmxniHXwzZvI6hTEcXtLREZqGABnQmEh286jX2zWGw7zXaXkD8K4zW5/XTox
KMlmr6nLQvKGsn84b8KVH3KM97g6v1nZGO20SR1Xw/lU98wO9pFPBhkXDjHN4PtS
NrjAxWFHTCqGeLTyNiAnLYPMjoraijgDg3l2f4ziYFjPuvfNocI7vHI1yOCPVm3M
oWDIxxQy0rw2rrPHzz9KZ9sEf/JZRgZLp9raIpu+UtrH8oa2JwBhmab8hiuuM+VA
HazHJsLut7+IIk1WEfAZTvJ/vkvnkC46aJn9ynWbUNIehsYZ/KWBxxO8RWwcURm+
BJy7yEAObAM+56NFdfJCOa5HREpC1LPoiwKZRla68M3XUO3gUonnYjHm/WfpS1GL
7Q/5b6Q401XrFBtg4hNL830b9RIe256LjpJ0XjIf5KRcSHthUX7peQHcldT1edtZ
y4J8E+AE6VCBcTBSPu/vUBOZIE0v3M8112YRYEeQgmlXJwWs+gc/MCJotmo3x5Co
h5sBvQ72XV5AaPh+8zaRNsnJQm9T/sSotnBQAs6fQsri+QK5Jbgo3oaX4zZLlkp4
B2NZEiqNEZNWiiq+rTR0Uj5VhgmRqpp1DgsXcXaB3gVkdrJsQT6dDPZlXLErYEmN
G0WBhfqoQnw1NJEP+K1RMAE3tLhH5YaNoJlyoZw01C5u/WGNUJB3QMDJRZyDMzjI
QXlyLel/BvPq1RqoT5aq3Oqt77HraNrn+eZ8EZU6MddDbPpWQr1dT/o/ls3NRe38
+SgVYFMp6dE8FYkMkiNhGFPXgIN980owj2NWmBLJoH9SxDyEoU+scbZCPET+7Ndp
B47orezFHCNYXtyd38Et2BrrhHaS96DTHTsfeQy/MCIlQfFaM36UzdBKuaWiqRfq
2JbuGHd6eXPqCg4bP28SGIIJdYidqUNT7rvGuQaAzAXksTqV3Fl0n1XSBz79FurF
UgsE86nIpq1yMLWinaSnLMcli6T3wAwXkO1VR+3wXVdWk8KZ1TGkcMvQ0SdZiehG
opS/n8+cjVIjXx4OcpHZInI3Zh+4qH2fdsDQ47Jt/c0EPzbo1D2y5Ejj4o7zhtP7
xVo35T5D0XcI6q2KqJkuf1AsQr3peFq++XEnxYr+3o4CVjy7ZcMco/kIJTCYEfn6
okAa+VyNo8YhsIC3ZG3I8IYcjMjOyiEvHgqgE5k24bp/yknFny/CAMTjrNmDhoGn
16rpXjLNbE60Q3nMeYOCECj+vxPYwQHF/zTsqLmuSLCgc8XN/YYf2BFrnS/sN17w
GglfhdImDbqk8UZaIfb/kGjYcsgoX49qcdaKZ0fQ1HmRhzwJDc55xDBlTYjrj+dc
ZgwkvUao7JSiqsYmVcwqeHGHTSrlS/Ode+antZlul2bTxXSKhfJ0gGzqPPjAJEFJ
m3xlUvDZZBnwtOhXV8MykcRqgNHNwR/MNWPcEh7bJRpnCSCC0N/JgLtsF6n9zCDQ
RFsLxpv0cuqynyENkr0NfWO0nSQVJUURVLf02W6fVfQ1bQ8T0ecaKZxbSP3ZwoV8
55sR71/RYzi0NABkewk5/KLq6UOfIDsYyPeaLrOWL51EP4DzG+lxh8dfbyMdCnG6
X9ymG+F4vS8NzLSysBM/Y72SK1qNHbc5CG/KbJGzMCejf0Aw3yfQNzmXw27famdN
owZ8rUuaE4+xjoyolaNCqPcaKDiHTkLSxMzhBDMBHxscLaWP0oZPRw3ZVEF25Pme
imQVIBC05PXvgGyE4n5XPy9tH50IdYiOtJTQqx3pYWXjN+LCchc0MQEajwV12uby
C9W325vCtzv3buS5HDW1Q76gHwFB3UlnLihE5yjp1sRh8jgM3bhZvtqPXG8uCClK
T8J59W10DGMTd8+tjEEOc+g8TAQu9wJWAfK1pkdzj2cAD61ZW3oYpvf/yjjky40c
NbRdPXB0JOdOW0DUY0xTFc6pZtfg8130rmjsGnO5EtMbPvUmXWJ2GV/AazLoqhY+
X7Vwi/T/ha7EpBMHWi/YUoqoqdngT0fYakBFLt9K2a2DsxfByKgfh1Wgjk/ZXQBR
LSNDh3IbNu0tSpQwyZbl/K96jubJv4d78x8qM16xVr2vhIrvG6Ya94wm9ZyYFT6N
zlPbvrAR2wGBnchfjJF3ACh4pdkO3fpt9q8mtJ+zrHigEc0E1vz0JwfRO4oFVHEP
J216JD3OvhJdB+HxfvE1mcs1Xl2ejTH0eursTvQw8Ubd70Y5l93ky/a1A5ccfw54
ick2alhMWRHCtw5RR+gVgJiAQAj1irWvGVNDf3+AV5Sksmgxv6TarOOBU7Z6qNMB
cAzHdiQN0T4WwZ0nCrxw8Sg7f3nYYOBqQrviDWH0klNAhjXk1+JkWQevy+wraKb/
lJc+p9PHl/8vHXYU3jQPIL46cXfkWJVQIOuwSYpyhdBYXsKnKjzB6pjG8GZ2fYp/
OePweFFCfKSe3uKCXHFL8JO6HC8g9X901q7BqSmUd6HUCPmLz/mnhf46JDUItw0x
dl9y9iMlpyZk1ChiIDXDk3LbnAIjoca0S9AlvdUkIW+lIPCJuYtBb40EYU8aCzbN
+8Qo3ZLDNlkCQ1Kiprm1zq1rHxlxEgiFfqG81DWVokUa7ZLQZ42XNGNSrVI3UwYb
JdOdEiay/z6XNXxpV8LgQeq+3OWwQEbaje1+vIZ4yhv7hAv4cGRNd6DSgsz8ASHZ
1b3tpPxPhZ1ctch1HUY1NNjfpX/pCn2Pvq2K+oKwes+DZjO6CubxIPFXVzJLPEaG
rAvW+s+bJJa+m0ZtFQb2FxdZBbdNwZaHnp3MpTIUgvKJXwiI1l2xDiV4upXUlHZE
oHqu2N+5LamzXDCq4nX+H+SO+9+d2jTTPjuP6Fk91LHPKXpO69gSVQLIhh6YlLRW
xhJ0j3FKZOy8KbKRiR+CyJ6ulS958wnnpE978LKVZFeYtf+oQ6RHiZuxh9K7LP9b
qYY/ZIN/JLpIdp/x+KX0/mWrPdpdOe4bkI3H3526D8NqATQqc5h0G22HV0AGnGNJ
BL7uFgEvIff8mbd7sUWq2ATwnpV/8R5s7hf2ZzJYXrjyS+T2MI4zlatZuw++l5Tt
Dm9gdPfPSK+igVpW8uNNvSj+G5IiunCyCUD6Tt+iT9e+szK3xQ3VH0cuAbRFSm1n
+hEBXlM/VecYN19jHvgy430WqFdJc7FprexUeMWnPm2Wn978hEyrC4lRlQNiim2V
NyzVXs7lUr3lDvRPg8gHzzaRWRrIDs1P51rBxSIc715aCT10WcOBcJ9vuaAs0RV5
dL1Slz3GjhJenRnBTarmx7OnHIr5eC9Pu5PBlIZRNTZ7t5k/wX9Cryc455d/lMIT
ZYaOvy19W+7LIm6cGB8fFCjAO0wbVMPb+ZKZHgDGdunkCZm+IYvk4n6cU+O0Hwkw
lkad7dLDEPZ1LJ2xdY+HQ3Dnr5+oV8gb6b+ZqwTNsj8Rz+8tdFM+npmMFXqlv32z
vJ33HhzT43bzq5dNyeQXD9uFcHCxFIggAT656AsH/V035/5aLxyZihHvaLXZNeEO
e7rbEvxheXrlM5MPgxxYVFC5II2mOYcUvG8OuzJDW0TII1+VDQ01RYy7cqoaunTV
YOBWEvuF+rdZVznUpq/k92krD8ErKXstXVH6hzu7f1BwHUJ0NyxlAyDOYaYB+mY2
jpNWTz4lih+OCvLG1Z/pwPUtYhFKdGuXCUZnLkQoRXcM2bJPvwHoeHLb576zLjF5
J+X1kBe8Hb5IvtqXG4kPbVZwy4FM4P3f6AF1Fz0ZN2s/A5mF1CKZZDoPhDhjGQQv
3F/E2x5MY7xLKvtLb1UE+hc64TnGUwyn5YeioYZeyzvDDPonNfQfxhnjOwtQ1QWr
uccxJU+0weYHuFqV/INN4CnWeunS44lQPSebjUgWCvDFqC79Z3M7GJHEJlFZCjXj
CS4ls0qTUOVDPkWPr0xNYr8LIxqbBJG9JLGAo17NYPQziR3xMfCi0iau9o5adaJH
hzeMe2Fav3J2BSvjGhAXEaa6gyJHO7pqYmXtn3ee+kyL1Lk35t5PjUYyvOykuyAh
lg7zw5l0NiBqA0sVV8NpBsrsO8a985TPBCFSVjwvyIp6LNxL0n2NdgDvfjmoBQsS
++KTOlouwB59nmqao3G8qOXCd0w8uKMn0dUeS1DbskgQniVi98W49Ej2fSL4iOGV
YzeCo1vhCj9OWpIPkHUQKYveF1D4gWmmjVnOgV7A1qcAI/3c0IAF4uMO0cKxBHXY
jAXflL5DDTZR7ARZvWE86BRq74sNWi43hJ4KHODVVxkFStmvdTOLl1xRYwZcvyUH
fCxeA1PCc0SUzyi5z2Hxpq8pZ8hvuqnr3483IqMrA8f77WvkS6dWu12y3dqSApj3
XRgLnEDqM7iE/cOJOxJvLTGn1SxnRz3o8HCK5LeNvMqzusqFZKiYcHioEt1yXIse
jpSMihelCkKLF6zVC6sE57A9iuotQ/S5YU3zsSWj3Qw5K/U9bsJMQpiATjNIT6DM
JKrwFOkypx0GkaXWXuKFe5LO6BYWV8nobzMPA+05VfuYqJjasFgL9V2u4UHvsden
x85x6jG+IqQ7uN5zwnn3zL1pIG1pyZBbfaQwlOGE86SLNYVShb8/3HsNrce8IPSZ
ov1Vfhmo1qED/3HT30Cr1z300/vTOFJZreBK3ZcJvlKjtKF43JeaU7cyvajegVI+
BrM/ukErAgfwcUlTEEFOwOsGTlLcfx6JxSQezf0QBrMeAKIuSd0Wg5mzQMbch/27
Mu1GFJppN0Xthjliwl1drRDTbtjrk224LmOhXy1Sp/LYfn2LTy8L4GeLWNLIwXkc
k0uOAYEwcQeLscJkGrplS7I3mqiiGwqVsnCD27xtbx/qePUs7dfqhfn7GVrTt9+o
iJqmEcJaPYGwn1tspsdu6vd/SdWZqtSSsVoKr2kjeWx7AG6TYmiPy8b17xUZC9Kw
LLx/ofFvWQa1MK/NHuNKffXO82gLBPGsyAKZne2k+RkkUeFHx5/djAZ0s3OFPHE2
YYu7pMmLQNjNfLx1fQTkWQe3aK1cUvYFd1C2ZEi0XylRoaQ5jzGi8KizlpuEOpBs
veWpPdlFhe6FfHqg3HODx8ccnH242HB8CRZIE5LOVzwtsAClhkH/AoXUVk1yUHwS
fdoXMOtrufJu6iWTKvH3bfmX0C4+3zROnXkU/2XuVQWAMY+hLez11UfBjpjbNqdX
q0ReE/njZCgbRgghtNae+9z6qxIA1tcAP36EMmsdOp4CkJWpoG+Dybwc+CIpxwmN
r/qDNSW6D00+bYkCw5kfM1RKmmv6ZVHV/h0wfepjjRMRLBAtpT5by+B5Ootu9Xv8
s27gIkfZqrWmOqdKR3VqXk0hRjYFSlS/nkFK0FzibNVdh55bT6D6XzrR0CM5DNr0
4iU3xKDHllZojGegPlE/Og1Ciu2hgLzxetTPe92fdcn9DVusLdTwWqyfg0MgDg39
JKFp1lC18T9bI95jcWgx/fI+EUsMWUmbnRnx1kbk1ZekPjeA5NzvpQVfzsX/JSpA
RIEfaTZufdJMLeT0TvfadwukRMPwsKDZcBHAIWWLq4NC7/2jlZjarDG/H7KPNMOL
YLOLh8AoW63jWn9u7CE8P4EQy5VYZr9RQVv26G+FwKa0vkcwzGg2gRzRajOoyrU8
s2V5Iz1Ro27O/QM8TWZXLHFb/oXRdADo+/oRLCgmwlP20d8uLmgftOa6K/HEZQXf
IIt1IHWM/Oa+/YwQVIuP59dYMoAXr+UYybqr1YlCT1Cr4sVwOzkRsFfQDZ/C3j/X
lHVKnzJxea28mfllzW16JfcC+nQYT+K1MPyZc/GnsD5M+CVN81yV+mwVZljvRs7l
4Cv+ZMrBMn13V7MnNMVs16N7l5cS7H5zlr6qsIPHbMQKzJD3COBGme58rok8twLZ
+kFpOaac5YAvQPCF7C9v9qgnFxtSWGCh6tnY2fUb6prIhZjSLFiLPkV/rXth4kKj
MhYR+hpV2siN2JYcQQXQUS4UoO84w/iHBcglai+BwkmMj5w/k4w0qv7hlnFF1hy8
UwUrWbVYmR1BSZiTawO8kfq65RW5kXIRe0dc1vJQbZ5YYpbnpBA313Q8NNMMhWHC
30eb7jVPFVr6q2AVOp6V4lRHsFmMKjgds6HDr+kqK2PJO2L8S+FZBY7GXEJubVt1
g3GqQKkkMGyCxtQbYllKlYjo+lcbjOcx0ZX79ONQ27rx13r4uNwE0L/EPd7WVnQz
wFncz8cFCDf+KK9igZPP2IQ6aEqdbS8r/U6sF5wazeJ1BkF+azJE9JFfx1VPs7TV
/ZmjyufFN+k4HlVMwKmMpmxlgEiMiWGrl/pT+fn1sHP94ltYjOmgapWK1fH6Rnqf
9xQT2Q5dZbYQkbA8E/pGe019tsuGiKxeEn3FrPbJBDLTuwcFEaphraveAtuOxAO0
koj+PnBRSYmtd6S+7zbmGhkBHBGoktsdbvMhGMik4sX+6w7j1x4EYSRw81b/5SFk
mOj8ABQkWiZQi7c8CoygApulTt58ojuH5qVW9iFgCSL17eZDe6x6Eo737BRMz//F
C8qe7lBG6El4iaSURd6XUwXXIl1GJkI9JASj6gttFi2+gg+uuxbK7lcHGLn8IuMc
5XrqScoBEfUwDLNRgkYzHrZs0fIfhrVMKJCgj3lMohdXAvCSceLMb0jKBNhhucqR
zu6rLgu94L1LMwTWkR/IK47zHlzoCcxGk4kpIDoJMYo484jOaD06iCHqwFD0366s
38JHLxt9Xq4jfUVZSyujT56DgzK8kcHF6jcWJTQ8rqEJlUovGKfnhlXnt3HeoVMe
CeJd4emIbOqKFqQ7yR4WAJy3oKVANeK5rKHngxJElR1K8R9/nMIZQ0A5Etpnk/eD
9uboer4mIPY8io1nugc6wjpIweUBzPhvbvBJ29CXg8+ifoBx5Vk8EGzNk7BVu1g5
sN2cYIBwO0nvA7jSYCIU6CqHD09tgIPbyNQhms/Pt62acYt0NWwu9qiFnktrsmDW
CnVv7HsqM1vl7KqBiRCbfFBaFv7OLhdc+InIlG4nezRIbst1NRxvwJ+laHt+KmPm
Jou+2pWApRZ7VB+2ZXRfk5JBUNdISk2ihvWQY0k0knyAs72EKfzSf/TXQtu4K8Xx
ZISfzfh8QpOz+qOEiyfAmrPvMdMqS/ez1kU53l0JGn5j6dKcI8B0XAjM8zQHtRdH
LloJzxhnFfzapjA1xM7V9PKr2OCzz9HRAcFfYIeg/BzIfTscD+4jeoCj9KNm3wch
W8GLUA4EoKpI+++Y+OtH58mTmbNFCevTkkR0VHjWFP3qVsDOBarMatwoVBBflisM
OwrFKDCgPpzxGX6uKi6vFhiTkLGIA9VewgTP1rxqmppVzCHj6SAIZV6OklYmZJZI
GnXmT80CMNoP3BDYzwi9Oaol5YYx6Hryk/YE1HlYsIxTARI541XT/QwuWG/rjGPP
c7NU2SvJ2yYuOmxNYNamxS8eO7w+dfxjz9IX0GjJ3yNoAQIg3e8L5RKvVERz0qqL
fkbpIyZNOvCuM7G5OhRzRr5PpPiiAdrLtx92fZ0kybv4Z0cmcrFx7ZBbYu4ZuHmF
XdSZIQ3ouYvVr2LFu92dmxao063ON3rogIaI4RW8udWwc1xGOIrb1QTzzEo9CYUy
zYdM3ZcIZFZ5g2n/dWvFKnStTYpn4HAqZ1P6tz2tqI29OhMdYGF5mlhlsTuZ3fve
YoGHWQLeYukzoPLnkKuhanBLgw/XZYyKmkZqunqiQSvKMmLD3mY3F88bB3tKRZtW
n/DONCOSzkv0idAbKOWuqU5t6eCTe8v2QyjDCbZ0tf8Xr2tHRTQhQ9NhWXWJce+5
71It4Tgj7Pd0gDM/3L5vk+Ab9CImq+slWTgqCn6T/xKDUHAOQRcK0Xgh3yJ9+F/l
1JM6oJ0FFxihq7Av+ddsR0Y2YooH9OzxqrrUI+duVy2iqbUrjhbqD4I05NgTsV4e
sGLWCcnPRJ3sITxiE/oi0a4g27OqWise/Vv7PFTDE9owgOwQYyda4CcwZwOiLmss
GzL25bffUO+U8nlyxbldE2nbIJqTv0AAXpSYpaNYmmlQy3h/S+fAs5EpiOVJvMDf
ZPn/Eep1KFGVm787RWjp5RvTQv774vRdx5ekGSDqi3LgnliMLs0ZlR+xT3VBpq5n
4ZJdyODFef0s7T4tYgNoLScbXvVwIc95q2pr3yD9u+qcuxcKbwRGTDS9HoQMyBl3
uvQ4BuOuIfQa+K3vmnmoTnLqD03tweRppsLgVsBBeJ84OgRyPzVTG3o7oRDuLxhr
H/dqjkMXhUTVBUd1ox9MnIoMtOAgDSLBpfmDpLoiAeuNVnbBLvZ/X+MQOxHBQqX+
Kt/bvE8StptKuCq9h6yFNTzDg3zZGVmgmePL3GbP8YJli1BjQoOKAfkZtUUX4cxh
KrRluzL8mVjIGqHh5T28aPUwFSBB9LH3F7enMAvos534If2/dHtZjzDCDl+O1Oci
G/SNooakjH6r8GaOziF9ZogHNTn8JbEIlxi3cr6uLNK1vZaDcshKHrtEi6IuZWjw
EU9igj0CItChsHzt1mGe7tUpZz/DiorYC26eDal4y524ptlKr646gc9sCXCA+uDs
o8F61HvModUJKOOuuvCiwFQOR/SMkPePZ212+Wn8QKbq5f9Z1tThCuL5etnb/DRb
wM4qiSF1D55dhKaEBc1JMhNN9ZFKxJ51NXr7PV7qP6jYKeXVTBXFsriK0z1v5xTf
f3UvXTN7on6F/xQTNWo6aTdGGDQvdn2goUVkf5zM8ykvsFrGcEZVl0TDVjTW0VC1
qNTwl+K9I3zPW9qvfa03vum9c0cKU/3obT7w/q17fs+vmraKNdLGqF5jrzfJjxiJ
SJG+mbBQffXdWGxKcpALsw1FhbMYIhrtpKSXvLI4O4aBPIyrPuuX6YpMcqHka49W
fuVosWedtbhg4L4T8W2kKT28C4r2lkupRjTFDLiY/vxQFT9rl4++WhMMOUqV2+2U
Cj+4dj864MrpyqAH5mLuuqWXyAoux6uMJEjRUOJLSmMcjWcWibTLORcGw1jd6gA5
PxWy7buyymfY6SnNCK6t/Ddeo6JpYviZTeN54FAT3CesrZ5VspdZNkPpUtgSUT7j
1WQnOyyRpIzjii1N/oCOf1QmNUoK/izvGG2BWhIYCyr8qcJBZPBaVqGCI3iNsZiw
JiLPfcr4CNTQpCefzBVjp0SPuHaqxDnM6HYRmz6AhS/fFHluGH0s/d77j5kB4b5C
80G7+Y95V65m3CA+TVrZeVBwlDBaBn0C352mFQeB0vrcB3sygf+9mwejfS6YApOc
cXDz2BqoL2GQtBpgTyPbRIJvPT4UqBJVkOnj/OKDSass6QNaVdQJTQreXf9w8xZj
yjUStJTD3tbeoRcq6OwaJ0NHpLlGaXwn1aMwu4Wa8dmhnz2HUUyaFF/L9Cdi/4PO
OmLEHtB6+aR6PEPo57xklmA1JibZ4i5bg5H6LzF/Xba9PXZolVtGT8RbDRn7kHYj
mTQXBpNoHlTC9vwEud1k+LUlVt66dygjntZJaI8KurVFZTUYQ2aPIhvv30HSRfEA
ufpw96SEZ+bkdvhHVTnS6ZDQeOPH+7S3+zc2q5sifzVImFBHJVw2vkhHCSZaOPBf
zMXbMC3dDzT30Cc92Jasc4umUBOoJPpeNGxusDo0a9O6vOYJgiHwOll8hPVZmEvR
Ivgp9/M+jcZAk2Cg6g6vEBpVa0IVhbEYriPA54YPWBBceYOjVvYrt3C1fC7ybWIZ
oxI+KzyCk1+GvUHxlVJZhmoAoWDupafOHyiUCGu12QAYhcBuGiSl72lZtSB7r9FR
apUTVQ1+WiYoiyCkXnc5BkZwVwvjTWeckjP8eutHYs8G85+ODd/D1909+YlIrJxG
F5OCiHMab4mqMdp7x3qnGWOd7JuTr0Ke9TcW4wECOVYxpRRM2GJezpaAviVEjth5
ZwvKd2o5P/h2rpkSNjebMK91eJW529O2VWqBASU813jjlsoRezah2LN/B41SYgmH
CD9QKohX16iFQApqbEffXl7FLljK3rXegc3IEGKVAbDv/vlJBPEUJSu8GTcHLQAX
qpmhQ75s9hwGr+byU1zR8F/HXDElqnrmqekDo12q7vGoI19DJgCFKkyycJZrf3A1
xOIBCXWcHp57QHacsPuazkivdtVoFtA8XcyW7Jaj/6G7DxTd3a2y+R2pX5RLm/ou
9XMLA9lCc91moIsIJOol+D0Fvquv9domiYmBFOF4usSFkoDaLPnaf5po4XMukjI9
cGjCudNDEWr5SCMSpHeqwHZ4yFC7ILhPL1bBH3G9sncYNRT0gX9TUxfupE5uVND2
36C6rfQg6b2oF5Zu/7gVGp7xUiPoQ+wryFS/mYkRHcfdy5PC7uURUqnM9O6Yc0fi
oq/1RHoGUST8eOckVYDGRU765zNxrrwCYQVmHa3zlwJLAi7WoqHKKPyAR/lKoo7V
r40iV8+N6lpx5V/sCyI0f7ZWguog6xsdrpJbNreZtWa3pwjRFvUsenBWW47gTu6K
gbnxp6OC2kWAL9yQ9Fme5i1i3c50IN4Vwlk84GlQSycdvFZWoH2R7qWGDRCtefWq
iMmHyf+wuWBrxLwznx+cvIQbCFG1Z/NvUySywykqzm+AR1QQnQ5KxpDK+pAxiTU2
4XIHrrWZ14NDi5KXeotm9gaIwgeV1wuTZAuTTM2ij66oBYk0GFSepipszYqrXngu
p6AwuetH1R/pfklC2tJOcgUy3/r/rXpOpJb31dEKgVQiXXJRGnX1oqgTHqMz/YzS
F7ALuh1FeaGlb/htLWa5VKStWoL2KmMo35yrz2dIFwc/RlSbL67Tpz6KpHUhJWvo
juCM8WcQ4+/GF9ntiKUBrQYmueVLxgpaGsBqVcpQ9quQxKoPV+m/v/kiP2280Tql
T7HrnI/gP3cS71s9b0k2ObIIhkwC4NsQTGxyFhaFJOlwIKoobOt45pWBFfUIR+nh
Npf3DQThaKD9kHt7Lzc1qJpSUouN70dWpACQKfXpxFlXmqUjkRRStqYvTv1lm8nv
mdosSW3TzKyn4hdY+/2MM8lkI7af7T9SwiZSOH9dAHGvKc+pc8/wsisCZMHolDnD
TcA5YVJiRSLJtpiR0Ae+uOtPWiHrRErPzh3RVELfzojqNSMSmz/8AtymsfJmBgYN
Wwk0xvkUd12fIP8Z6NP9vwQ34sVaBLNuiwlT5NB3Mvh3N03hj9vbucBwUOU+D4KD
B14OKTLOBGSISYZb1RPtP5gSdcQ5abgCBd8JwYHNSy8V6XybwgPZP6EBQI1E+CyQ
nrb2w35+1kNbXxYpSQx0g9qOetmPR+LUlxVSRCSH+D18uaNAuZ/FcyQkGOfzk/fz
TQi1UmCzeg1XKv65z0iX3OUxuKp9X2PpXjlzFOemhFrgSITO156yVtjM8tu3b7NZ
cAVIEV6+Kr5SAyjv2wjrx1zxLXaVJduVHyf05Z9Q/8D5Cfq8JNoFfrf57jmrScrQ
4+spngwz6q5Z0KnpP1Bp/SaLwgiIkdkR0V8M32aXOzpeovO7L14RhOwtXNTyiBED
sP6KHVY9XSmgWJy4LR2mld1iOFrSa8Xb8Jo6MjZor3Iwk1J1BbZPBTPr0MM2gKlM
DsZVig+dFbh79ZjQ96Ee5QHbuA0mimf91BlJ9QEVeOTcZObOtclZOoNMZ9iEgs+o
3pqTEvoup3F3Y0mcurYuV5Eo//GJgDHlwwFWol3z5tUrbxeAyrexeyWHxdH4OhmY
kWuLwYNng+GpcDqfwe6oqfvHvRDOjIJc6QqmRAbpQvTtsTRxmjwHyIun095xQGTX
PcDFCkGDriycVQ2SVTmyG6rl2zO8g+uCyL55DBXPJCyaDk1UM4zAKpCvAEfO8Uc8
MKys3M1KBqG/0W8lhi7PBMLMvKJGGtn2PGh/7jnXEqn40MZ9UekA+oHSNxPZQmRs
M4S3iaLDXmFRSau1JRrboReg9iIjy3huDH9pOiC+M09EkKs1NtWEofa0AawYwUki
sp0bvDlq2YTwmfjYcSlbwUFkKP6nfH/wX+BQMBH05nWmW/5tNLta3touh4eK5jJY
hTMfTohJNPNIkOS/j8pvkobKHgjCn64YYK+1jbPEek5f4vLeXyBtc3CmXlgGtvLH
HSBMBgLZtn/UYaQ6Y9SEozox3ckDJLLQT4D17jZvmVX4kUbFNgwX3hxM4ZzJ+hon
FbqK5Y+Z5nLya/dVNyYaBhT7D+oFlCUqA1lX2LXRujs+uxqzCjpialaCTqoT3WKh
TsrYWA6+L8ZuNZpziWQW1J2XoJ650yfbzr7m2sTRvdsyyUgXsjHXur9gggSx/5Xi
kN4i8A4on9ae5BwwLTlBKPyuhtq/8QO/vsvnkbDt6lT7T2Y5tRoGy2T3bVdRyTry
VKKkutk6DT6ndT7GmiKGJMI1ODROpLNAUAJK6MnHIh59WPYLkW/krkpvX2ZFB0VD
S/SLPbn+qXp/J5gS5osUkRvJYwzxk5yy8M/5Im22le+/dwPMv9qpFDyuxtERDDS3
dm3XMqMn2Y8VgIPMfTJ3UNkN/+lBLikDL/spTXTQVqv6sACBZhi8zuZqUIuy1Rlr
sDJkCh3KhDG+ADOyW1zh5tblFXYLQ1pplxsfy6gtGAVDJXtHZm/BVwVZoXU3wpzD
9yvDoxt9RjV1Oif9Tiz0vbujVDpufW1evubr6OGLGIWwbT1NQPBomnJeGPe5zAU7
Busg2yWjEqJMddy7FJ9/kzrtNi3saGISC/sCqIRdZjezDi2ExGfc6M9t7KBHZ9Bi
mI7S32TXMNeGBLSzomh5BHuPdC9q4K08tahxWCZUu3r+R3X+63l6FW/UJ0Yz8ol9
J6VCAJoxuKqemrQnQ+u2zcM0Z+l/mN6DQx5uCaItGnV/KmlKRJTti5rN+UrEfdWw
3SS3Y2jcrH9JB8cC4ygHl+dHJqvsPNudJ/kcgkYjU1zc+G5hceGQ3FS2L6pGKgT6
ezax+lskRHdeok4O1SpFWb9RIXGyIbKdyFYqBTMlORjd7XRkMLYAc5W47zSQW08q
6FLmTveBvF7z5BMICIdWUpwJ42ChaeZmlN68FRiJMTKIQAww/4Bue+/KU6Zg38bJ
5E5P+nuwmP0+wxKIPihkerCXS8zGH7CZ/SrgZ0peYMhgzEvieV/OpGtGNCRJSCzy
zxQv3YaIAh+p1EwUkq9StpAg3bo+ENqA3rtVBFYO7/1UVvuqRHbuRAH3p9Km00VC
DGQb+5qst1ZlEQ7Bg/rXM8BNu3YbPieQzOxMVa9p7rZk9SM5a/8mL9NwH/YS95+s
GdKMsjhd8dn9nYB1XllNFjGwwvcT1Rd8/oHgn1qHFO043Iwqd+JIfPZ1m4lj0uJP
QAnxeoz4s5UpY1YxKYwwl8E9LMTdHcac+sp82rXK1zEP1bi7plwy7Qek6twO4904
nTFvR6/wNljn5V8/eYwijV6VbcL5aJZGTZ7BulovT4A4BkOvBAr3kCDPR75ctwWE
7obWu/wIGuWfqfm7Ed4PfC/yzAfc4azk4N0kUc4kI/zzy48fj8Js1DNRE3m8q3OA
3I76QFM2FBcC6XH5chfAc+B6oH/AkRGqF5TmKnY5MgaXZYy7y6vC27QVl8/jBbVM
TEzw5Tnieq616zLpRH0cWMMq3azsWnU6fnKGXPEJxbAxu5v/NJXnTmSD4Q3RkLzP
yQN7YbjagN+4RSkXRGAej2cMIDrUk6yALA6ZfzhiIc+Irr5NZ8nyVMObPrBvnokD
xHC4U5mpwX++e+x6sNw/gaofMj4iuKeulICK7TzXt2OaUCiiBLqPWj6awKNstFjv
Olwfn7Qzg+mq278M+Te6GvPiiHeY/fulHOfjxbA4I0ZnG/Gz0PmbVQQk9ronRQn/
+C2j1hCKkYMn9VIHE5Z44IZkcERJlVdaoESF18WHu4WgqGNfRtNs7uZWf5JQIo/I
xd4zPOqp0x9a7y8n5plGBOkfrssTlUuhcSYgedtcwFdQLZer567zksRvnT8RoGkj
HwAeNFDSqSX1tCSOgRF9NAtVvfN+gx4711ADjDDPK0rtwRmX9a22YnHqFYUI3EIk
MDqonGKC2CIW9C+iL468EtHUFTEMC6/rNO4gwlaFyyKCO3E64/WsGVIL5Qy9yy1s
fdO56eiJecHCSioVzJASpLZ3XdfZSRzgStFBJ3mCS+UuwL4QeHwWRyzz6tmd8Yao
l7t1m5DsTnjdCgH6Z8ZospqBhI/L5TzL/DSQW3jd4oxuaO+xBbIychtwBVtn2rpy
yaMD8XuhP/W5/LHajYf0uyjLCSNq1bfEPtRFn3zKFXn7Ton0UDe/Cgrcwa9B4Ptu
rU4Gse9mcShtKCE/F+4kkGaBEQLhtpqLbkMYYYmqm/5AtaSn3lj9gC5aQ7CTrLyp
iweHC8Kcqh2EQP8fgRw5DI81JKeM4vQGJ2MSzowT9qQ13XkDb2kJVYOay2GRxgVj
Zlz76uXjQZWEPIIRswrA4GtbhhtHkVFTelH3xyL5gGGzkADYyINR+7BVPXVxRWjo
pgx5Vl5uxv16g0AiUn7gLhNhrB+cVzKIhB3oDj29zZArb8d+jYD5qgmKfDjVXbQ6
5NMyaDpWzEkSGrlsd5wXQF1GFGdfkiYEomWrhVY16ksktlXWBEikLtBFprXgU2y6
Ev8pgio/ZW210L1HC0s+KYTw3xNAWI2B1L9hC8F+n93k9gA1BFJfqh4pWJyW2iVF
PNunq9X+ww8vXLVcR7vSuRj88z5iIedRLK5oYx3Nk5o0TlZtD82fnzoZFOhtQ66V
3PxE0RrvvD0m3QsObJ0ym8SRpjxfURfav+ynUS9jhB47QY+tV3GsVJVsajLEahQM
zZIHolJNOnlSUA/9EAi2mM32E5INHvRvKUBFqfnsxGrShNQ8v5uDp8fu5jRiJycU
zOo2L3vBEb2swq0POG9w+XxAGEg0rE+Ty/65d99hDYvuVh7GczUPZfR4i5YIhwSz
uv+2VuuqII/a1nQmXZ4M1bsjfgx5OBUw+tB/8nSSGc0U3vOXIjoHUfZak0VIvUFv
Ephg5s1BT+gVbrLhNKZVfsiclzRZZQpjVoW2mNcPuQgVI8uXpAlygfQ19sSZAsn7
5S0mwxb9rip1wqs0bCZjsInA7XC90g+qMbx3oeMKPsox6ajjHTELwNttugCcifcK
Wyp5RvFXaw1nqtwvGByqE7Pe0e5ONxLW3C+CIAQZWBhgYXdWpdn+5EoHavCf2Ksw
SG2iL0ydh7NM07sX1soWx29nZk0tnqLaHE3knKJPXE/JyYCoFz27v+cJf/8FnPt0
h1X5Wl4+qNWYzOOzOmXyZPzBEsK43Zuq5bb4LkqoUglaNzrUYTBNkaoIenFSxFWC
7IlC5tuibwOFe8zymFBD6Z2pGM0L4Doh88sw/AIwDcTQUdvZnDFhvNqY/NSV9oIz
kPoD6jFBkj1O3g3XVEUj50HqCQkCKUdbYd6T/o1/FxRjP8pXMoIg4Lv4UgaHsLw9
YJCVULZgxr68SZLPZkPtFg7ILBKiFyGE8uS8Qi27s6HW5kuEqTI2hddLj4QRVUuK
67wHzJUNcA3CQ+IxcBnFuySAMYYkMSdPuCXALtYsqIjkuRjy9cp2fIT41yHxLC6X
yqZmUHWbyyuZvN2Jwdn9JoTclQ3kGIFq9P/I21Y2SFV4Np6rHI4VthU4UWyMmykL
fHuNTSfpEmDyGEbZq6XHGopVOoZW7glc46cxCQEqchlg1C9ak3Of84DxWlBYSgS1
udAy9/xMWjimzJO07Y27H2BYuVrxuD9d3hqmEyQwfF8bV31pzM+vz6TCYkn9WI0R
057ygDYMzPFp4HRH5MZYvl6qEIuCyVPj7sEML6yVSAvQUyduD6ulQnjZ37NDnCBW
zCvfxEqfpBzy0ag/HRElTz08NKfcBhclYx7xWVgzOnfl4jv5LLCjwv+DWeB2MCg0
6PRQdaKXr824mtp0boKFbaWrqNwDCnYeacFA2eN1YFsJzK5+loxhKkwlPOTaYs89
eI7VUIu0UQNuTyk9QyUHEXwfskIN16ttsxup0fq8eS8JmFiXkcS545XL+p9S6sIB
YpR4IaudpaLLE9Xslu7QA/5/8eMnKolvk/wkyZxYXiXqa6mxTmkoPt7NFG3y5vgo
rFRkN45/w7wjeymSmmuhFvNQ6jzB3VLhUUKnn0DBeNVhtlSy89hPdjlmxqJaRvm/
JcA4p4UnL3LjxRp+hIxZVTrC8XDUuU3/BFZHei7bpo7lH+5rpyZSHUT1vjSG0W/G
RHmGN8djxxpQ5h+HtORvC2bJv23QZAytbd1tIttagCFq1sBqWO96zszE4IwuYo12
wuGmkm5VYnHFpkzF2+ovZwHzwTq8BRx101dLnSFj5wiFVzBOyrso3ckqx2dCU7Dm
/FvBzOuRVbhHBNTCcPIr36umwJfb7JbXEOnpNg4gUa/bQridNSgP/Njxw8RCQDh4
38i3C/2kiY99hZ7N8L3uKVOBt0zwA+Ugi553Ak0C88qLULb68f9eN2tKmoTGmUIq
XYUKJxVPnJMY3gU8up0bBqiyMnJVA9wJYeivIbu3E9IuI5rn+UOtUSNEn76+pFK5
5fOWKIrAWK86aR5FeMDDRRSEmLapYBJXd+odmSG9cbcDIkrNra0xU0nUvt+0FR7v
Q+ewdhTCukyCeL3tAGMRVrAASOgvBbw961ZeB4m4xMp89DlIc5BCD+FlnPEM8XF0
Gs8vwMU7yA+JBPFcDYC/ZOzFtAEt3F34rPaPqoAYu8/qq4xZiuNoTVYTa9zP+BFG
Yq8gJZvKK/4FFsAj1JYwRpMVXzKYu0wtJQariugHKT0YiiPi2RxExJINRij9ypJl
tBKGlgI+nmK8eaqGMx0Ghk/jVeu6I7FawlkrCMzIK5nBJHRRMgYGj1in2Fng/vs4
eYXiVcXXyququlYGi5qkq6piB8U28m26OvAA37NrQ4dHv11F9G9hyHekkytVS/oS
Y667Tr7GmtgyV54QyYypKYx8GlDQLMoGY542r3XCDVhzv3IXh2E+bZdlovVgR0On
WaqZ8gVNZ5p9MM9AHFs8T8qEWAyvYw5kPF4ZrIv2BAXepNej/nc9Otd+WeoKeyI6
YSkWtfb9OC3g+QgXHzP1PIEX6cKRhkQkqjOkr+ElyfnzyKkgpZ4ylwUZQ5Zf+WJc
JTAWqeJ739p6KpGDwMKIQ1Xy9/qNJTAowiPKKclDKVD9a0YInSsxOxgfFEJ4uM1t
FpvOlbrajOJz/VZLaR+YlwLzZXlaRc67cH1AEajQu3l+Bo/gmF0Gf520BmH7vGh1
5WrAbqU4pEJAbMiN+eqif09MHIbwfzix3xEkSX/6/9/gZPGimGnVlr7mjjgoSQ3W
fT4I7p6QKlvpVK+B78ZLZFqJzQ7s9bOjVY7e1kXVRyrZyRiZyrUP54EWHaneIlWt
dfQjJH0Y+EHT2smgSITqTOqtepD0ju+Ptra1ej8gD4geSNLgpjOlGTyFYBH+PKgj
zuG7Q5Cw9GbUgbp6jhV9z5Buj1uw9xRNt6y2Sn9wlc98gQN2tYQLVWjNX74BIbST
Jk/VSy8zcSHY4J0VPeLQPmKoEWjEgi7PT4F9k7bR58XhmT/02ltmlzuuXjH50A7T
qnoJIkCioNI+W/+gZlRH6gfmljvt43O1xoBZXuW/NlAkkwsRDOWsSgaCv/dJNiqC
Gc3PemSC81JGX4tnQQQI+hf2cb2EbPnH34ZVVgiN/RH3ioJHtPwOsTOglG6W5TqJ
rbRTdsOwezA8Wfcdi7AERXqp+IA6rd3qHsgas4R6+VcZql9hPy7JSj192yfcETyZ
AAop3yhRaUmzroeIilRFaFAm+gDB6a76EYsn3H85CXFjVxaSjROAOEXPa9IOaFKh
RYwjR5NqibqJBUrCX4yyxCLX+2yXqoBCpms1ovfe4Lh4xdNGTEl02iJdnqOGJLEz
IPN7JfT+sZEuxAfcFHdDjsFLgEcKM99LQkvdG0ISxsMhciGa9mc46E/iVv6hp8je
VUl2VrxS8ydVJzIWSTE2iHPXR/utGi0ir5Ua4vX4UIO8ZlalQUfAtLdroGbVNSvA
8QAN3SfrWWlgVQY0PAvtvwDsN3t0f1aTUY0/bcQoRROVh+IRUmDaR2HNCd7b6ED5
nkq+IbPNK7HbAJNKaZSM8Ew0YISy+ZJfFog1zTVMPCDCnERKZVIVfnpqU1d2+hVb
fT2UO97wZKOWDGaLAfTOBxFLpobjxMsfwvmYEd0CiYN7ZM7gGEm1YOFlrq9a9cMX
aiMuILg6aPzKFcXPhcHoYU/4oOn/FQAmePvs432TlfoNZFjhcNtDxkgGpmvaNLUk
GTGOZRUhrbI+xHO5pUwb1HwFpkatLQR18OSDqcieUBF6TQnc42Y78w+ASKAA6yIT
UraErCHNtBlqKigocjMQAnMox/wTf24pppJolcNic3B6M9DPoJd9ahYSOJqD185E
VY/6OPPdSIY4IB1HJcJT5vvzKT27oKdPxO6+VnIlxf1TIfDxPZ0sNWlZr+Gu6p2L
B3FQOueLbDGbR/p+PGPf0LJqL3GdDlTRopDFrZaHTMdTTphOjpZe3TN/y8EmxdA8
osxB1WPZ9m4H85XmfVADPx6xc3rB80e6kBnKSU6/1PC965wP7BLoQYg0/EQs9tmI
0IBxR29YUCD7YjRnRcau8LLt4a8XMbikWwpe0eMCjWh6U0tSm7aV8XM7psBeTAzv
aqcZHHUpBUC+UEs+2RjXmqVYTPexpgYbokj3RD8q5AP7nmpHOnlnNvCjOL9IXlS+
S3P7IPoLL8EhGpXkI67na+7NeKOANhhRZRtl1Z1ujo65sinX5Sw3gX5r7nAdL6sA
KupSs4Wb8hSs+174jC8GxJwrLK2VktrrfgSgr6Zx/xPHYyWywV1ntoQIF36QjP08
g5TknJ4A1xveBBzcadDjo2QeBK7qWt5pgXtmGARPEx+bYniQGsG9Y1LNOaV6aVK4
fZvxM6xvKr7BFzEpXLnVgRfqj/s+D9Sc4ZNXLUCDggyCAbaDoGpkzJZ0Fm/Gp7vg
riHftnY6lopKOzIO+cX4CER7sbhO4zUjzwOmgKS7UgaetXVs567slRXWQoCat0mS
wwz8dt+LUS1o6aEFXTGEg0pWldsZM7TLR+9g+v3xbTYUlTrTkc0Rt5lw0s6yxTxP
N/M4LuN64aBxnPJfk7dXin/Ki7ww25ssTzpK+NXpQnPJduBMFXBNXHH1RwrzWvIk
+jcLPXes3kyDv3NmKiW+xMNIPkQIm1biEnGMITDTCBH7UVaWipe3TIuwJjy3iXLt
4kdELIdk2UKmnndAgphsto9GmkzSsXeQQn520co6pWGmOx8XgGOZNrA3DqHV3Tk6
cbVxSQSuS6jg5aRdnBDi9Dl5Myt0Ps1X5GLHFmUvJkUrgAKAqc5PBncux/xJ2K0y
EWyTVOPLXQBo0VutUYfdE/f3q8ERickBYW8rwIcgwu2PbdP48Uh5xP2d2z+BZkte
u40FFH7ftLsbJuFnvzLaXosvhpmT4BF6EsU9Fri2amp/f0sFBeevwcMKgmPpYZqb
bjj4GVxh911pucFeXa6yC/eosvKutGTg3wKYIhDGVqhqcD/fvKtQIKXsblsiUfqw
liu39zxcsEZ6qxosqGbPsMfu5Ef4KM5dQiy6Eefrf6u1SdgbM2INgKHgfxQA0zgm
e5N19Mo+u/NIwpOo4k4cI2IoKqWV28Cnoauh19FsvMcyGCWrNZKYbcwElkZf+/hu
bsfJ44ZOhV7HIKFu0/N4A6lOwPOdd6UzW0Pp1ezmXiiIgsDbOeaV6lXlm4Z5bk9A
3lloceL/6a6ogX8rLemK/25fdEiSrt9t0nTqXr0CqZ5pwsFtHlhn5NDbLdffk8b0
GXHekKu2e3UY15HQdc60Gf9b2IA1tuZX0aVL7n0s+K0uZifQpqzLh19uLPhtcJca
hk0VsCUYDrUJSNctrKPEYvd3ogX/gAsbYB79v127LE3aG3MYsXucqsBcJledCpqT
x4koe0pejYA0AiyZtXncMpEoLLKefVfEPh2kwQ2w6YBnrlryck3ZYS3eqKxmjei9
kt7shxBaw9iIyvrxrefOMLBJt8AhVbz+ec/Aq4H/su0C6+LyJgdiFqNc6ye7gZ83
wuuOYfXm6f5367m2paEIGlMAmV8ivELClLljk+5yIg0mvpaFCKIGptgBav4bdPcm
d9lJ4g4IPYt3vJUnF8fQsj1EiKxOujM4N6phukMds69QCwtrxwC5u41BXxb4Esb7
9R350wsV7mZQmonRi32btWOzSQJIFdSShk368nI2jIOeStjEiPuqX8ux3s4SkpmA
SoJpdtSNYU193qIl0N3HYMXpZ/6nUsqxTGf+ctzshyDV/neIdv2bo7zAkMPmk5MA
l8+R5fa9rU4epftDSybS0U+AYY9ZZD2KXPSBn18/WUrEe6arFeUXeZzzUj8Se8Be
JIToZ3orAUHcaCFD7c1wqEgkxV7LvuxlREdzWQ7ncXhqVvg2+sf6a2OhNzs3g1pq
1XJ6yPdjk0p3sf3Cq62Y2993qUXnumtxqhBXVifIPmSQjbqN78RYnqoGJb0US/3x
cGrL/JwOCIHzjDszwsuDZAxCXHjui3Wiq/heIZeKh72KniqpmVUTNUJugh4La8Ga
PMdGVSWe987mxbYRIPRNM9C/dx6A4TzCDOq4LH2GAJpbyr0I1W5Ax8nrEboCySFP
73GXcH+02YlmMk6DosWnsRre0DumtLx+jRDGY7b3FEI1ZXawab12Lau/QRDkDRzH
At+0Dep3Qa/g8nL4R8Ep/2jzTKOABZCVQZJjcd1zxeZ6Se+m9TBCghOrkSwfujNk
WiIdYUfIGeyifIYcWM3Aity3YmDTC90Ustzny+pazk2/2L+P42keMHTOZ0xzwEAN
AZhNRq5YErv/kk0FoRwIOIO7ghYfWVsYzvtn4+Z77TYJ6L9zm146AUivFV50t01/
DpYbW9ShXOANj2TZUp8llPwOKwJnhlNasGRyjYxhM1n/SFt6qLt6bVNhFMI/496t
FywmKOgO3Gut79meoLgPvuofUvRej1T2xMMW5xs7pJo+d+C72PJEGzunvTMQp+cr
idk26k9+MdzNhXh1n0p2jgvzCJL+Bp9PnTbarc3gJtSsO1tDNjalO0Uv0oirB8fD
C9VZNVLEO8VjmiNBEXWploObQaYli8o8Icc/KOiy4BcuDq4bLIt19wcSu9IIdrRJ
l037gW4ys05kn0bk9O3yQ/i0mPavMWi2Icp9Soq8rKRGwlGvkQUb4/RANXWMnirY
DEHbyq0J7g8z/EDKHPz5RbuBk8WoBZIol1M3RDunlQersskonSpeKapcTyMGk+ER
wCqFUCNXo5uAl9PR05aAMbvkqdqQ/3mZ6xEfMBJM14vLW+ncyahLjOmQyLXgQkOB
Fp4qsIfVnDDXg4W3dewSWhk/47ZhMHZSrdfP3ht2Ajrsh37MUhNPBPS454pGfxwb
N2e+1+67rpBcIMu7nGNGDdkCBZ6V6wdJS1YBiXI58DOtrBqUqLpxFraO+86TX3ja
pYSALMwy+dKk5QK/COrU6S8VKWd5UZ8hmrS+bGk1CwZCQswW6e4buFGtauA3nYmA
C/zzZRJEnS64pVGu5rNYEawrX1S6pvRkL6Z0hMS7SlAkRa11NbE78pNsd54oWljP
18kHJZU1uvDgjOaVNCjEmX0g0xQDT8a5eb4P5tj3abXfkDPPKMXj2eFAVSHAX502
0RLtYTBtClM/WJIHQEgRN0vhD2A5v2y3kiCR34e4u998t4Zep839BlS3cLaWr5eE
l+0jrnnOAltXWx4fD+3yGqBeFtMx3eiWfozva8oqaIGpiqepJeYWniunViVx83g1
ISBYybYJwmY2Bf5kVvT8x7WFuMyThqTTcAi0hzDF7larl1HrPkrgNpAEMgVc62Kq
6Oe9ls8aiNnJf9qtIs6mY7uHvKALiDr8qmNOJIpUQq5c4kf2bwnA3Ta4+/ekSz0C
NjaT/r5Pyj452yRXp4A+i+Qjg+wfvrrLTpghem/FzZf+x/7hGb9t1zTGLYhkl9Qq
nB0Q3s/if1ieISXrbQqZyYP6qNGTFGnhbn0ftHoNeGev1oPkdfjDcKQoreakj0+A
JlnbPQe6vNxDLHYeqyJLxPmUrCkjZmogek5DH33azec+3NXJkJGEDUKVmqZLFCjZ
NdKa5m9sqCjA7Xl5xhvo+pdfSu0IiuAAyhT+d66tP2CTX+UqjPrvCnqMdDWjBGIS
OtlNJ3fGxZpUBjqaLI5cO1bO+jwwjkkRPwQa0QyfTS9Wi72EtsU1wAx7cTVYx5ya
TmT0MU9Wqh0vX+UIjR/lDr1fwSUoP8SJa0a2PFAJX9FMFdyTY+5yZEibrT0dkrXc
2KVCwNl7e1iioNP2guDx76lJXLV27yFq817oZF/9A7yYMlNAJdHKvddbwewGSJ7b
4Cyqe9Tw1hRRQxdullAM3NM6W1HzmPoL4MzhT+0/uIlxpXqsHrDdCq4yo/WSEkLL
7Xz5BTSDBIMjpSbO4agsyS+zYJlTyUYGBlsAn49B+pWjUCzo1/+kzDS7n7+hiGlC
OcSIOKas4VL5zZwj7P/1gkQZgn9yAwlOyfqK0No3GONyardjKoMj09BEDe2FQv3f
CJbtvPufa2IMXavOl/ZGp/2YDQJ6zCn4uzvQNKLlhbYi1Reo9s0QrIyp7tCpvZb2
kC6TWxfVgZEqe52P4xW+RCk1CgBigmCJ2UQ3c5NvPDqyalF/l6Zg0YwmH5uCoQTw
ef9wNA5Hq0guTWN/Vm2T6uUL8p694r1CnKtlxCnTI3t4xUhUiXPUDwMQvkTtc6Dn
Sc6fBnIFg/5iw9zWS9w8zd0UK5X/A9Zut9qdve88rfSFeuUH/9MQRAD7cJONMU/i
404EsAv4sK3iETdIge5htv0ZPw+MNR2yuQs3g3w8gg29t5DOSbvO3t5Aa1rXKYb+
LrwoNnH9dsbKR3HXOK8gcZq3o8Z40ra/aSEkySalWIP31gtiZHxtAJ34H/5ApJGU
is/Yk6P10w1Xk15LYBD2GO+2j4QlYo7I84ROZHVuOy0zrXJPqxrdX3rh0ID2CUn/
Z+xkv4FsSRh8mAIapntsD2c8Vhr0GSBChy32vQynJ2PeRmxn+XCQQZ/zWRvQf+Ce
CDT3yMxmne5U4OAqo9LT9RDvufNe0AMVX5eYIz2il83WqbXGFLls7qY2qZV7fag6
3INRX/Up5wyFoOw4wrsrO+EbhV4qOlyXkgZOspkO4sWxPL1/fZMCE8Yq17NODbqf
BK+2nhVBzy2zfvSSU9G5dGVNM0JYmCIdYAn6SACYjBklviHKj98lfxjjqm17wqvY
K8U3OaTTtLUoYCEZ7Q7TNUTrQ3ZOkdIvnuBestpmqiQaRivwxncWiMFYkrcplwGL
pXU3EkPiqRd86qW//RtKRdQXpkrhjFjcyGZtYd+vFOsCZwRV7MWvIpP6/stuvA0K
EfszbnM/zJhyHqV/xqyCd7XyNvxrZEB8XC8P9lvWoBcVrlEApqYqN94tEa9kXMev
nTV3TJWe0XUBdGcZF8luNALfCOClFJ5ayGoZYFg2zy5bcaWvdzwlwaoSOqodFCni
LcmavhuFAKCUxFoXB1+qh1jFV4CwWO9UMxDxONsF5ZIWIaoxTOE074TTuOKYVIfk
btigynwQSVNZ/Lgr3H3faW+N5cZtQfIfbFL5RpfYo9j3fdAIR9Si9XY2YRAJyDY7
riIhUU9BM+trYkghgF7/P2MN7wx5zCAIqKMA9ACIfyD8nmhGsXfCOUZDE5qeg5Wb
gjoADFaXGHx0SeHBWcdhIomIB1u1PF+2w4dwbA3+NyKSozmMLOuMqEEYs+OoqMo4
1EENntzWf6wd1lRzgPtxJoXzITgG+lc9xZ5pQ50ItOTqeCyYtKfBdV5FE6xY0Xmb
aepcwshFW9UHss33z7CGpEdnrKukQBsxV2GcmBAANrTyqTCPgSeAYPsdAFYtuW0v
KBreBLdZmw+ssk49t3Pzbm+onOW2agajnVByJ1v79UU9q9SSKU5mFZTQ+EBEEFAb
QmeKtWPnKAnvSoDgOH5uyxemiE7eszbneSTMY6qH33yZwxVxNCKDe+CUDuqn4qHs
pObt6RlAGKAsasKnfs2edO8HnO4G0uK1AJx0Nor/IlomhdSoYoj1ayjBhiIgn/tG
oQKATqRVWxk3icL6YDAHpBPKhpADcj21d03MOG/kmAE3aBwUCz3eCzmE9fVi9ExB
BfDwAROqcDbv/kcZWen2Oux8qLX3Lm3549nh3I0LI33T1zc0XZ7ESFBp5Fh357s0
gyxHKcOlNHBc8uq4QLOS23z2t/IOpZ5olNZ6kVD1UMDxJPvggt06kXM0T/bnamqT
D6OycvKvocwlCyl6CKnn1fe5QiIE0ukhbAhqzAkL7jJza5l6u5RDYCPPFbrPU6sL
/Hv1nhXz59UsCwR69jHQelggvMxntrYuuJOWQzl6vp/tA6l4WBT6y7JNQukZa+V6
H6SB7kUeqqARWtxON0iUYl2HgNFwPU0biJI+DQamDs9zUjjf9cYjsKTNmwX2C1Iw
35Kg7a442SCDM7hUJONB+E7+yMudsZmnF+8U8tQFCxenye0IE3TYDLJQWykYqFFl
lPy/ih9aAHm0rej6dhxKC95ZWci4p8mVVSdF+entu3BDhZM65LwJTlIKWCugPR4D
dQxut0uAWhLs2NVJ9ATJZbIJsZSU7/ErPQ1LgeXGz1pcFdg+sYEXYdV/LKcLCvGu
Ympr3Ir/pvXcddr1Gwho/98knfTBLLW5rgxeylyEfpEauBLn1k7bYza/eoOXK8nC
9WlcNJ96ca5rC57V5gyy7bRun17Zbta2vqYhxgbCoj3EG4c1NVBphz9D7uPZCO+d
cdGzIoLg1q6tYLLaCLpffHGc1IC9HoVwntP+LFt9OaoyC+22HPltT6FjuA+tEZ09
OMN1vcf2Kw/e1RRDikUI04VsSnXcszxkWfh3arA38SmACtpHzhqBG5zfQGzenmR1
Ln3wQeYBj7lrRhvJeiP6olRgeEBLGe/FR5LHkovvWkDCzyRroWfswwo6leBb2HjH
xCe6wZl5sXXvMdiSiO5EAT/YbeJwWtWgH0oYpU0eyby2NDd8QY3W4QlisWXAMwMX
b3Ev/YciCV6URPSLJ2Op60/gV10ufIv3wUZumww2NqCF+VV97uo1izK5SC+qLqMd
1iYMYTOdfDj4uJ5Eva2I+76i2Q8+5ONSiB57dKZH7C58xsc/HwTh2RxBO6XcUc9N
mIWHTMv8cEDIq9e0wpp6bNDE2evhUt3K7V00Jvvm0uiUJmEFEeIZYz0IcX0P9Pwg
Y7uv6MrfYxG8LOU2/f50YBLa9o0w7F8HSLu4CeABK4aB+iAjPlU3u7HCKMBoMUq9
fSSrfwKrYHf9y6pT+ZVBjpVVVD+p1dXlYPO3VJ4TJyF2hqtK5vnkQDY0mPm/2Erj
BK84cm8975fgdcy4xKWPEuq9w1Lv1o9uDJg1taAi5dgmlfu85F54DLA1GZshngjc
qCIacPxLxTU3cLxZQzmTDWpJdue4ndHXIlWqcZ9CfWS1gSv7Zty4lQZIEuH02iz2
ydwhTg+FCmZr5fKgu0KhxVM/gov7o9/vmSaFMpo7me/C3XT5fFe0tgZ9QvEqZqN9
xcLEEiGDtj9/94FgYs2FvPo0+ASFPNa1AD4Wd23nJL9cbxOUlZzSJVq7HWqQLkMA
RigBJjTfj+x8JDI/KyaS5gDTH6quVOj4GmEAas2eqDqSUAbhtJk+N4ZQheAoBYx6
OvCOGSj7gBjnOjUIRsMRqjwRmTiWRTv9xgkGastg0GJjL4B0IHu+EQMRk/IOiBiO
uvE0OdYf8IDlRRwKuZZpQHbggR1sapOA15JqKetfbyhK533d0UCJgj0ETr3bHHzD
/cB6sFrYUdTfOuTmAx7HhuLyXBnEoicM/iVrhRk8Q97519psFmpRRRl+K6M54TMW
k71mAkkkWuW/ADCzg0MxMT5dtC1ic28cGzx2l1TtLyT12EUkWIVhjE0jhF9hhkZu
oOqS5KuyZImwi65d5Fhrb6VYzQx5U7GXV2czBWptRiDAIDjRL3OpZ+c0CZdg3muQ
fWzcmN9nSdSQ0vXUvV9p4odxZzBQ4wB3CuZlZ3fgcXw5UmyFq/U0s6iNeQzvZd9a
jAXALPKwjJnRwCP2SLRyVVGuvApX4rTfNlpdJVSiJtQE59rt6Mzco9yZKvbt6IJx
WgdgWWYgjSKg7OuBMl8y2EgS974EZ32RmnUZhKBnaIudgKO4gziVR84y3kXLifsG
rq46M85hUJ2kSOUe9gfHBwSfhFL8cBYVgyKH1+tYwut8ugu+foYqAHQxzdLJhlq4
+wrnExc4ZfPxly/CaaqFNBw0xW05bNMaQ7ORfiDfKxyVd//kjVjDmetRa3BNr7Lq
APQhQtZJZ0tiL4geZEB4CrBggDJqdUTcwO1Oclf4AxfXoGR5bMuXXyfJMWrV82zA
1hngWS53LLlgxekmtQfkEoqcVyiMUKSmTGMsccsxQozNw1K7d2EbYGiiGAHNICbU
0EUnRVFuzymMV3qZfi23+331Vk0iBfoqu0ZkK0AMhdDPNt5LHMMA+ssrqiaHcqx/
/R0XBxLJZtehYR9xchh8LRNPBF704xs0GG8mA+yVSyZGaAAkEIHWfM/QvCYUNcUL
2b0t8nUods94apmE6iKV7TgOdcVJqx4uxUjSU8v0eE9ddaH9+nbl/OsCMUBzSAOZ
YZh6hXxoJzvrZ9oQjN3h7t9loEriVgyBeY9qSGPHegMgvBa7dZsWsoc41YRov9ig
08EmChMd1VONP0Rh/Jw2T1jnL07TGgynnTH+e4I18KX8uLDkEiPXo3/f3iH0csKC
y1jbAnpJDOkCDRm5DsEGrPsy1S2674+2Z+BIsyg8R2fsRdPDN6REljNkOmzwQ+8y
1MevKDA4haOyT1Mxcx3EujeLgmd7fATDmyKN5W2dS9k5aLwbpxGqM41DjLDKuNVy
jQL5lgLwZqja99QU1id7V5I7vdtXd4xLIIeHfPtUo6D7//W20KU0lli8B7EXK/8F
JxCT5ICT3MZuOO0kvcH1W0oj5G9u1ozu0qfKwoGc3YzdqOlxgBKL6pCFrrkGfH1o
iyITs5HAnuVfO3ebkmlJLo8UM/qY8nmTe3fTYAJGdI6s9+RYD/EmfmV/+G8sUlpI
zIVCfkzQfKLNj0EfscRsp9DZKAdr/Dd6dpa9jGKQ+YTJU3k9ZhjJJKZs27tbsem5
/klyDeerg35++uZdBko6XL78nSUr0RkDtxtY83Lslw7And2OId5rlIEabhsN58hP
vXGMP2f985E9zNgrJxbHsWcO80Yx/4rkiUUDQt8atkuh8VW0jJDKKCH6mb1BaKg4
CAt3RY13Lq7+moUwSETlYKiUazcwEAsz5jPJKEpDx0KX6lpNr+16sNJ23Rn6SrZ9
+RNJbzWPYsLRSAzOFqwjlqIRXv4dWg+RbVUkAVlFEG4V0JAYdu4WrPaHxTuQTs1e
PVeAZ9w+7xxTp4Dx+5fn6n5jHQDnk6/RJBxVo4hzA0G8XYdsIn9+/D4gaFK0bAjt
oi8noGyFl6O+AvEn/fr+5Gm5BbRNhAglzvaudeGg9ueZzt2cMA62sEKgKGzfiHqb
7qjUlMxhHQ+Yct1owo0Ysq6PC9tYJazrS++57ka4nTNh6RSKYaHeCU+CvxOBNr6X
cdtzgWwrrPWcjRPQBJvMVcp2QeNRdLsLA51Iy/W7wfBkU1ttp9WNa5aI3khG3980
chSZxF71vp7BSsrvINKtaosGcsh0u+HtuZuDW3DIQOQ/4TArA4XiD3nOAu4TOGr9
dJJflhY8Jiab1yj8OySchAIALxHyr1RLtj9fwlpLjanGpa1KQKuStp+B9e0HlvW8
4SE4TdGtWERauLZQZNR9SFLfMy2+HgCr4BREz76Q6G3d4BmNlhp6XD2+vsJbYQOh
6faVUNdAAbN86QnSRGIbi+CfpRVobBkZ5apQEYGGiXqkfRcSjEeLaktAz0h0h7ya
1d7o+KAEMq1uvE+6hhAErxEgfeP0lhWtFfxzNB/TMYLXTcQMFJdNfCNBdTau0ll5
PBgVKmULtbyopawpJlasn7Uhho15FC/yal9IA3715LRwwCP86PNdv3Og/lweu13w
njdD/8W+Yhu9IJhbh7B4xTpDjXSp7GP5hJJmd5Fn6Kaq9wifQpVrIbvNp/626rgE
KNciphJTWi60x2WSv6642iqQmr5N1XeAI/16e4I9ceUjomL9FVvipVWWTMDCdC+l
2PoU/woc7f0G1QtUdvAqyDRQslzU6AAfJKyqabDx6ZHD+jQvdlbBMvX3aCjyiB3m
1rsmW6XyQTtifcjKDuguLKffVKY/FlpHLW59oHthzhUgGOWnklplSAaeaw0+7ogd
QOghTd6g14WkLm2XaKB/broCLRgrzz2/mANmPlLu6Po2dKnic4QWMJoD2lpBjN1J
24E+Ynbl+f/NoSHi16SoMV2ycLXtn0/+i9swOGA4IpKjMJOTmVBarvAS/Y9wMcxj
zSaVmHgEFNTUfSaU9Lbd8FYrbA/sRm+gMEgWZEXxr6y5DKkbIt9rjVQECimEwOyN
wF+ZqXOcjnZ2U/pSRGjpGrgFvK8idlzavN+Af7ZroQrwT6fX65SbDqD4ZANtzCC7
IGf4BfyhrArHvMqfTIeN5Nl1HQ2ZBXTWxVgkJhEmFEAxuaDf78Mzw4SHgs9MJoGa
cgjTBl65GUHlaBZTodQCQQZI55/tPEyzP9qDWMFmGL4n9j6IJNwwkZv5Chap9uPU
ewSD/uhBdJu0sd6ReTDCeOmVHJVEuUzbXHhc4hl/iqe8sVl+bt1eEGb7p7qDI80P
xNvKaRBB/IKgYgwhusISXwjXhisZzKSxq/ScWxqTzcXW3fwy9fJBDmcSTod82GUg
o1cI3g9IUY19M0EvcIhPlEHy0IE/FMyjCbLSyeKr7cdedSKK3RmG8NIEb49REdVs
SU0q+1K66KdjgcGXDMuY5OfptMMdBfD5GUnX3ewLvm1yyTGM3KaWtE80qQQ3qAnO
t2NYHmfVzXsvqnQthP8bT5bgOWl8TjfVupmg4zGRFfZSb46Yw/8Z+Vtk9gKHhNLx
PM6Nk3noCi6hzALkBBXMsXgamAIVUjbK+xEA1unWKFKYwdvl9DkTYFR7XwrtDHqK
WAWL8gmi5sS8O5ghUPJrl4bP2ehUTN8RacPrz7YLhjziFnebv++FURELrfaT7to3
8Sboj1S99L0mcbOFFqNjCl7QKZI6gVd3qrUIf8IIfCG2cXNb2oc/TfH5xgSPLFOZ
UddsjTPtsoD8z1Tm6/EaosHMJlJceq3KGZLpYb+d0Mwdn6dzhlJ124hA9O7TkGVw
DDdPUcaxuAgNhyzS9CBRr3hMJpE/HizRSPyXISzXOs2UTgJMg/uYGFwww92ypUDK
/xpkGukojLytajw93sQ/aJTFeyfkW4t1FbwT5C3hNHEavEQaTZj9FsN+OhccJTLq
E5oOZb1yXROd5devGy2ZZ+rfUREDmqsAIuaByJHU/phJknhCOamNiK/33vSCj1Qm
rHdTxaSYg0Nay7Atea/GFPnfM6TF6yE/9QnXUfrSgYr4175p5IoXW5h6gPRLyfj7
oWecJ4mIzPPu+OVpsS+gb8IB3+QpRGNZ/10mIVkyMgM4O5O7ymNJFE4ciJluUlQ6
KlUAvmLYs05OXbgNap5T8yuNCbfmBx7jLYT2Jmwjlf5QiF9mf2C4VnHmjhTgxSM1
GNNNa6wOXJ26L+htJliGFxChvosZGMRnKCxFuZENcKXHH96AGV4sD4RUw+XJ5rRo
cLIoMqEH0yimlJ9F5N0yaWhiUiWuiIGNSaNljXqKxEDuAZy05ol+ZtJDYpp5TexE
AwOcLT72kU1w9g1bk56QFrgEte+0hi7KWonHGyXOheU9Dh2NiQmuEUYQMes6nbIZ
AnVbziT+RvKucWUTGAGZ0eZjyOCThrd0WDJS1pDw4QNRe8bOE77D4IBPzDviacGA
dLkTkqbh6Ec8BiHxp527zzykh7xkIQBs9SetHsKqKZ8GJw5tbFK4e2SW1wJAaKIJ
82DCkE9NkZw4vWRah3oTzsaxJNY7UXKHVjWtf031CP9nlFKGZhPC8RBMh5FvDu5B
vtEQbzpq27lG+aQhTWmMOB+GjQgLEY+cnfNzEhu51Oh3ztJgHbA1qP3BH3mFzzn8
xvD3MXKldIOTw58BiWLo3l9ZKWCCPRKu5lMVnk55/6GIuNAfT7MtFU5zt1IeSU1H
i3OgIh4hXKTrAILXA9pRIpTN9WBwLEbPzIv1u/Nnn4E3D5lTgnsxDhUUJIOC4w9l
WBp8qx0v7+ZCwzmCWIhZgAMO+7ktPgen1u0SWjdZIIT9s7q8AteDYimKVTD7p/uL
uy+p0ovySIG//TB/3bKLQSapx7B98lltVIoz/BofkEjExf9sUkSAcORGdbi4GTTo
JXwdh+jy5++m47SJ9qYsqtANsAP1tWuk3HN4u0bUkRnBUqHSoRr0/UEDSd8nnnrV
utwLUWCGogWEeMZydZ6r9psfe4mBOBosv4/e6h+4POjd08yOxj/17MSoNzow5Kgz
ZKSgutot4uRdHysq9U/0RhcVn6aYFbqE+c/nCn2DffL1sKUoKqL+IU9sTpD+qVY2
KZBcRNmFNaqFVtlEJDk3xwmfGJiBwUBzX6T6BLowl3Pbfhw3zO7sdBh0JfxdNKmG
ojGTsocnXOKZZhQHP0mCEWm+joMYwmPUUm6ReqkGr7HFzhhQwA+Yk8ywtYnyXu/j
VvTZoZe9c3iiZP0AqpqKu6CKyr4+Yq/hf633ZNoyBPRhj5qN50TjGqEKJqPbKOo9
qaUPIquOWHXbFH3o8m3sb8Dad12JhL0xkDQfX0FvDtPPBM8bV9pezklnQnXS/wLc
79zAsP3X/K+eUOxCi8ZFdZVq64f+msN151wSv0yk1kq5sQLhxEs4yPUQvQPKtfkb
PL6DstH7c//AIrP0D7Ed6QOoB700iGVnMn11I6lUe+N80M17kNxxzOl+OHs97kdx
A4ooVFu3nYbq7NjdqKDNXoIX4nvvPxzSmAP6J5MHgtzYQwsbED11la+qodIgdNW8
x0YpYG4P4HugAleLa+4xC02rqp+USe89eiSYXAAJ2JEaBWr9vk00Po56Pc9WmMnL
Kz8aklrYsh9rQ7vOdjni1AtyBZGNQZdiUFTqcXNboPY7cqwHS5jUPTplqU5I7WkL
cfm+faU/5ms6wrtTEk/rEyrwEQHVFbKiXegK8JRvUfaYuGSfqDQ8js8yBMBzIQM5
49TwjDc3V12twYFPOCCsv9ssocn0rxRHOfs/lWusVgh17hRg18kGJJ4q7OPEsfHa
e19E0zOL718fTtUThUzZMl+6udn2rrdBG1tIfV6Nm69YqpHr1NUOEkM8/J0MJiSG
Nw7OQkU9C0FveWTQ9HzbNCYQezi9tBGlxFu6x5LhkMdxm10RrZOL8fCdOvgYS1R2
+n+rsnjxRJLtzBtmEYpav5xljCcIQAQ+Vv+LHjNIwIzWahQ8szaH0mIqwX9U03A9
T2eUOe584oneo9B+4Fk7j88DdaPJh08rTsZGQ91ISWbRw7P2JD8BGU7D9vfT9Ln4
Kk49N9xI2u9409D4XkpHGBu9oqElf/BYzDyCVTtu8wTU93Ktvy/WjM1xWMYgZ7Ie
FP4TlsKrS3zp9A5NdJ7qunjGf+7zJk8DrT99SEj8aMXX0iwacz7M+T7nOqm9uxcr
gRhtUKsnT8hG8mXRQbbxfWwmFtpvQF/RBgEcbjQCG2w+yB8d9HskLO4Zm+HQjGPu
pBxZsILLcgDJAAGFK8UuoXprlgIEkZi7XavKjrxaOoH4uOIfpKXbDVXpSa0XZG0Y
PD0Q+vGx5wk1dwJC7VOj1+npUV+834bwrD+KZbioU5gGoHyDH0L16C85BWkumt3y
c8ABvvrTvkBPiNnCUfUaZVhja1ssLJBGYzPqEnhnNPLmH3GKyAEXBtcu8sQJIEy4
qwPHS9WzmEg5TfPrcCQ0ZJTfLakDqTfcurhpN66BY+FiHI0KotEClzYlQSg5qhkS
wF0G8DVTq8OGKffXGJ+vqg6zflHBYMGAUXVBTLR9rXSKItbxdrfQQ0m9sritrNtp
Bn8VQ947SHkoOlYoWR4r6qhzZVkmqeYtKs68fa+xr2k1CSOPh0jAGdalMzYVoD/o
b0RS9axZuRP/rAiaTt84yArH3YiWHK77olSZAN1pRuABWYWRztHGeTFYnoMcLnuu
DCnSLlgzXtRDtcJVc43RZHRxhITEqbd48G1Yy8e0q4VLcAYMxKMmOfkk81szE6oV
lESaGrxWJZV/A34AuuSK9TvDNuh7SXn+z4HTtzhPE6nMPT+3RD/CRGvv6iLqTdU6
16Xpg6+gTJaIAvFyuYtXkMIIYU3EdVE7431Gh4F3JoBRD7824vMwlL8BX159qfCK
DZ7+f7yTxGlyHjoGlt6c2WddOFR0TpkinlsnkvvI0WxbT2YjZiiAqw7nDcu0j5W+
fm6S5fCiL2oiy7Pzb7KHx61Z/DmmvVRdSnxE7KaAkukKYeOadgDC9wQfHDKOsn2v
a9soNt0qxVAlHldegoPeiCGqSjiYZyHsBeo/9DZghFcsnlUDMCbg4Hy18cXG4TR3
ZOcl+/8YCoMK22UbXFy/wwb4v+VtcnKtd0Nwj3mfGfSiKLmBcJQHGbQPCpzQUPg4
qmNfNh/iiVzbXqlXQbggP5L0v5OB10Fdi95fmBOY4yiornbnyN2rpQVRghJGCy6Z
EZx8Lnjn50hhtGM2pySbpy4J69PW58dbl345+sWxy4BRSKtc16i8sX1gQtBL2LJg
Jq3LwrHzizCUJ28fXvi34DYwchRCWNnf7U193bWU73rF6pgcTeXVQwvllox2q9QE
Sloi1cKxaRTKPeELHqUGHbU7RchuJk8ocTNz0R1pC+kgVT6ojrk5yYKO/GgIjxry
iMh+SGM3Ljuzuz4FmqDLwcBEBPIVqoZ9hlkL/EJF+Qc0cn/JSev4uRNpZodNZsOq
vLxoP2ehHNFdlIyUk4jF0/6DUA9UfGOdsWT1zxoXpR9EZxfHzSHipjXcdyXASnWn
vJgly5cKh+jMvWQAA0JwHPo71ulf7TRw6XG+/qeazpLzqCFeH5/IUSk47pHzz757
3Vol1JalsrM1jOzc4RXPN9tcGbI+5kZHbi+/GxtOCdJ42ch3Zk25VsFgUY7U8IHp
iTHMf1YTl8MPbtKMPvvGLCX5k2EMr68xU+7tvFI8Yvyb24rFcw+28yAhgiVSnfoP
Cn6u/KRbyIiWaWOHRP2JEOxbmWLh2GmqOiTkv+KzTpB43WveatSM8GXtxdkxX8U1
on+bOAnAfbkZapHltiz6GVTEQ0M5XQBcmfjbAWLjg99t3OeCfnGmxSbK9YuSzSXd
D0GsNAZjWi0BFjKk8bwaEwDeR0M30b14YR3HIAKHP8qJxzmqlzP8wm6SE4E2+7oF
rVmrSnGbKH8ZG//7ZUzE0I2R2haV3L4A695eT+sePaNSH5gUqBKumHNKAQLEt0xK
3sOExkREvaNU507WebUmQVfkXaMJ52uuv4EBb88yEDuYMKYczxfOyGNMF833wI5A
bN04PUNnbGfYm+VTSjhV3sukvehQldv2mQBJYD111/z/or/C7cWlBhaw5l4TRA3j
b/AGZU3G9qripF0ii+2Q7Zo56uoGYFUTPKHNH3Suka8IEk+XXIny2lC93pm3DEiA
aaJRmfBeq/zQ28gfeqatOYUcIf/WLghSNX+w4nOJpxjHnxxwyoH+9+aplBHVn2Uu
kSKdOS1E17NUzw8TB8Sh1LJNBI2Jhlh3VJQtujjD6inKSMTpJT4lUV4dpL3BxM6/
772iee8jO1jHQCbQWW86faa6vO8L9lpQq1hTspqV5PbzzgPoeChYu9UGcwKMPjtg
j9+Ww+3nTSxYcmVLnViPDElcf6vW4Q8p+bA3QxV3aB1ZS7U5n8Jim0zT4ntvXlLT
v+n+IZPzAh40fUGyVto83Dqy19xH2zJax/YhgdNY+/fd+ZXH7bu7ghtchjaXvisx
vbAZdEMFX2rEg3vlwQKPtT7n11OKZFhUzNfb7kedIkzgZh0uapxhWwHVtP7x1B3E
7SzRG8ECQx7tsW5vsr/+EC3mHNligCG7w2nhixHNGSFU1oYXcBDah6+EYhUvNfkK
tOUE3JVvRRu7HQ0+yBV63lkBe/1PhUNss3LPUhbzHOmvOE6zm+CjD0180LO43oCy
BVPXLH6G6rfeQZnZTV8pQHQVWNRtAw4eHAKQ/nHt4P/v6n35ID57XGZ7C8tPt9Pm
BlJ/Oi5qoR9c/Nn6o2E05e2cx9s5iLLTw+zymSGz40gtKdtsnFJbyoA61mjgWSdV
N5pjpX+LYeMDAOW6u4eKcZxMWjf852lr426jLGQli/YxlUunVbz6suGpg1LqJoA+
IznHGM1MUPjXNqS9VBC/Bza/O4OY7h1LgNbTNHAvI1+NYVQGEwndZaSongjszkmf
c7j4Si/hYvxmF3t2Hrn5wbiW9Ei6Ufh2s/nLcs0qQBLTNMZ+DGM7vkyFEhEPm5NZ
Dcv9BWw0KylID0Yehum8uMzpj0lDdPjzcZvYVbBxYXqzs3SqYwtVdUgsIGmS/NV7
wJ6c8RQHJ8MO9mc7MMDR5Lk5Enwo9b2wirKKvlomdSlWFo5lib7sv3NfR4Yo4clr
UGNVxdBZgscCT6M2Jv01y1xlIlxWXFGtY9sxOODRn/RqIrCNMozaHWeRRZuvdhju
KfuBkX7O5dflq36WH2fYyiFf5Iol08q4+A2EqyIMSO0whw6pTRaPjGfBM/KESLym
rK4uiQxSQYZAjRKd6ebUWiCnSt7YeAjjIMVeD5qxRaJJrt96mTcn6m+OGWa+7xUd
3waRQB1e/VpKtljRaNTmgjcK/PFlMOkjATjKJzmQKhjQDRJevff+UK9FU9eAWZie
UXa2BIPiE557yyPuM+XhwQqpVOGd1xCMWJkkL1bS9Cn8FNlfls/vgMo2bsXGYkB0
cYWSg3pwsxMk2B3WhWwuyL2zVfAcxuwjgQugQ02vXH/2hBL1jHtY5GwFcRnLdo2d
EkUO+16c9aXOLseJYnXgFw553hw9/f26ACYqITJw5xP+XvljiFZkdSDJzTun/+0V
R+QopEfkXNZyQVkNPeYGn4ZgBhCVViqlDmVliavV8qhBe4X1uB3lxERM6i+Mx5S4
/DUlKFe8KFR/bf1f8Lxwmqw4rvcm/CbEgGiaZGShYFs34dLpEsODaWVNMwfgT/sR
+PX+5U1PQG8yxLRpZ2AqDj0dcm0Gb7ZBMlAj4h+I451k8ia6oGmNeOPeEVsuefMF
1f6Mr/L2vP91gJpbSL4OY53QwgEml0wGyg127/9cKP2gxdQ5ZIVCCDNkpxtcMdq5
f/Ub9Gnx1Vkj2MZDoIuaEUBzm6gBPBLiwTWrb7fQSjBW70GkBKjQdvEUTBpH7m2J
MSXU+kmb6it6UetGEh+9FueNhyAgNDO6nOs0T3m38z6Wgo8BEEooOLMDXlkAssJe
Z65eipxSHnM1ykITnlsQUy70iUlGqRrI3c8uAzmmI4oV0xn1/TvzQeGu+C8Vq5ij
L0uXXTSVLaLlyhzXOy7wP0HSiAtQvC5piFOeh4fg39VfXeTb6RFeXtETHtZlxX9v
CFJaXpJOhtIAgJYUclFcq3cUoVIMtimlLk5Sx+f8EnDD9fIrDzBvT13iYOcHYT7m
0batF/Vqx3SIxDCUDb3zFV/ZsZ7cLqxzpYaGIb7D2kOsO/SNHApuEZ5OOS3fEdIC
Gbas1aGQ7Jb/qZh1TZwaJcMmIDdPYhdK9MPiziZWqqwW8cT0k5jEpnU5cTySrrx4
yTZJnZ26bge/LHOfUFqwdMTaKUIbkybj2rgtCgcNvA4R+UNBmJAA5ot2Rhqlr6os
dFZdR4nnNumlrDhQS2YykQtbufgwr3TzE/dYAh3dAHNWOdjvZKWRxcwj0TFdMUc4
Za4olUMttCy4or6bsazvbLNMMeVe7FlImFQL3iQds9FBRQXhT5apNDCEkW3IIqpS
N2xCpTVfbV1oQ+FGsS+0yw3khxeBWk4GcO9y1iPL/gCWdZP/oackMJNDS2x37Pxv
ftpFlrbWpmrp5GAsPBXDPPEUplqMgY+iU1Tflx5YfOzuTIpYIO9nFkvsHMW5AXOm
UXvtWfFZ62BUKunsjWUvDpDWyw/MXJmkZ2NTbC/WQHiylVcyz9/OjHaFP76WHePP
4SMn6C2OIhohRyoDEQdjb1r3UeflsrpLz29gJu0vU3ziPuFh9M0yoTlQGpuhaQB3
/lBqML6VioNwp2dngsk1/lcRbgGIWrzWUKILdsbbZC6owC3oMnGkpPX1JoClRKr+
ZaS1uhX/9Vw3gsiIj1gqdNXG9pxZc5nsPN3oO5y7qRcQHoFzWe+BhID2OBek5P1O
8GtPrFYtyaBGXv9MGheEYdn6M2zmd++5Zm8VB2Ml9pAYmoJILzj1Aq22WFgusN4m
+PGVna47/xNh/cayCIJ1Ih/Q630KF2wvo5ti+/6siZGTLtrhKk3hYGl8R6T6ov7k
Qje1TsgJhEBh06B1lHQ/Kny/sg/1wWekB4IfjLlsbIGSjXA0jR8T7YcpbAVHalKa
2ickfPv7FFOjr+y4iHRI4DFcH1tgqooKQkdsLL/GK2Nwz1qssVskbI8hHjGGMyxU
aDYMf8AdxZARJ0Da2uely0UE/kLYinb4Dp5R3pHJinHEQsj+eryoyaYva2qN52JU
UdHGCsPz/pS2+ypHzyq4Z2h8tS5ya7TC+fh/eQs48YVXupVFPcq/c6S6ccasPV+M
H+DhsOVUumedVQiQAt5u6aL4Z4U8No0wAS9mDyau61Az9rJQBXM+VUCET3lFwwlJ
1lsp7/dAUM0xSYNvjR1+NBAdX2XOTXN8zclp0hTWtw22dRP1hCW4ceQ0C496vuUB
IJqWDJP/rgOQYaosKEnqWRhhG0N6+WgeWq73O49jurQuH/bpa+UO0ubYtq6yCQDb
kevk5BKUFwePQhfJEeSGpyyaw8jc9nbooQ3PeM53B/oaLr7Hf/RJg5Pf54ReCWpx
5r9A/jArCs+9wUuPyRfauOxrjMkVmO44zBOE0R3rpP8xw1sVpkeO4C2S2Hb1ougw
cbxRYtjrSL37bEBzZTcFpm0BD/zWHaigpRPhudl13lb5/KRtiYwxvEz2pMFRuyEu
6sOArXabonAJ1isWS4cnEF/qWoLkXkfuRsMJxLMG9fFKZnT0A0fuBv4Z7CXMsAHe
RYU0H8VIW7jbafB65F6hVK3qx1d3ZKSTowK4ifeIZc9r/HYk+BsMQAxOripCc39/
xm6fad55lJFTQBSvyW5+SqA5vwVPTWW5uza0pTkFEPd1twAPa/JYSy01h8YcG5pO
x3u+MSzsMWk/yUWeBNRnhLGSvakGLjE9L8APkf7lEpnHP6PCHmnrF8XGCHzo5rTz
nNAHXkaJt8KM4gCljc6ox671IcLrkTTLW/bqsPevDdIqKY45SgdYttYlH3oxKYPO
noDx9l+hFg6Gp7NpXqbpt+Cm94bne+GG+/kG5gqzn9yJpsgqP1tlmlpV+sfELo5e
Olgu/611z+Tt4i2GQcq43ihyLEVqk9b/DL29CuV/gtHvuYohBItX6d2+UAbjekKL
b8LkN3HHDKjGYPbQOaD8C1v2kEvkqfajdvxomZwShfS2LE5mhOwM/fa58yfR3hJt
KdhIZLaiOwVPmLtXk+sJWJ5GFLNRs/sg3R0UFDFV7mSHtKcIVC/KTULlm3MA+bjx
H0hiBh2A+xWXMOLqDwcJDRI9qmGntEnjp/c+sVf6zyG+i8DS4kAQGXSVoVsfiK+M
z/L6y67GptTi3OK1kC5yyeg8OJBwn4woBvphajeO6LjGvUSAtUzskAsJR5pzYwXN
28SvMvNLvSqAiRmev5MNHnmGfb5b59+AlH4fb7knMYP10ECV6yqGgIbKg+6zbBY0
shBH9nkICaQ206Ti+i83KdiVRxhmq/EMMNrtizNHOEf87ocEx6nU6XDbQ0ZeVMYZ
G0HtuZCMEqJ+OWA77gluqKq5gmXN2utx/alRpvUP9y5/tC/5nPc6c9zQKYxu6rhp
rQ6vM0+8Iq4oPsFuUxWUgWcU//LyUP7Uoyo3IHNRMiFBTIpEFMWU1wajQAcgwtYY
7+BpmqImq8KxXxwJaiL/MxALKEXX2IzbUkK2DSHxDaJ7xtSDPBZrgqtWTttk7afJ
kGguEQPPriCEd+0srKCSdffTNCHGHifClawp3k5wlnZbMnAyitMvFhm1RPJM0rYB
AGdSWw2DxkYu3XRRW+LcjgPnYiGxZ4dWji+sqg4Xf/LfS0NxTu/jP/4WKx+oc4RW
RZ3Hx60/mTO/Kix0uKacymg6eZC3qgEa0oKsr4AMDX0VI2+5j9SimyglPZrGZ1nk
qZWkaqG+Zp465raCdGn50SwSnIPdT3/Cz7p+sfaa91XC94X3Ekt7tp7ute1Nkn5A
MQVm6BhhsUlu5/qEglgKVLDKgRdgHkko7hqO/RUoJ4sbrm28r/xA8q2p2THo9M2z
9iWrA5StwWjj46fvQoJWTaJw0+nWsAwY2JWBGYQX/inog/O8PWi5iPOoXmiw6FI1
Z6285FOOXwbIANTF1VoWlwjhvNjcjha5FSyhw8tf6bFfLbTPo87mpnxptqtig/Xw
Oe3XQqT6F6fJ8SEx4AZULQ+clxZj1gYiVcW3xyHHWrloljksianHJ+WeBleDfbQa
M40PD/KDZESUijWLyuH2mURV2Yw8lJ1GaWdx3R+en/zunFq9Mxa9lIziTnVYO6hu
wwkkwy9MueimcoQBTblaOcmdphu7LsgFqGIg9BMn0CEUNtxACXJuemHY0p2YYAM/
inBAgSx8tMY/oeoS4QMHu1AJwu+u1iSBD9Z3A7MGnbmYSJiziT05xCLG+ckSYiNI
1WiT7wkcRyceYW1Ru1gLfxF1W9e2b9ZapNgzMnUBixz/tJYS1azcbcO7irpOcSpb
BBTirJWHm3HUDOqxn0dkc8I59/qfNE5xroaTVfZnri4cWhR8T0VrFPlo45nIHvxs
NHDFDSsd6DJalhtlseYZul8rHtvwwxng3De8I4G/5VRMJHj/sfuLV08rmOVm/cOi
UMOBonKIU3b5vrzOezivhPc8VMNi5Qj78/TTycpt+P5mcqQ8pxWT3xAhGSYO5/Gn
J6tId4me++dX3i5h021QHS+mAoowkcFQ/ClqlNfxxH9l3DWKLHT0MuGfuv9OeCV5
AtpxVr3ye/PDemY7mqOINhPOxUQlau4l5NMpLwZKoV8U9lV//mZTR79dY+3GQEv9
YHQIIpTbhm4ghKJYMPLtv6Eqq+mDSU44OI4NmFeIzs62LAAc4eQZJ0kbR18nPUSk
GUeagDCMlezrBSznUOYaQCsyZ2Y5yov/eI5nCesN8Jy2DkqEiN2VfZsr/UVV4Xzr
X/h4bDpDJlqs5aZxmtQjtlV6VHBnPU9usX/RjilSY84pCcir8Gvn22RhLbKRzXtz
ASCXLlhSW8a3Y9H42JCc5iGDGzBKhfOvIpK/vMoPpANEsv0byuKDmrJHcxVyEtON
cfsJvBRGuRX1mM4stiUuZk99NKs124eWU7tbI2BXJjEGhx4MU7Ajb8jv2Jjyz4ae
ra40gYNPsN4zawpAGkl+lBi5FY3we1tD/eZRamb622+vw8TN1fG+ZOKyOa/vlGLf
D7P5t4dr/f/0AYxsnCDfLrnMmCCMlk06WkXuS31Pl1VciyHopLqzw9ZFH3vkuGLZ
pQhJMJytGHOOeTVphh0rE3yOoBHMFwUfwNA1pUXzy9PnNg9ZvGGDv2EDWV+wJJ8B
U1xIMdM2B+0BgOync8E6QXks5uxgr5n5jXLyPX6DAP8dOxq4vLEQ5rEDKzLflyIj
/HrfX8WoViIx8P+/lLrV/Bt19sPYensDUKCB+5lj5IMlA6QfULGfxKBy63AQ8ZvU
a1LNLZj+4a2QH+DASWNp2o4FD1690uD+Noooqt87z//8VgKb1Uyj7lk2IZYct8nQ
3v0KtCCW7F4ixG3dI3fpttZvtUakGEescLjxI/OU8anTo6VELWWbHxSA68QvBK6m
GWjxQJbfK8VH+FPhKOsx96d5xtBx2/1XrxvDeGU3sdY0Irn9gm0YLPZ9XdTfVLdy
cJPWTdwVyZ2z5KLDcJDu5FUYJA+u8rFrHjkCfxn8JU+c9G0wMhQrkeqKfvng0P5L
NXrQLYorZXYabw8xXq9y7Xs5cb5sxn+wq8yBBPYINdNK0WceVnbB3limUzT55VKF
GCKgg8SczICa7feB3Wb1IKPvsTMok5upLu0mWoIlcus2c2BZ7dDeJ88dOOcpzxCf
XLk3pycureEPPgs1CmxggZR9jnxFDaGjsreL7yXqHYysj7CVFhgxVRmoAbTXhBFH
D8L92WtF9qvqFJVooWd+PTt3K8rA8dzwV1MvHSnqF6/9NXsl16e4+v9Pz3LGYiJ9
ci6JDnsSS0IM9GO6rJzRJ9v4gNjjWd8Kmgu8hym1VE3KdMofs8h/l9kOFTdPp7vO
HOIEPn3AgZCVaFzvBN17vInRpS9+d3KanDwplb7Ia5ejo0p9kZ1FZniq0pX9XkRS
xfmKfApAqLSbNIQgiLLC4GAsZ92TgMTltPO4M6L8FWB3eOSAUP/inJbXkwlNG8t7
wRB6aywrz4yRDVYIgZgaYo73NnICqKYwUJVzWh5Dv3lmhTKZtF9KzWF6aWUZAp1D
CNFx5z/p01aW4X7dLezyBtUQbpZeNBfKua/nJ3nZ0rgs7cSNiQ9T7D/2wurSrNsN
atQ/8NR+8Wabh4w8M1+2ndFs1aBVEAqL9UN/FA7expvtGVPKRco/NAh0PW0iPiRw
3lbErceff9C1pl6PzcEKOrsNzfHAk2YiKWsteO4hEYdKpwrmnIZIn83VjpzM7VHd
v8Artfh4AYzsSKwRtGsv3xZWKlQ/Vgq6Pj2ZuWFkpi80kKALgeVihrtc+WH3NWQ8
4Rd1r2aeGX7uivTMPgp2rFmji0llF/JL5crsdKt6aR+fXr7dN/vy0QC+PNgMLuF3
MgojX3SkeTuiIjnwbyenRFrXhBOdt4crp+e2NquhNMTa9tCg22s24nzRGwp2UTE2
QVzDVlbQJTzeKDA0p1eZ+13SptNPHo660psymsyutd22Z4ZOU1Jv+tIA4SC8wsxL
zV59xgT9JRDgG92MZV1nTbLIx7Di3nflETdWZsFL//AgSq4lAaV1iBGbUW2Qp+vG
Rxcemf7t4bIuIKoRpLqrdZ+snFYejKoQTCu3lawGIqSctxHK2u4XtO/bdDsIseys
BkCDC7kMYHCIBYBEnqOxQHsJktVM8WYiVdjUN/KnANm9u1P+z89tlk+qzLUFgTTY
SuuR85mai0iiZbGaZ5QXC4ItoORdI+wEC5fmrVrMPpgB0Fhk6Y+piVVwGvf9Cm1T
Ur98yArBhKvhnVViMOU6E6GbMyxiCnOFXhozGeaHDoidxhd1tY91cRcDWnfP+KS0
9ShWk6zRCU8PEVR/RU3P+l0WkRTwnw7co436PdmOFFXUvTff2a4Od2A9DLw984aB
SyIk2Fn9iI34GlictxfrXb5fD72AOFWFLqouaO7/Tcfu+9UTY18fgBWvnCIUQDe9
gspBjH4mdCkHQP5gYvS76ljbBmC9cwQP1ySOhIQ7h40f0PgCalsUtGygXIKFPM5I
12QRQtKDQpqy9eM6qICr1bm5pVjjNsI0fWfUHZVKf8dsfv7ePOn64tnAegsZofW2
aawHRm6dg2bi5mifXvgDnuEWMU1j33k1eq/A98YubvuUIDPjpJTlENx5O3hbeqAI
l9nA2e+eo+2wGDbaiADzWE/HN/G88691JizxQBVow51nQ/xPT6vSdBwgVO+shd1h
6U45jSqNoDtUPXIa6VprUGALZTj8nR25ltp9GHFAlKOTeAX94d/X6y3TiR4Ox2/A
gbo43yuOZ92aAz1IJjxdLFc8RY/9g76h4KpP8nr3NPCDGlguMrfBhw7NyS90fM0i
mwdRPbH9ziXytdRkMIgFt5JwEFeNlVKGbydpIMTSx/CHfAJcyYaF5uo0/BZdFKb+
/ECK5edRarwiXCsDMmKzP4ae8cLdKeHTL4Fv5XVau+WfOlDZprBdYSQoeJ3C32Ku
qqaGo3IY0Yau9+uZ+EG5jnGxFsFaN3Psdy9nYFDrJOUT6DCAw/RI85YzDPqZhA54
aJkMxZ40iS0xg6IcimZRWOD2+qYmvmKyPeRlsDsmKoBYYvRjP/M0mOnM1UsqYREX
Cmeb1oCWxxXyRRemCA4nGh6mA3xDh2ooUyMI7z49JK/cvfi7QjZqFWJlKK/nF3HB
v+qONRIw4rBZV/NuVPySXtoBmJIqUITpEoWjp+bT7jKmxjUKiY+DSoF5cLT0Ey/a
I6uIS5O5gCLDsdFg7xDQKdLj0XsMF54LWZpXsnS/FHOEm58E1MopcWKONA9TWfu6
ITmjSQ2MbwEL5D2DHRlpm7DUDQ9fdu8ICr3JJOsHKORFtYxnIEZbL1fDDmLP6ULQ
/9lP7wE89ICrOJo3exADawPUR3WW9Gn2aF+jhEN4cosc2MYbqsQqpc4bfZq0a0yl
TIIQ23NrHH92aLayCUHSZaJFtsA+3Ni0P7eI3yivmty1IFkYZwPH+6nW2RykY4zT
uvq20tKEUR4+zVKhP6z5yVmnJKYWsM/Sp2Buyj9XsK1rOunhmZANjl4EgI1lk8/d
0TOopxTOsIIqKRvCuXe9dGC6tbJrVngjRWRPW9xZbpxbqTDgeqNWlXq4QShQ8kiz
mu66t+YjXHiupsGjGh4E2lr4Qj8MBv7Waja0zvhNu3v3lts7lmSD96H/uv0nkulj
9A+XyZncF2a+yMI4rvkV/ZypJ4SvIrWWmBZEu2uh8vW2imOtjUq3gWhDomAYMWJZ
VnnO0f37mhX/Xv0+AVQZIRqPTqzZ7RD0gOWalc9S6sDJVWVIbBojO/i0d2LsMT8r
N/PlO9ZBslmeVk6TKH0bTGjQ1YTmCGS5um6PPnFGL6z40CBCs4ujK7eabY5GToSP
wndfj/JzRhL8rzsmwguRkURJv9xxeVyu/yQDrxgRdbu47at4mVGNXDfXlcA5JKCG
PgSI6Xx02sYCDBhSi9XoCaWcmBtGCQCBvLBbVfYyBNQCvuIyyKv4rSapRxwBVYEq
qEJV/bO/+F0LB94x5/fE91RhJwMO8LxsUoXUXsrxbzK/QDUA8Pqqk35dfOc4sA7k
vQ2qkyvtAjf20PhPPeJd0exaC12k03JV3OLkveIO0ouQ9Ucp/KnI7nJwcqplOCRh
EVOFvX7MOWQT0WsSJkFun3XpmJ4ufXmJkca4r8vNwIlfnpe5ss815jDR7IxXECUv
F750w4Lg3vmS0aofItdWETS3pBr330KPfjs0z2u8u2dcnot+dIBPwZ3ERynUp5mi
/DjlR9ub/IxpyihICFnqK8vzLBz05SoI3fR+WV+vF56f2Xz54ms0S5Ss6zTe1an8
GX836qEZ4sReToSUYyPCJL+AnM+u0ulJgSMdREXiHSYdDloaAvkxCw9ItdI+hd62
cItTVCJ7A43Xk96FyFlyHE2Qr7wRW9wc7VeIQDsRu97vWzcn5+iV3SjQ5H+ZoYJq
+lOiCZK7ZBqaocym440mjCOJ1Yh0LQZRx9g+tnLhbboflV6h7A0p7vY7z4aOpH1z
LFm1L0VBA21jiK+jxhAbvUy73ye1e6k/gE4cvL7h1zjoNB2o+L02lFlqNczTTsGt
ifZxkaAkplupZBsTuT4GgrQK7lrjfrXu3o+cOVPw8FD6mNqJ+QuIWNth6fySvR5M
BMpH6vK7IoPKEbpX6Qo8FxxvbVpfzhSuooGjY+kpT77YnSpOsMrlMdZITAtwutho
s7FoVdR54O8vh32x/yqG9bexkp5ARNmNiSMVp/Iqd/mfohpjt7iFcX7bDQ6GbM7M
4F5xnb8AIfXycXoyMO2bsjP2qAFnuVjmSxw9WjyQL1WABrS1omO7lxmIU6fEZaS8
em7R5imJNme3muqN8MXwQ5UoQX7rjmig/HwkM5DN8Pf21CsIaHUa4N/3RSsmyqVk
fK4T56pZPyM+CPgciTlAZBxK61CkD4sdhepkJtK/ygao4BK/2x1PyykrdO2lhUPB
Z66IdmqD/oOWJvNapSK5kalze/q3h8gHkT5WQlkq8PDc5RQnfFjVaDZKJDh8a/Ff
GcHxzt4elAVMEmIRRrmu3a53UOEc4tPQ7OdWSR5BrkrkWm0YkzBY/0NtdvlHNfrS
yZVqu/yShRbF8jCQe0R2lt7boYRRsxEIuGzlZz+r0Rj3hgymeXe0BVniA15P/B9l
EKnjtGSWJD9l7uDYHlmAo2Ns9Yw7LCYgE5gtDh4khjbwaI/e7qLxEDSAcByVK8IY
pXGVfVwJ+Uoapt+zp/WKSENeBFevRLInJS04ygVP+Im3iLUhd1Ue7oVs8wj91T4e
3HSyhco5lOR3MmpEacvOtLBZ+FbiErhEtlYPg9zosCwdBcs+okvfOABcm7B/OOoE
/VK2t3Wu7QQEG86aYgeZIVtwAll5hbbuLzwSEsPAHCvLGEqeD2Oy0aXFnxWNLnyt
9XDNdIQSnSJq9PhTVPG1eOm2RjQZ1C3NCMLOFVK4mWwrbUaxM+LqePK2DmSEHcXX
gvALXtQFCrx6WADdkmR5ZRUXN8CzSk9DDbh58Qw/nPXCCaxqoKOV4cH2GkpXDo7R
vTVQSsx34F9g3X/M4k50eD53kZNtR0iDHt1jAXvgKpLiDT2yTXRDeoukdcVqFdUp
xe+gwiSumvulJ0r5k/FaJJlsn3cqebU2HbCFaHuJeJ8HqJzx+TDdbH/6L1+32/ut
iPm5LTZuy2buUyhEpPjRqR9uYNeZys2IFnPzoe647TWqe/pjzNLAK4Xs/X6BsNh7
5RofC7SnwhTv0uzhl+wEC98N2B0qbZ+i+cOJfOsm2Ik64BXgFqXVYmQxyZn4ezXg
agNxb44WX91vQiHiNWhbZsav/lW7A+W/Ncwo+VNERg0ZU1AqWCmTByCqrhHXcHV5
0hZVjyEfUF97LAkurRXR7ZQpo1VERFfO2m9zUoqHeYouT0HfDyBozd964E3yM6Fo
w0oJeAuOxyLOQB16kTOlElwbnfY6jq3RQ11PA+cgxhOo2yw80SLNn9CvYLg+XdUK
A5pjwBVQ+LmMW+Ha/8adWCdFraqjstjq5OQFdBrckw0853EF/1pPgfdABqmhzI2A
kG5w9vmvW67imQxe2M/YQu+LD/yq3pgHhESId/wthTP9UAwdp8UY79WBlbI5VpnF
6GtzsFS32wummJGaS4vbmB/l2EuXw9sV0TwrvrtNz3O7K90EAD59TReGcrkssZR5
XdUdU3xIV0KoVhPuqfRXRfuUEkLnhOtEYScce5jaHs/ouVxMd6JlMQv0vDxjSScC
CgR1i2yhPQqbatYkga7efEQgZsncf3786hFM+M9PFCWR0WeQloM24lpW9UBjJZHq
D9zarLsXaicStFQggNmqY8yls5VM3JkfCjadmyREQCjgOFpl+ivyNUnJt5M+v6Co
Py1Kn1ci/iit9cDeNiLZBl3qRCulJVklhLN1fUBlgrVa035gnwRkmu44LtkLeSlb
uIbFWPfQb8RY4kZICfJb8cTdM7e+AQRGShI0VkY9+thT5fKMKjqW9UiVxxKj4M+J
R33+/GZgYgJSU2tqLwQtPnQPyWHlyGNop/X7D02zqaeJD8Yzfbc0/TPzNdUz9irc
wWd5EnrJv++Fj1cl9eRqUGMAb1Zu+wGwjhkKlcuHyJl8x9E0AuUzW68V6mHpJjpq
FnS7NsgT0Pi+XjEdnj9vNfSjy2XOS5Z4NAQb4oIOE0G9plax7KiTSDyK2Vyj/RCl
i8mp+EqJjjx6fz/vbmWcP5kz9MsUk8c0hVpYJ/iT6ocRciM6ye3ZAmzDQufKUXUy
JXRzgOlieBRMBGa6h+QBw+p0hLsBuKc9bwC90EIsQ3blJZVsS6uEuZiAQxm9bfwV
rocPb4+DN9pwNgkH2PAlITYWAfZmOBmqlqgCczuGngwEIoGmNVuN1vBrO+070pA2
cxMS4xUC2YVWWocxtmK2Z9AgKtnkxEvVo5g93j0fYUZ7/h7n+8UyUtc7+blpILEL
BeEBVCOxYzucZz/b0kNzBmVx1q9QYqb5Cm+vqWU2maEqS5cAUACrczxawey0rMVq
eMCcjoTPH2ugcl7/8f9QUZK5GEyLor+Of71mrabQ813wKn15KpZPn7gYP0SsY7gH
0/ldZc+npwzVmfsmOOvhslh2Q0Bqqryhh+cenuE81xeT+4cpVfud3KEVH8s2yUsR
dEVPoCgGZZffVViAdRAnKaAx7OUkomj8iIUaDZebH3qp03+32NM0yHGeo+CU7rwQ
aTTMpi8jLjeZRQ9ow55nLnMa1SDtKCNQVmPT1XNH1djY7PdrQ9+IZlV0hL9FZmYT
og0slYo/BkT6TuvozOakQ+DdJQLoUp4Hl5u+mGGAs85PF06lVwMwtf55Qt/u7IFC
PFUeiPjiO1+PXA7wvQvTaiuXzir1FHoh5Y9s3dq0TpLv0EPGyWp/r4SEJlekv/au
wN3aW3Mj4QhzBtnll0l7tcbauNcBopJMUt9zlFU3GJO0TxrkutckJ4AY1PAlemJx
uGYlMji3on4tqqOFKBCLbwn2EFHPou18yFX4SlKh80s5XlS/g+QQNFnYm+wqfHnW
TQpUez2st2Ngez23RPCybct+a4wqyhdMMmCcm6Ydxn/WNuq9zTlPD3+eZjdcDsRv
KOqaynO4BuoIYWhcU3iHN2shWkDRlXggJlB8d3EncOUx16cB0v1UmWu7dQlmMCto
LZDdS2Y3aiHKmRnfUexeMpwCE8nEbXm7PXddGbscyW4xrjFa2YJOAprtyCro2Vty
xS6y00lrw+sqoZw5fT50VHPv1NpMk5FKnJOyaE3E8ZoqfJyzK32HNaRYiZPdNYcJ
Y1Oxjxr6ER7o+s+2IJxaM7vnRxH6RysITVYDwX/l+mMOcwcKFLfijaFiArxpkGQA
xoHaA1A9QTAoYUG6hC5SSjKobVBQN3L7GPVSkq03WQx14IEpUSsQN6CJA9+wK5Zo
Xo7fVOnMMld9p5L4+WQ0yw/227Y87D45RgF0D7G0z8NDaKoEQdisj+gHJ217piX0
yAbQHZFB9jp+iLuCqq1BgwiL/DjJnH5srqCy1CMtorASqVRp3Yw+RX6CkeZVTIgh
zRvdZtTgc7WzrayVJNDB1CT58Zoc8sN/3tMsTQd9938D8eLNOOYViaMNeT1YzyrA
gbfbgrYamGSu92phkee663JaHmR4abQ4kLF/ssMtp9X/StOWR80t/RyjqxzFJH4l
WkL1oxNpGZO7Yx1N6TtEC/Q+R98MoiOLg/LIp3NEFwI3Mi0sqOQo3cCaAuKkd2dU
mOxbgkb25VOsKfYlwATpcReSDfH42ORxlTxiVRUg6RhKdA7bIM3rQg9S/xbrsQ+A
4Nr3B+foFvJEYldFdFEVLyFd8slLRl1NAEHzhNzIpGq+K8Fx3ZZ/6EndbdiR0qak
rB5kayeuG1qRcqGjj8vcAweywvhhD8pNjR6luHBLk52w4lKbdFUwt4RFSHpDRCAn
A8VjhNNgitZtVXBi7eJ6Dr2GNoblRo9Y9nFrUlrtbwl03rBgqAt7miMqWdwBesMl
qBMzX9Xp9MfddjYqqAT9omM4YUBAvf+qQx+S1KjR6WlnY9sTiO9P8YL4aIhNgAlx
V6czarTpsmVaKuve3ml+DbLbpxLoN+PGZ7m5dnoYt17wsitS8zbjZoNcqrMYt0b3
qX7naE+Dq0+7VQwfOCJ1e6tgRs5YaVoAyKY9S26Mo0lrFpGWIjqu/DvzM5NGfHER
yelB1hcRxYL9eioFIc1t/PW/Ziy2eqATDBybg7jPim1R+II0rzvNRdO3P/QifvUe
X1qgRQGGebzoWYVkttfEIvVZIQld1eTO4SYPeiUXDS5heAjTgHkB+MOzMw7MNzFN
zLr1qF2DHMYGSEAZbINgwBboljrX7lw9vRgSa0xn/785c2vMcmTw6Q1PRzxoDrc2
1QFhbfF1Q0DWH3kAYOE1Ubt4QrKY36yQzbzc8N7K1zu9E57KGAKQu+0sropQzynN
ECRZMYdj0sgZXdsi/CUVvQ3hFMltqgtLWvhLjnxoY7oBdcLnbER1eoBYMTGKhxVf
xf7FVeZN4nBxckvM95TndKqUGaV6PCzN42VjT0HG3UJ44St6+MHpjE1XCGHZDBNd
3/8aSFTaZRSw+iJ2GCszJRNoRXUz3krsUD397utqEKdM2z+BGKvaKYRRhwP4+0lC
/tcV87LDcC2Iu9RpdOJHV3XXeYwSFU1tGbcZ+/e2gOlGjysjcAXHqQHqyT0C23xe
nUDlJw+hStlBR5daleko9Olc/k7G08NsxGarSnAo1iBJeLU2p39Mkd0knQsYukAh
89k+Hn3MA2vx5YNtXTx12dtR4RgwA56J93S/+z5/3sTOg8uJne4bfJ7Oy1KFqEQI
9U46zfBFIPmhfeA70OqKGrUMnlc6SOQtiD7s0D3z3Jga7JX8gZd/zmQJaENQ3GTi
4uRNCTT/7A6Nq1KgcUtEEYmQfEmAnPiYjYiJkF9TXLIbgLp1M8fUbAX3bMKkTld3
qSkROJC36gPGmq1Cbh/odq3J0aWuIbzO34ZHDlwlB2tP3knJfzUGjboaSQr/9ttB
U5XT3pty0VNizKfjU1cfXjlDoIwd8hgMjh5/MSvn+dg9M5ElU7d8+Tlxga8IJW5x
DPszCR9/F61CCKd+bQf4qvSKooZZc8crdG8II4GlO5g3aPJqqKjVvo3P1T5CWd47
pdc3v3zXLvu8YsbS93LQ1d0gadDFFEkSNoMpgFy5Ag7N6E/GQLxEDDIgcGK1qPly
6vAevZyDhfD8PhGj/GcdvbgHvdGrz+Jo5mkLBYXpDARHhT5fAJrbTBg/wkfcecQC
a6SfN88kFZGJ4t+S1TxkW9GAZJu8SZN6o4v8+jqpD9YYPBkqaEUT7la4ainenJMo
nlg2UKTcxvHAilz3/140OPVOgYq9XKcDwTD8Q1vlnyGjIxLFqHOQuhcXyb4Bh/ip
XCY0KCgkeLF8iQASla5O/9cUf/6n2UpQs/b60Wu4mvpnhAh36p51xYFX7ZpOz6M8
IojLCj5cpNI8CAHMQ5NggYPJhQ+xSfp6RhC6Fyh1tKLpsjqzLyTIlxOsBswjfII9
aKe3icu5osIYYq52rEPYiSO15nYIGwcJ67Tchx1MFD4V0SIOTJQUpQ7F00lcztyv
cDKzoZ2kfBTBk6s+z7dlkfNUeit9f4Huo6JpTcuZN8rDi/djjI+42pL0rsmV3X7i
mUUmPVcCmpfiK2Hfbe1flleuuWfv9qRm85uENl4c6Scu5sdJodDdpV1cLYQFZBO1
7k62VL2TbbPqwV1WYqePBhqZQVfwnuZiWsnbcecAzRkw14PFrrD38cj1ja0qUkak
MI0lSAQhmAcy2QyNWy2Jt/s/bJ5AK5EwARajuhQ8052UpxziIcwsfa80Y8nZk/bU
Ul1UFXJJBmzxEegk6SFtuf0WLQm7j80rTfqUEPbFP7SDw5+H1CpM5ovljxA29077
oqPzu66s56DMqod/3h1zZrHkZ+L/ogW3ZWfBhXL+2J4p0nHBmLilxp26/bFrNwph
B/JKMlzd4nir1n61gUn4EnL2CQSnBjPhmiOjsxEHZHxXtC2Nnx2BaD19CJVtwQ5o
ot5ggP9WqkMV832nN4M6qvkIBb5HN/fo+3gOU3OpXWpSd3eYOM4hnBNewlF4rGtc
8McS95J7GAuUSkuy/7iXBAgAXX7BAWE9Pq5ZFC/fXfOW2alxJlaHAssGEWl0iJEQ
YlVZrmitbvU2ex6OXBg2F2oGH81iZL0staBr1hJrdrBSk1rrSeIt5xHwBhaNEtx9
4WL2qitSaG7PlV77aNHrN1TykSgljrjszeNdeJOZhwPD499NFheBh//3CoaRO07D
B/CufCEksCXkZhGZamfmy+oNdCDhVgiOYx5Ag6UJBXRUnjZWHCP5YK/NR/xJWpaf
snZkCNwxrm7dzEGDVJhjPFpOdP5dwQ2SNqw8mVgk5gsrrkzV+/afnxhFLyIWz9Ml
OBbMpiFyqESR13tpaUY7pjEDu1Np1h5E0NepBTbtZdy0YHcBy0N/ESj279GBx+Iz
oiFJ1f/v7pTsZ7FXIVrW0VICTNd1vQ70Cglv+N68nTkebVJs4czvVKq6C1rklULi
EgTvru4MgJr53O1cQVQYNqSTLm+65M0K//vXY9QAmKK4lGrSO4LwAQSQs4phNFLZ
ks/HA1OhYWTI/tbxf/Rpwzu1evywfpYLpNf8Ay33BG8ov4W7QAJCGXaO2YGvcg9l
OjRmrVp5eOfXC9ISRBlffCJxYlTqk7Wrg0DWrf3+kkuo2/9y2qsmJpRjg7L0HkT0
hHuviJFUcq0Ior3l1RnBeCgiRBtxVFm9GGOCeuVYqxzOdVLrx5/hd13MDtIq17FH
CwadhXbjLD6hAqZiC9mTwP2BMnnOvXiWL8/0azIQAIuvEs9hNyGthriGGrXxDZkp
ZxWjt/M2Y4wNob932ls8frrVe0WoZByPDV3d/zWlmuLPLWYWCONJUWMg7k1UQA0V
PuZ/AlJPBkbObcgKpQIdjF67K+mwhBRenv7au+ipg2KePCaLATMfWTSODcwE1kSE
Xa+tJ4nOtjiRhTWbtAFscnf9QLcRE0NO5XGGZY1tlaaqIX4KzORnNUqbKYfppGpT
88ZmmyHMhYQFklwHb8pKGHEQ/Ni0D8JE2hBSlc6GzOCZ2sOc9C6r8qDJa69nzTKl
fTx0NdEyCkfpjdBLkw0m+3QGXz2uo8Hs8mZfvVeBTEzUaPCtKTtX/iRJhVkt9Sun
UkkYj9yt2Qmj4iv4PyEVixmBSfd4lbeJzHSfEQLRHNDQLuMtyYZGvbAjBfTSeaDi
y3DSinqkP4uAU0vc1k/hj81jYIXq/7KkwKSbK44ix2DVorECSRbIfx6dHnJe8k86
+ERYtQd4lDftgzzmfznsijGX+0+jBZ6GIodjQDuG1o/r5brjlMYp8XFelTDbKyWA
QaWTNG/7GRjF108aS2vu9wFHx4dTq6qqtR+KdNdVqs2vrrmDDt3AXssaBpE0/3eE
ec3+ZSug9HOm9d3QwlmmhecIGxWhMbLoYfARCUs09dxOZk0+swxkvEU7KvCjm+uK
pTSvIc9Uqy6yC48I/S+WcwtqGxd4oDPuikmPkgmLPddMxp2ivKHFkOGy47ubZUgL
7bUCmeN5LSTDee/jZeWQIEaMPkfQYzyArkmaA2jU9WzS8xipf5MxFWLWrpgL9a8S
Q5K2eoEX265a7BoeOSq2dSiueJr1TjUw/FCgb8l6cHIIEkXKSjuFfVppwPKxz8D5
Gc0qfR2DW14CgLEHbLKeMZpyl7Mh5NJ4PZUxJbKTB6EYYX9qbqZ3D8C3DHOxMus2
RCOulKEaucrjwQRbOH1bvRiaqUWkDMk/fY42G0cGc0koDvOhuIk3EcZEJEUBUIgS
L3gGUmRgLkZ0I9z43FbcmjBNFSS8gisL0slqZ12cV+K2gTfk+/uyffkxKHCiqIN8
DUETH74oTiGe0Y3LgbymKld3q1lgD6rX0p8qB4Xs1IRUDdPzqjuirsjJJ4OkldkU
Dz1jxxV9XTEQz56K07U5C+tUGH7co1AArR5AKuINt3pQANMlvzdalnKs8COJFg6B
JDoYRc4kpH0xUwksk6vX9KBtgKWhY0aEPM+nyD9uaWJCksYwXYx8dktmp5tfwQqU
OHVj84MSgCSlh14TSAqdPWwqS8jr6NjXFWpVctS0o4v1xpi5LtZPajqB0+oeWJW2
/AjEyXkITiiC0XqpBFLTNkoQa9s/KJFWgvO9xmg7xtMiYCIndVdtQOqLD4xw0X9V
L0JvWMhiQjnwjawaQuVcHXZv89ckO0AqykkDvoERgCP4nkeWGTa5RKwKNmn0shMy
TnjiiXmvcvY6PGztjr5vLYdRPbz5TkyMQRbA0fmsO5iCfWXz/Ba2Xy6LvJEKfY2U
orUR+OwQwBXHKZR6yaeSKHcGlt2G1BuWzL17+2xJfO1M4Av0Iqo/V0N8iGHsRcHI
mEDQFkym0qnGKlN8Jx2an05TPVbkiFxkVYHH1Ju+HKm6sG2imYJt2TkBCNU6IvMT
IyxMuUZIKxawH+mGBJjZQ/FBXmFs0a3nxHeX2mt5LcqrfzNKmWWQQDV1WP9eWJio
PTQwDJ5UdtqnIjf/2KUlUjB7C4173LWxQ+Zz3sNtS381yH7eDWf0aQ/Yl9mhCjdm
ccZ5Htf8x8PBdwEEq4wDCShAm76ok79Z+CbHwCUZcVsy94ifRnx8dtwgicN2BMm9
W5SMTYJ6zDA8nwbXOECW1R35hFlW3lmrsg0LF+EYzoFHt1bXr0cnVg9eXqSaGQ5E
1ICiWbLdKtkKC5Or8mix9rkSKYKfrLaE0Y++bllHKnsMloMSDkx0QiQ2UxKn0mf9
AXxrEmMuugjg0DdqKu2v66CfdCOz/3NP4AO6FYDQdz5SdLxp5HKhAd8BxCnsg2m4
YS+xEeb8vxM/rj+8fvvx2Eoc/YivxwPBWt5ttLoRxHgLr3zBRLCTUYkgvOFUBAY9
kd7skUe6SMgs8H6sqwOf6Og0RYqqcqst8cz4x5d9ZEgwzXwUcw3bMsRgisT9Pz4S
WMAujk/bTpOF+HXgfN/eYLAWotRXV1pMb61paK47v4nyGOGth4nXez2c8nw4Eo08
c4QfbWe1XnPm+GKg0OD1wjKmhGJP43aSm7Gqw481jl9Lufj8DKpD2N3o9TssSlcH
hdzQwWIYj60Fuw63xLIoXFuWgble2wRcJBM/wNkgTN41bMOTeFk6yaAgnTKHKPWS
4bXf0VbAb8OTHzULqklPjiKT82rZ3lm10VZjeZc4TH6cMg5b+LCVfJKaitjXojg0
SuwHgfz63GMIXHeksLeMonNIFG3lbB8NPmv9BbXWzf5Y4+9OrKnhxhTU2R+XOBlO
Q2JkSeu0SFfNa2y2ms2P5PplacnSVIuqiDPY9wU4skrD9K32wJw32Wq5JlKBlX9z
v42xiLnwbkgI+91U8QYWFCnyEGixYMdNhWrcDgzsqb4ZPlwQQVzmFdNSNNxfVuh+
IyXn/ynLSUHohp5jsTGvpJi3r1vg3EI1Th+ywYZqE5ZwPteuNOA7vd3tSk5UNYDE
DPVcIxfYmlPIskoyb07wDb3xlk28bJ7yvF1+QsugZZJknkuN8D0n6V/odafnfVNc
RiHLMv0namzjzGsvZ8PZtEPIQAQZc1alCQ0yaKv/8xSRHza1MSO1+t6yKef3Thuh
h+cNECMhXgNkPbDrW0tRPvodebivfg2sniXF59sP0zdgK7QTMGjJr1+vKNobLeXj
wzYzhUrU6MCBpOm0muO8DXC4119stcAmFxbjU8b1T1bsrGEHY37WnpKMnEZxqD5b
xoX1JFJ0XdzCc6iK+gsDEpWb2tsbbg5BTnA2QVeGpxBrBH67mxaOdPEFijNy1J1G
n8ugltR4I5vs3gNC9ifatqTidWtPjd0vitHBnvHDXugNUpsQq7CA0CyMc5jI08tI
ezdLUryu267I2SnEKocxb36rH0k8mLdjojrcfGJTjnHjqfj6LAGFCRa/c0GOBv09
Q8kVo+/ubEUWJK5t3VjnJwhH7K3pIUN6O490QJaeasgMRFFuG31EZuOnDp0NLRoy
ogv1Mc/W3ndwLBzrQMZ+VJFNl5BJF6062LsKj/BQJnFUJOTsS5UqCFJYLaCMF2dN
VMSUu66N+JTViiIWLHMaTT2zS7H/OIJkvwUefHJ2iZg3RNJMbEe8AsZ9KgNclgyD
Y7jYJg9dQMr14J/KxgZnL1Mrndm26JZa03m7AdWB3DqHHMDZKXoqgz9fBuKL9SG3
4dgC/JWP/s5kyoz+QHVfn+hnVloWqKjyfRKJqXTCG05V9WYCAivZSJllA6PzCdrI
7DMUtfJDsl5x1mLa8DuETh30B/k1y+ZJWXLHD6zDO8MrpYqj2OLGovNvDLEsIBuG
1DdUVAFZawGV9l55IIUe14AtJlqLU2ydXqosE+p9d1eVIkNkOm7K3mpT87ujuHsg
SM3AGRkXkQRcC3DaIxOyhTIrSzX4gCgAvDWdBo/WfC6ilecW2n7RKX4gBSAFJOHP
BTwS4IjFEbutrgbnmwYkEQl1uB9aOw7TXLSk0wx82U/vsX4CGPVdUQ89Ev69gl3l
iNq7LtSQmFxY7TjgsHO8iNz1Lu8QyBgKYtEdUqsS9fDnj+YhlY+YH2u+NLRUTYuY
vvh5ZJMLwvG5C/0eKt+sNU8wDVqJPureVtPshjXfYTUfrnfFEM52cmwclbHMf2JU
4JiEa1Yk9R9hywPq6+u+F47YJZxetlOrHWbrQOt7jhwcx4ElS9gOaIQMxkQ5qYAl
uyYFtcnPM0IamZmeAKbJ7N/j1OujcKZKbTRYoodS1tvPuPmLZ6jZzAEH6HhYV4uO
1rfl1i4LOw9ZRwz3OKLE1NULV6ieQjonD2JJ7TdjMrBraqMQ9PqxqkqvcAzkxOxK
6i0vAX32FLFNIsdC08rI6hn4geQy4Hq+EPxFgiyHcNSo4MamldhV528fjxOuY+vn
YY+DF0r9KnRXsE8ZrQeq9PhQTX0BbXOGUiuqdrfhp7tAWIkKxZzDA9GJcMLDcP83
t2Mdo8udvobJ6Ud6T6G3HKINHvlnrebYNLrfKfBMH8kKhsrsdH9hl0jYewjGarta
oaH1wMlWhjaYJnsxbF1KpREKGQj+k5Md231CWfebmJ2e5mrkQx5/H9QVJ/PqW2Dj
0mulZWWXijdHN4ZjeAHbVHkvCZ6rTX7WxqQOKPURcHsLBCac5ah8onDB6AgGeI8b
jqjNFu4zzeo6Thv30cNLB46qylmYZ5gDXrayIHxzEyDEd9ABdg8Wxnn17i6edDNw
+CJ9usws8fyAeZKU/YOvqIEoU29N7IdGyIM0adFrYw7BqZzZqpYjsNDD0npUDnw9
cNKYFZ3uYThsjPu0TY/h1Zi27g5tnLaSSPYlcNPw7IF+pUUDN4MV26KRvw0MJoEq
DDZJu8VY9z4MYTH1syvR5PuRtsCXgPj3/YcCxfVJXcUCvF2CxDegNPcWahO0N26S
N0YZwTfV7lJjfmriiDmZZJo0mWBauHQrU+mvwpqwTsXwsUyGYCCACQaferb1vo//
AduU++vQRNghqnpMSEwIE2uK6VT24UdZ7zR42/mr65fyUgV8JlCtiKV8V6eWxU8O
aVVas2rByQnEI4dFXeyW7MrU9Ys4OsykRVjUUdOciRrxMBFc1VpEJ9d7ysvNUYW6
Ii1wLwOFcvuPK5HSvEn9NHmfNQ25r57XLlFUbMLLU01oYuE71Rrpa5bt4OdoSalU
Su6N4GaJawXURN7DqG6nlGiL4VLzKK+sbri8ZIWJ6SW57Zu+dj/IhUHo+877hiDe
UR4d1Qque3cmKz/VCC+/p4EIuJ7OouziIyI29inW4N2BAk2o0M4JUF8TDP9iSAdO
LZLnnMEYp9nJlVP+dZfO7X95624LqJ5spn4RC5Rg35D4ar8lHBU8sWqQLspJiB2C
jhsh8IeAi2qwB2dD+NUel/0c88AzbYtoPKMs6I8DJnlvdzT/6/CE/QESbFGoSisQ
8bZ0JVlgU6K7A1DIbtNJ5/mz7youpm2Ai52am7HC+QE9S5fMp5c5rKYsKB69NvQI
0Hn3LZJpUHUy8F4tbVN10O/Ay41V1EmwLYxR0ahMuuM0Si0ghvw0Lby1o/MG91DC
B9Ff7rJt0tggZ286JROM6ieU8iWx2kdGH3sXeirxqEXCsfyyhwxAtSdwOv9yOwnf
Np84QrxnF6yKw3tPhDz9RDDs6+zbmCQbMtsBPesomC3k2Pl5rG4YVBgy/m93+8gt
6XlGExpCmIR9cp6vD1/Jv6n+7MYH9TKQ4br58JLR8Wvb/94ibqrXrmMy3IGF6opb
iiJmrTpgDj9fozD16I4xLA6i5KqhtDQ4Y/ym8rEVW/OzfJ/iwtgtgYrgZ5bPGP+y
BOnnFqcLLXtbEAHWDnVo5F69wa2M0ERMKwWu/L7in/STi30EanZearm+PgpKOjA6
+Jbxmsb0mZytTntIEpijjxKrwSfriYeid1x0uppUY4uXaih213LWN+hS0dmRgp9X
l41xhOsFii9ZAJ23fSAKDXsehmHzkzD9IbKbiTRzKzkj8kW0hPebS12Si5o8uVQA
2s4zFP1nnzDoCeih52HUziXuuo+GFp+lETMC/U/mhpCEtmRUsCDLqKQ+8F+JaROk
ZfNYyFIAUDFvGD3hs/kGp8ucs/XVRStCEcREZzUIXlSd21zXB0WPzJ9UxpsNiHzt
CuE+peNlZHI8yytUPBUOCgc84Dnhuyk5AzkSU31ILwn22QgoIObdqWlAPuST8QKk
YsqPn5gzG4lD1JPDfmjZwC2yoEuErOIyJNiJpW1AYf+4E1oBESigBdig3pHuWaNl
1qmiqaEFqQBBygZuzryFgE4LHowv4yX15piFfIWDPQxjpfL4kqzASnf4rGwB2Gry
XsAU+vb5nwcGkg/M0sgP94X32y6dgNQadH0e0t1qB03OZqBNikvsdUKqw1AC0FfH
PNOh7BUcl7cFyKOKUl06RwRvNUgw4Uw+6rKtlhywM0Lck0KdRU5Fj6idy462i5ZZ
mL6rZ2MC5617vvcJXD60mDeOSgxo6yhQTu4tUdNVTZEIAdiWowL/PQGk9Wk3upKq
za8sNKGtNQI3Z6fyoMR46D0aq7cq1MJJHcwhyj+LpV0H9ZIUWBUaV+L97mm8DSbh
frCnBjIa1iYbJ6XboHoXBTznAFe3Lz4uV9zQwFJaIHN+KYb1UHOYVg1b+YSxL7gQ
8n5e2fhfeurqapiQuDH50Rd8V7LZvXjbgQp9tUz6RfLT7urM1KjpEMdU3WGgAkJX
m4mKG1+4uk9F8igLHULKuqDbS5ApmU0N1SJ5j0V9mAeAna+fh9Gp/4/T7CgoJb8E
xfMOZWsTnjpW8ssOtFlUu8ueUZMJsyniLtz6/UtVQ9A6rWT4KBxrVnqWZ9RhMJ34
Q+wHv12YpJcfMqJEvcZ7GsylqvEeXz7AP7Cdpl+Rv/Om/pxFS4pbz1hJY+MMSzhY
YpKNbMNkznMHXBuJQkRuxnOL4hBCj3vK43BVuDj2K80ajQj70UYaM041TJiNe1XO
J2z/ndpdum/tJG2OliRlrlr3ldSv0V00xtvKO0O2ZlBAGbc+F0qaoSzD24tPBFKF
wEuygBq1AqFWmVji7xMn6CTUyapTyKc67E4W7m19gk3660T7OkMag0mf4Ner3QtQ
FXzxX+WOrBZvs9xdNoB4LKwCs2MY2eUH42COJQHy9i9jjyb2ANaHZUis+YS6tb95
WKm2dCobT+rs9iUaseF05RtDu3VMzJjb7dba0GlIPnwiUevPX+GBClWSSbdqtR3J
NYmNt6u2fVyFjS6SQOv6ZYCEGYWrcFAEKtKIfiDYOGe/gCT7TJDVgok74HttRRZD
A3j3tBYZJihPPDa4AMH7P/8XpRmMtnkBoFGUOUBiaw80OLk6QXF1SYDtTctPWe1h
zgn4Wv3AccpBltvZpnCS0gIH3YQ11RLwlNZhtFyCPWmvO4TOyEtule3fvMOlUGWu
8n8DQZG/jMBZQgSMZ7Or3rFKo7XPBLMaYAHjCYEBx+FutO6xhJ4RY6mGtiff9BgF
r1a9dzfisdo7hMDnRUH8Phw5tBz26O174ZyOtmf8D/rw8NlWIFDNOAVswex6VzRn
SL+v83wUOkuit7C6XJGrlz2fQRvfejkfXLs8fsYgTlu17DD6SO0BA0idRVfoR+hK
xfyKmYdKgFJGSZvQ4Y9mncINDKMlQvT2F2pYvDP4TqV7hZl27YkwgPZ2mVnC3oS5
WVfC0cfX2LzDA/1bdW6P5negeD+pddX4tx4+hERKp8e9I1XXSMZRffnz7h4xjevp
G/ilIFNr/zGwrcNgfBXXO+vix5KVgb6N/AuxNaeCK6YMxgG6hgI1FDc5zOQBA8em
N/I4Hcm6NHw8V5T5kCVVcHlsZ5YrQTnfS6kNjkRs9AQPSk1BTuuXjyjLy+rxd2ss
w6hpxQ1M2jBts2BG/3UTpwoLyEbCRVWHO6aLTCTtbYJV7CbBHMGpr+Ki14cDfJjW
Om7mDTny9iXHhJUmLJL0ftGP1CE5ct+52Jea0IBs33RB00xh3onfwIC2mE8YuQXr
sCsyJDPGVG+FlEKVdCEOCUoZTqCc/o49AbJ9U+vy76eMExzGxwA6QB49r+b8spta
becyK5Szgppsg1UvtoHJTZn6Od3XitwAtLp6ZrVRF8+5arSej/rQUtGUoSZsaXU0
QgU4Q4tvydvfVWUBUoXPceK7/YCYUpZBEELVZC0ZKTvHe7F02l8FsGl2N1LVaqF9
6MKsnK/TVCija6g0FXuO4hldmDmfrx39FNcDdrw75yUcrHSd4BXl9zrqziQq9TCD
xOraOQdIFkkgePz7kxd4C/gLorq9nH6oVTlcV/s3XpMk67wQ6wr2eF0te5ktiyB3
NwWMoF8DCTzxRAzVioCpwIAFUW9NQO2Yl0IHP2QLMllWS+xUMpGIEDYOouKuPVEp
CruGKAMNTPehgsYct3s+xg2zxTzj0dB0o6/Thw1/bhxShHTOMsAtEZSAlzDlQ6ds
pvTUX7yATvwjASwbsCiDlouvYghgsczMcNm7Wq6wl5WFGYeKeoosERzgM7ouPrID
uWzeqR5ApcVYqYMMFiKdrVSG8U8/hWZGPHpUxEHXKJ2C77Ckg76DsTKXssJE0+mQ
2ZGpExUV2pbfP787MEfigSo2aLBgbfU+DBAOcHuPwEC35PoTKq0Uwj26y3WLaht0
vqbGWFgamcyp6J9Xx8pLCoZr/QRjZJvYlTi1NnpaAr4P4TCoExCA2kJlDdmBX/H3
MIlCQWhrom/Q13fubb1jW5hc2NRx9EB7YvH09NOf0VHHg/kb+QkpACc02xcxpxxs
uNGoxG5Z7q4YK+hMegXy7h+e6P6RVCELZsVRVl771WiweiV2Smm0ZLLF8gosh/d+
27PTvp8TckCv/5VyejI7FbnYRwDctCA+e6Ogfvg6UVRmZMfrBuRQvBeaOFNT8kYU
b3Hd8lSC0CGhjwjN6rn0Eb/DaB/KWdi0tgBrN6jKSanBmxpFr1dPO8QtqI1WcOOQ
zs/Jg90EbsF4OauSQoc9oWkDLFNiKtkGxwRGY1to5UnLfj2q2YVUuY0DP53B/ezV
TY6mhnz/iqNnpXvkJ53HI2tLAmSgPkOIyj+xcIUQIe5oW/ek4fcWG7ErHYTJMrGz
37nvrMWuTi7MPx5Ttz1ss103x1ZWgreXqJ9Fo8kUo/jfDaKHDJnhcmbVXaxCOYPG
KFek0/h7QGMIapSWBpp+4g/HKOpXeLrJdNBTaV45b7urfcj0FiMPJXAUmZFHuMCh
8br7gEW68fMiwGKSiPGim5HNHILiWt8LVffsGkEn0oLPnO7kWIyyGaLC/QCqBxC0
V2vRUE5pNGqlq1QKdMBwPNW5FWCPhlW3AKdGEu9P1XfF7tGykmNErsIqCq6zrF/J
B6GI7MArvSuIi/w4hZNJSBQrbrub48l31RZ8ZTqWr2EApeRXIbU9tcgMC5HOkyly
9fiVeWjHcw2qi+l6x5C1yzJXKv+N64Ig4p5bATlfK5vk56F/n+GkSu0Ui2od3+dP
l4bj+lNJb2zSBL9roqX0rRw5HechIeYCulaNamOB+bM1YYfRXo5WXwctIsLZCpnc
FvDzgcilPyjwdHOBAHcj6DsnRZqr56fx27Tfc8tF5plJt994sDO6UpsXi0BQGGVV
xV27DYenJL4aMcSsN70dGvW1OjkFDpq8K0/z5hhz/iy8KfYMqsFcAr8BugJSQVh0
hp6N43Rhwx7OA9qlLxTOEZEIYqzoWoC82xQyBiwQPtOSIfGnHU+UUQnBWmGbzax1
pEQiFmKTIPWoR4U+DVB3ZR2+FCtrcwRxm9iOTehNGPFoYxXQYd2tlIk2d4UcUPTU
XxzF5B09yaxibaTEgfebuoHr1UN+PAxuhtBXBr3Oxxj1JULL3SnIsM70nOcJnWNz
lElo7QvDA6tvliF1McqQ37x1kkvJIZlYgnQJ9AlbpSomqnjL9Aqll5AI9wFOuSmp
bsEJj3A1M6g+2CxBp20MlDC/6ae/cw/V+5ApkdPVjdXuFElMeLk45BMbB0ki2NPu
F6Imgjk8fb22TeiDo9nvecGA7Z1zyCNAhSSqTz+o3Bu4trLRl+EtxL5oJUrFug/K
ns6oYCVupXYhTVIVdUNhrtzLx6CaLZ75nzxVkrVDsDdx+D69iSTE7BUFqIeyyaok
LQZDMxoqX5/mUCKC867GzICnVjDn1VUn5Yam3KaeeBiUD6ONZ+p4913qbQbHz4sO
MlhQb+cien/DmUpXvSlKPUomFQAKjzzYZMTwjCFszWM6RkIxuIn6R2iA4kxGUEUB
lugZflupVQ/5AsnBLvqIaGvvTdqA/CPayZBk49kK1E7qlap+ONxilMiwAVARfdzK
1CmrUMC21NiZBr3U09l3+BUIdMjUVHunHhY1fbSsd5x/xb53ktsloX4d6iFY24SL
klwIZxE+dVJPR45ZaTFHXacOKNzmQCpUQSOK9VBhlVoKVF+2q1Bo7RD2fF15Jw0+
/EUmtDUG88JnW0PEmNj8J5dwRvShzym/aYtM7VS3uAD+aLb7NaRaCtsD/mZyCK8Q
tsReyx1NtLLO5EQjdGqVROeHHdDKoq5oI1HgbPVcrNyjd3HAoWboBe+KX7JO+mmP
l/jxNQtrjlCO0/eyIA0KFn9OvTt2IPEH5ULbFSKL6p+EDjGZ14jTQvvzJuOwl2k/
yR5+C9dyxCb+L3A7t+IuxI6IAPi+8oG4jgxE68Sa1zffhGD6BHob9GOdYrXbmhPq
a30TONqVwh9tvrvyrluGtH7u7jV1se0xLsaUhCTs7cWOU3MNAcVaSQ6sLLDt9G+v
tpPmVAJdrD2y9AJf7JbQpmW5OhFiBc5wNIW9B8th5URTAPZqieDOuqFcRqnbkwRW
EY4bN47ylwbo4DNF9F3r2aq7UZQiOg/yJAMKWNtsvBQOJXnIhZU98I6YdzrNMGrb
nBHmD8pMMmMiDblsJsPsjFuKpO0QqmH+XD8Sic2huYPg9eP29xehnU5tDUJWHMkI
DoZoVNOJv9B/QnXMTqQIw7i0TTCfwy+UJzfPPX+5oNyrQnuRaLaAi2rKBemXwnPq
+A2JPYpz/UpHpaitH5TaCWwJfmTJc9ZdTX/LDv/domjAUBOcU5Rlab9FKK54+Yyk
Qlo/LVxi2ywBcD1sM7Dn93VDToQgdSlWG9nBRTX8D7wmBLS+hCsDq3/5vK5JdCcl
iJZ1P3AuVOO09NrkcX56RJ82kyD2Qti/HLAQaOqx7AAQyNxnsJBS500NJy+LCt5v
nXFJwr+BOWmny5t5H2VSjkO598Wycq/fa9HZdjlBb8MsVDKlHL24muoC1CZwIhXm
3/qzMRQsIGqASA6+7ySZ8doUmnpAzcexnfAmpXaI/6qzQOPxltOTN+DcIQNzp/k8
2QjwcbqLkKZZ3aNKzIV5zlYuGk/lxLelWQ7Zr1CF0QeBdCYt2kPpK+kK4y58ww88
IbJQeJ0Clw8UCzfrsVRVLYth1agtLNdscpU2HkjZqYxpoHeF4O3/XJLBdQtHGdgC
0F+PPCOjfnK+s2djOSCdFtfYWkkCPWO0gwwTPx1e7NPCbQBnEz1qaTFwZYlPvgJT
6avu3edIbGxglKfqxsLkhds3EZMJ9ZCQ5VtTPxOvM3oLNodCPgtZAYBLcogsuwiu
aUpHhN7n+kFFEBZqLR9xtIHSWq64k4ZQ9wArM1FVXH2JZQzrQ9HPOZZCwF5bdPX+
mz/egfFIWwsoWT796ESsqsRRodAIISE5gD6x8UD4Bg7CUUVugLg3hgltUOgJZLr5
qhDoFDk5Ly8myf0ljgpSLFcrZEdAIRVV/OEsXaO5nqDP+nIpte0Foix132OZ0zOu
/VjB10KnZQHWNcShIFSMIb6QbcRHEpRllk5tkhT4R4UHpEkXtmlq5/T75e37dFbN
m5kOwJbL0Thf5T2LBpO8tsnl3MNkGS4Nl89uDDXxK4Xqhke2Akq84Wm9SQ1Zhm/a
L58ZfOlgMxCbKnGIX0pxlcBrA0SmUE3l6YTJQ5Bzx+hCWjDw3FLL/Y8bv1pYzFaP
y8mG74yT5LSTMckiij3hlhTWr67JRRes+Pu6T1tU+odA2jC7ozEELY0iC65hY47O
sRTE97prCk7sL/nEOh2nqZHHFnbww5nSut3hrkSNw/64bbl5pRwMk3TRbcUnNDNt
4lmmYsw0bzVymPc15WOhlv/P2bMYsM/0jTACutdzdnL/CeH3xU8fCAG1d0RXcsJA
3iYDj2RIbJsBafpAlUi0oMVos0rJPVdyYMzSjgcAXj5GASQqsrdqf0juwPJtsA/Q
dW0JVuywOqllcrXJSInMHx5Jt4od9alGt9M2wJFK5uDZn0diTWLUPur/3cS3TcTE
fMVyD/JHP3dhUQkj2S7mMBNgLP/mnta2ZHcdRHlX+gnyFclkmt2dpYxBZWWHEih+
EFgCeWGkG+THP/76n3my3ilgPqSzkUQfop7Qg5sq2HZju1xlzYF+yfBGjQgQg5Y5
Pw41v/fAvneua65uUEwurQGSGrvHbwkCYBKXJfx8xP7RnW7kddzeuIDV+fStO7/I
S8KBCGQ5Tjq8gsOmQLMFpG/xGBvm1zkGRyYp5pW6m9xJRVCkD3yapUbYXclT28Yd
HBk4IWRwZadRGfsaYyQrejoVXUKCZlEZdZ2heU1zSBddnq46O12Dbnlk1veX0lCM
ue5pJr791+rOtJh4fiL+hkohJ4PjUWkG3zRWnQwOlT7gw+uh+2V3TDjDjChWXNdk
rdu2Xa8OPQ/CcBKU9+NziZQHjkjlxiigveLk2o3EpMFPwY6ZpfioWtFhlyf28Pvi
A5mSIiYTIeCXOktRdjrt9sv8x+NJaB0n1r6Ucdn+2F3ql3EL6obkYCoEY1VnGYST
JqasqRXEj1r0Ym56h3BH1+QRmAvQsWlbQ7KR81niLoj714mZJRxvNoaksZH2pOrf
+zyB8Acij0+adSa0VuA4f0c9Jm2kDAxydbHs8KVu5a9Z9ygO4hIR56n9PArE6VzF
CkxZB0zMaWoyXVDrtkEFoO/451HMRfkZC+Bz/5wwemGk9k/d3WWTzTFFM8r3K5cP
jc8kpB44eTUAgCE7SbXSLBlLrdcIjjyuiFpEc485JBxQBIx0qHVsBzpSvtfXP/LP
AfLWtvxWtGdM3OgzEHwDiMDxU1dCqENxGas4Awlobt2JauhY0JKNFuajpe+UlU+e
l4a9JTONP3Du7V0SWWtCuFxk8Egal2QT324Ntrf+y8Pqj7Ay+4qEwMGxFvznYIB4
ThOaFv9JNmenMHv0p50HW2KuWz2xpGLe4j6BxcEIMPwHW8iBttNq/n4z5Ie6dq9d
bxtiTeUcB57ZwYYPNtnnw4PdQTfSg61yv+PE3axypaZ51NkyDUqpJjnwAt0+guec
/CV968GqwZrTj0OsgKvJw7qZx2zvQ5h3ZIfz3Silaloatnj8uW80nikBAwpjhNuS
5EkO9azvNO5Y45XeNKRGBEvxGC/243DEwo5AcL3mvfIY/8OvsYl3eaw/RDc+PpP6
XMeYJEPoKDAcXZy1Sln2p+BVU2JQMUljDq8vtYGXHh6Q/d0d2MAjhiSeFSKMTJyw
7jq7sxQi9tPMEs8SiBOcds/cmEkYexoAYbSm6EdLKwrIwHcugVZ0uN1ilwqep/4e
8AZu7wBoyUi/Ew3bzKyj9wp+mqxpdYGdhamg+8q18Ou/9Kuv+FXjDeq3WCGs4of1
XJ/J7I0KfGVEJH6vvtZ0ZtrURPw7kfKALeUT0vy+CPsgRVqbnz623tAZL2Gx8tbW
+qcjShq51kxTBCSzX+A+yOBoLEy9W2F3yYczyZRH92yz4odPUTN9kARtnir8E7zR
/rq7eOOupDZ7D64mi3daE7bWcoxKMB/fTMEp8Pm9jF4nCgk08MSRX9NN+JppYVr4
iV/efwt/0EjbRv0+y8cGGsreSp98Hn/RtMwsVHD23X8kBbxCBPC8BtzLFKQgOlAO
VyxpZEWEEfKPu0W/ifC33JBEP/AiLONTduQrOOJecQ1v7hgAC85SwdgBaI0BznBm
+8fIE8mn5rpA8jOstwrj5wPL64O/2gvDNOZ7dqNSoGoGaHpDgRYqNxChl1qTRe21
0rsh5L+SHInDeSPt28A3wuo8O2RjJaiHZyoUDmrQoxG0wSGDF2yNNxy3B4Z9C/60
LC6pGjHvgW04dfqurB+K/Fp0OHgbQIPTrqpikD2Lv79iBq3egPfprY6qRFEaPSWe
/Z3CGn8DrvQAT0U6efJKrgvhBNrjFN0v/k0WWe7EYm5mcUnccHt4CU36i+NPVLS3
5ExnFcDFB7GIT8TUYXoeWMotRLLH8Ma2EeDYOp+7jWkx+RvQIM97spPlR8+3G8K/
5p60VGhTzOGsWSdD10bmlRQc4bjmLITRAVLHHCX6iHtSq1mIaahVI6lKfN8Qqhrb
2z9by8CR2tVP/KSryjJe6pBgHQ4xuIWDJOYeoO4AYPv+xHVRfLBYIwLZaW5HTmV6
qfpdZ6o+gh55aV6PNQ0O0e+SBEt31YzDrDJrjt6lRI3V6z4tzL1eFxLRGtuTwaXL
fjf6/eSNgYaeP25BcIdSGuweyUp1/DrDYsQGoFE+Jf+Os7z3m/g2RPII9nk/IeWP
E46OGEmyFKUCcOl5zQ0y13tsqSJOn815wm6GvEMH+2KXcntQuPcPszDaEUI0C7EC
zx9BCmSidLx3Iz5A6F3Ly4bJOawXc/Z2fGlqNmkOYUPjWhW1FpZgMJpp95SPU/6A
AlkyTjKYnf9vGm1WrvKmpEh0v/qxlfnjkGg0XjY5W7HA3RrGPE9Os28NQfv5eMl1
kv6yy50BbJ73bmChMRxLdhiLfPOtUFW2jc2UDeWosLfzmIAIRnmmgZXSUfR+Ygmk
0jkwU2239fdXRvXzHMF9AHIaE6AelXv11IcrTyAkFQjiaC9eW6EtDcFouS7Icu/o
ZeOEJVhr6HISoJGJ3XEVj5LW5quV6mkr1EtHDJDaDVKgEa/MPWbM4VOYmO9wIvu6
/q1537Wabrter58gLHWXtTJMMnCjYgazsU9Q6XQW9sGowG4jXbP5uHVua9ZLYpNF
97XySvb8dR0tPn2yH1QPO59Q30Y90fddU/0FPXObdBf2kaUBpAmY/tGXY0b2hUOk
pd6rQmoujINWDVAmybUyJvs+y7VO1uGpFKmRZj9v6E9yGFHwFKDHNMYurGZ1Xusp
+p7LBVyVUN4uEFiRIqsgonZEWDAsyooJHwL7ECvqvUrB9IumSSWF6ISM0FownpUr
GFLyMj54eSlzJxVLziLBF3gu2FR0l19O9wZl09RTIHKGaGrG/wvXw+wvI2539zpc
K+Q2LjgK9joV9SKwu5TqI6Wo8E6hwBRSpmYAAQ1G2vzUxsAad9KCTFaKAOQx1l3R
kLNTdht+WysXFjB6h8sK9/eh3LTi6oGfw50t9YZ5G21d66UP+TczsUBXXK20mczV
wCRVKRjzoLcB7XXDfARQYj015/XgHWpTmcLnZNz/PD2I+5hrEhu4G/41mbEMr2Qq
e44AwWLbuaEh8ttvt3MyOAbiYO8Ilb6tx1jgIPeHWgMQB0eEv7V4nE0zdFxuLJnv
/Kmuhl5giO69pEIzTsfaYjnStPz+BwL6G/XbOF1DK3ScRA4Z6Fth09vqqgmz5Dj3
9dCHQjM6+VVHapxPCRGeU2U7yhmYsE7JwPdj8cPI0TjX0nF7LJa0KnB+6BJuhtS1
tnllGuEIDv6MPrP6mvNIsphKshXONNeG2BpRp8X1AfRD9ZIkxorfBTqS6QUB0mPX
xtsiFRqY7u5euRSCzvOfrV48BSI5z9hGVtLBU1Yfn1vyxYUPaOZJu/mQ70WWmiwq
1bXJaLa+e0nB4jBKvTVZmQqvVfBzzppvCv/zYvOjndroBg17byhsqKrdG6sCVNnn
fUbr6/RyIC12MMWL0pH5n7hwVTPOiYVzdRgnB4pjqlr7FzbvUAKOQDoapEuoeBRE
V0bPl57aWUb6CtOgvtAHTUSzxu3prw1TVuZoksbwHZ/8b+VSaXNRNurq58IMhAF0
35AYQ0TloNajt5UbosEviDvNGuvVI3ssHG+0XWN26wyREuGCBa4QyFiRdHMpcE5W
ZnumxgiJhwO34eFKjj8VkpvWTm4LvFrcrCYyu0yEJRAWvW6cvy5PJARlC+SJQOqf
5Yc14QLzXLFW9s1aKX4ZXKJBI2/k+h0bnJ47bfjuDpgFN+OlAjurVdDYYs2TBybs
ax85rJL+IabpiLEvmOztrLwrFSidY9JPiwYKmC7Q3TlQy6yv6Dn3VD1JPYvNTYrX
hs/KuL3wFjFZLytCLY1tfpui/iII868EprUGCRw/kTum2o5oZIPYuqRVwByvlG+F
gRjN3a8KIG4Ez+AGTjYVblC+Ilq9aFOM6nukjIoCMbQTIeqNevwTqDML+MNvqb33
Fc9VCSIXnaM9f0zSYhN5++1n6TL1QYxoWtQlkY44z3+U16b3WNcioBq+EK0ZVfP3
1yQ39nrY7DV2PegOlfiuu1cCxl+CHf+4LLNLoCdcZi2XqvgPGBI3npdtqqJsBJW5
VaW4a2CsHIPSsHAejPcdQ+4YcIKMObmFjLlw+6bK1wIJV9tRWOBnzKn6kZ3grL+1
JhKPs0dufoit9a6mzUVOwmSZXwAxnKCXZzHaAy4XhiB5OJw4pQoPTUM0AusNe0xv
+hs20z/xipxGZt9+7MdbhqDclNIjGy+H+F3wAkAjNOQLh0QwWynrYxbmMI18/N+G
50LIw26QfQhHsg5uh7QWwEfILlLgSXLe3ENE77+rZ+d83ERJ21hepsXH+bdAIYq8
yjuOQUE3gtVh2aJ2h6PHkK2+tkU7EdMwkxkFg9KLESA63ek+lCTabdjB5YdF0RRq
rPq8hAiTKf+Axmg/ZOsIyPMxYLsuEkhCsDUDutAUlwBWHEO6k58r8Faq7rf/kUDa
q+0ODvVn8bUi5Ef2Hm8gcSEEtPlq17c/ObuK6hncLdFlbnglCytswalfuBmU+EWW
TKu6NuXNJal3hMNPJa3swzJUIjK0QUu941s19FsejkJPI4V4X7voiOvevF/r8uyf
nUjA0LE/X8imdXCpkSRMJKBnI44B+bmv5WNdEv9fV8IfI4SaGF6dU03MPPJ3zUx+
hwbovgf5T4ibhCwGmJqP2Yg9vbJ51VcCq5UlRMjwJC7JNTmufTnnjUCO0/j7FWpB
CIMmj5xHgVaoqAcuRznYzeuF4/QWjUoAJ+gdOPQzZIxAtj0ghTHRGcvwh2lLDWv5
vIXUJyzKzE78IQMo/tU5/E7FiTayZC3wVdNiK4p4WGHrziON/XTU1bEr9lYf3bRF
jTq3lmLD1sJHRQGWJNfTkDR9Gp6F2/cznWhbYjSNsYozmH/0DWliZI7Pl8UTq479
Kn7deq1Z3Z5qip8zIftmBlZ5POfUzPUbXNoFe6kHLUkD6MmSi79s/yLn52psVGy0
LqMtTBkv/BxsMVoO+tYm9Ez+erALopcc7PBGS+ckPQlHzZCc7i3IOiFpfepJcBwx
Mnf0jsOpwwc2KNHehdIJJQ5ShpjX1HlvlVdJWmQMnc7pG0t06KGW6xCjVFTwLzWX
m/S5lyuZ6rTybfNikhAMM2unud9NWtFn9Vdjv8+Fhy1syeHuI78+ejFEzij6gOtJ
Gz3X3mcsLMlFIp6VyUIPNJQg/6/KhA42yVck1qaC1ScViJO3zEUAdD3VGKFt/83K
F21y0zdpJhNHaeqcUUL8I781qs+z3R1XcG/RFZryb2E4r5b6JD/fwM6EQslqcUDP
K9KdiPUSTxcnjBYzRLYNjKHhtqLwNFbi9GXVoTH/lilF7vqkn1fk8K2e1TRcibWQ
956uDWXHFUSAxI25tBRIrinQA5jVAOTl5pgDTxjtDzP7Xz+wW4/SWerwqAnUkTg7
VCDpjrFtp99/585krW8zJkKTHqGpdL0ZJMWqB+dAh+Eq9ABhS53J1eu5b5JIg3C9
DY0sEhkbvQyY9EtRYd395Wm3O26s/qksI3TmIdA96rgQU8oJxCh1girhZhNUE9Xj
zyPZL/zD0RCe4F84dO5CuoG4Y7FFZSFlLFn9MJ3q2q1C6pdEnyEeM9/+mqp29JFr
zv0VSjmw5bg4QHXwdoyHtSFYH6r0MtZkkDXrdiLe9Aey6qN+d7iLSCkQK3dpV/1q
lOxPzWRiXb1nMO9/t7aK9mhkyyv7OIT3N2kx/2BgfE9iksSprWktF2Fe/J+xbcTq
thKCUdsWy8bRBYRue4TF3XnYtWol2UBpF7ByMKLe9CTGWaTAB3uDF/uPVGBq1tD/
wYKo9a0XwpFJl0yB1Mt6iNjCZHQi03SththexJeddjrIflA5ocJp2u/jOidu5cN1
wFbY6h0TieEnHk1+EVOlPJGdbysQoSzTKJH1pI8ZM/XGN+INC4UEilqaxoEnFUlq
l4jshIKPvd5pRneJwhET6F0srP66/t3D8cj7H9bOCEjKFNeOk39n14A0E3nRkl2H
apjT4GVwsfdamOyD9H5VT5xvNkQvEgcwshmbmFGWgm8lN91sonW1U1Up2I01b1w3
apZI2YvDE0LjFaeCkzSdvDKKFN9ierq5ESakf6XAapdgejLP6oRHe0ro7XGxeIwt
fZXnQAlkx01PUmF0Id+y5zXcgF0m3CpapvnHGdU7i52V14ernCcb1eiX59j05xwy
m0ECf4wXUwIB1wb1lM0SeoBQKRNgL6p/p0hhrg62olraPlN50RWQnmogvJ+C06Ql
mRtsX5fm5/qkbQsI1MbrCZGiNiOkLxQOHG9xXcuVdsckYGBoxDo3g5BWAZdR9QKQ
ayzVAnaJFLxQmHsP9cC2REcfvf3oOB595B64jZouvUXQTGZzuChH4AFnQ6Qkvdmo
Wd5z/yiDptSJvwmIpL03CWYCa/yMFfZrOS8532WivtlGPAtkwWWyF9cZQ3K3VhWP
s7RI8OtNen/UYHieFBtx6d8gX2zKKa5hVyHiFCL0kaYrCZYiOme+8mKYP1cdO/wy
01QMwaJMrz90pOs4hAMvMDG5NT5m+B/ZVu00WAXfrdNfpsqGY/05lqm7gW/5vuCM
5Um/vr0Yv+0RpKOHloRESppLeeW8s56monjF0ZOphIX8/vmkzKCzBXw9h6aDusY2
DtNTSeMwt8JBhRo4cc6EDe5hI3rH5pnwICiMUyJCGtp3FY3zU3VrEY8tVyfDuUSG
CTZcrse/wUyMFhGrgozjbzJv96M4eLF8bYfI8SAkF7mbNlFPRrdGmc0Y6SXEq0EH
HZs4B1RTrGIPZqKcAsaFtro104hjLzJw5GV1CKWOkBzTPdiqxMNX8O43QfX5AWjx
2cAXr9exN5Y/mlHBdDPIy4s2SpKrHn3HgYFi7NZUDyTmdgOES4WDeJRWxgIM60Ef
JZlj8eDq13WyB6nIt/0QZd3ln/5k7qXycizP+RRujYL9fz8KV9KH3u4DgbToXKch
R329wUHXrnzdkn2FIYYKm0AiHk98gu0G9vDTBf8LCrBwysQJ+8hx25MGLzGM/3ry
deqeeNCBoY/V6iILnOQknN4yZ7I7oi6qMuCZtRUaknGW7LuEdItsRuLeizNMB1DZ
je5eURShLlpx4M+H2jNFDPzNd3YcOSq95Ir02pIRntf6L5Vye24Bw9mcbGq3QB6v
NdKU4JQzyFKokpyaBk9l88N1jKKFmvousFXp/O+klhxxhUZbGp/EcxhkaaPLwhGU
a8u0gCpAAKSU39z2T4BiRzL2ae0tXl+mZ4knLn/DWmJMqA3GtZXFqCyPaNPZszgO
7GAHEP3TVSJ3LB+BBky20ctRJjJlypP8TwJqlF05T/04EreUQDa/0xfwJrk9JSrB
DhbIB7IHTthTzT35rF0PU3mngaoTn2IHfeuIVhCc7FcXILt/q75TYcVZtK0/z0Dy
MOnDG7JA94ZmA3QocnW4umnMBzZa0FvQjIbDKBR4a+/9+5iFLykb3xvBRVCbaCwE
61kCTpmZhPKF+OCZimGJBcOjXaV3FG3w8oKMW/23kzraddtJsw6GaMIqnrrGhY0H
ZQXox9UKCA2EPNtCarH3l+Jm8pqRIocMTfpDa6ZO3GvQLQIa23apHEIqxABBHKE1
cNbkaoQBZiFCy0FdpeCtFOfE/WNQOVDwEymxTLOhHEiSecz534Oq56RFPsNU/hfr
SRRvF7U/cJsnj0u36HQFGtHogjI/Y4FU/N+dS9tI2r+ifk3BBTvl2aJHnWDhwvrv
a9KhvFyzYgDkIF3yZeSun2Mi+mEldMnyxk6ziwM18nUw2gcZCUQPcKhnzmcfYwkE
myjHRavAx//jp4X3mHcGYX40hGCj2Q3jq+LCwmG++v35ZMGD4rdhuAj9YEhSfT2X
94asziwyIhXlc55LMP9XuKeycrz3bqerev+SeGC3qaklRFGNVwUSeVgdb+H8QQQ4
Ggruq+dGW+ZjFSwQvQSHNCOXLMQ5m9bgYA3Jmp8MX1sWS3fFqU+Ev2sO0HGeNxzQ
GlfBiECwSskjv9kb//zny3n+VxTLbVNiITBJUY1GbCBSseN247Ljh9OqSJ8Sa1cB
MQ5HaGnuWuJsikcOKdc9781THXE2hK7pDEuyu1tuJCYuzAKNZsMBjVOxQT/rRFRB
R1GrTKq3K3/aWapKSO/6JjnPKC8TNsbS58gZMfUZX9OxMItcHBmPnATfDm/KimpR
Z/3g0powDZZZRb9ppxMKNjtur6qEKTrzKxQpkkxJi0ljyUD1xvE3ex1by6km7guO
WHG9uZ74VlHrCIyo85gfdtYmOLod4YaBM5bUnAzlnVylVGJ+SHD7xNLwyBUK7HqK
/lvJzruvCsKX7fsMETTYyFgylKF/dQs5QJcq75NY22muS/MqGa/MM8zUHHA/P8xN
X8UG/JT8A0GGcsQB9PSZFCLvJmXRndeugKYN8yTDBOhuVt0T8XFDNoGkuXJGNCpB
9uz1FGl4uiu0J0NP5GZsVLJwmwPsUHrxEpAyntEFSu9DzEENSb2k2Dq7ic3YcCcf
6I6eSTYrCcyDuQqzK1OLqXmqlGZw/sfSOXuIhpd7Vgb+UBVSX2TfU9eh+oocow/E
Xiem/GJSIcI0XnbzIJxrsga9+Ra3+TAtemVDdiaEo6yE5+Ogd3zPDnNzxxeTyGpy
ZfL6Fi2804e2ZuY4RP2Rfhtf21+6ko3b1dQDHHZSyScg1vb0JKwVYmyCDQw0qGUm
BgMKUUYa/LlCEc2ZYk4nKHkxKB2lsXgKXQaCJuS8wrlAe0wI0g+NDiYn7PSFx6ca
kiANqWT8kTbJXcmQ0jNQWvyBdDZtMktcNTHPqFQnSG91jNWNacYQGYtXsHn6cKT0
/JC7UCmCXIaeiRE9JPPo2by3feLZt+Rbb6cNpI0Rcv/b9s1E30R2P7ow8UZJjkPy
4L5/ivyczGLW28UbkwAF3Vq9ZPrUAymfXg8T4eET5yVskZJY/cG/cqL7hGb/Vn0v
uwsJDy4BOnMc16hMv6X/XoThDlE0rAMxvSNafVAVkBaix0s0uzKrPH5pUVA3G/5S
vFoWs+CicwMiCrDoZgs3eiiTSFKL3hTdwH9LGYBH4CBKgYxfLZk+pOz/uk4E4TDD
gXB9efCQeYRncPwsU4vuOzh9SMtUz44e7Rvy7SZW9WHc2PYJtIpMNKcky5N7xLKq
Kvey9rvp6ssBP82NU7CbJGCPytHD0kxyxhzEu7ZPo6aU1hCZKvt8pz0dQWUim/ck
2+damEcDUPJWzL67AVeMN5SPGuypv4JMOfsQ70uTA7194GrAk2f6tz30CkYpeKf7
iycGJmm5MLO5kvMdTIIVB/4yzvVUbDjRQbGi83Nr1SsGYaaR8ByFzJACOigWFDl6
17AigpH1ahTAp3Huc0ctjk+aM+oEYUE+FNbG7W2TZaIXy8xaW+kK0UaiBmmcXB56
6Qcfd5nT7MefboXHhxfU1WtVmiWNuw2rTVjMkwXUUXQCepqhV/mGaX3fHXN+uePb
tLVkIdyFWUy7IEpHMCU9mnx9lxw0jQiGJScB0YuFHp3am7wyZfMk5yJkOBcTBim4
bZT0jLKkTQKdtzbw15AM6Du3RHTDD9BxTQpJv/lh7cVJTJ9aa/mugkgApP8yqEPZ
z5rtf2kTS1ke2vm9vlVJGAQ4Wo4QmmunbJucIZy8/4cPxLc9+j+KwbQVINkbAXgY
1OaxvGwxJEhqENXpK/RWI1q0PEFa2vBqRuza+svhQDO6/Z19QQQm7+Qs3gNlyjW3
zm1MXQrwrbFmJEHps6ODDohDBEj2vqc2RhCIMbGFTKBCyXcB0MNMZZFR8wSFnaqA
C6TerJpTb7D0NSJVKIdCb0/DNzwh8kzV7022CZ0FqJjS1ulw8Gt7vC6qeb+Yvkhf
TbQXZu3kyHNfjmVqURzf/Ur0JxD6Syk1oEFHEFBozdoMew8j4BmwB+LykeUGgh9E
9pCwYFqMl+Hr+YaFenRUnUUly0bIwu+yKuSO4POncpSLAqRGh1CxjC7C8unekL+5
Ej4l4h4xqMxDbSHH1OSpfp/kXeqK3kaM5KS4L6TReoRgILzLh/G3ohcp9ewApzH5
iiMxI8MebfDHFfEUE5Kv6kpp3K5OaYyR8duvFovJKmcxS/X61+C0sl5ZBCdT4pkz
brVZ7EbOjjZrwylRCi1SoHAKUprThvX9y7qFr6Bwwz3YZKEf/RNyKFtVQTXMxhMn
QFx58QLI+GJt+eH/zBmPipsWG20RKqiTCOJI6g+CcUowfFWCB8zarSg4xlmNadvv
j44VNtwnPJ9k/PZXNSZeaWoPL5EG8NRGBsdpkgZuJYKsRGS6N4Hbywnhc4oby8ek
XMk4SvULHiR7LPuVGOILMXJMkh/raRhcAYJS2eHSLD6eV+JuktuYNi3Ys/cwlZkc
gvVUQIRNe9SOS8PgsdBPR4ImeD8XL0b+CcM52uyMbZyu2oaQCRpbxWOG9w8B09Y8
jjN+SdYQuzqpPz04M0+UwscN0CI0XUh6uHUzYmLU/ZA1DZNwccLxZ8TcAu6CxMfe
Bjh9Zc/NfrPsa3QxL0kwgsN6jjCbBbCoMBoJbLzXWJpGHtX2VK7kXNW+Rga5OwEZ
VwhqmKU4cC8RoOwplt3U/nOPknI1bRjxYqljYiw0/+LglYIwbwo5MK808WZLBctk
lngSXydsTlDN7zvBTZD+Uqav/jRMFO1iCDvBxNZuHXTrdBWokPnEnFHMJM2+OME2
Jaz5lACKN693wPSyawbw86lOPa3c0IzYemfflxPddtZ7ryGXjbLyvLIsdw1/U1NY
lbnurqOo9+FZczgxyVyksaD+rsf1lGkMmLqTcGu8tpRMKbLFENe9wUTtc5zvBEl3
1OD976LSGifrG9OR9fOIxNUoLucTek6U6Ptd6ubQX7YQNGqKhbPpo1maUIknh/gb
dP0p5LPg5OllEafpEMR6Y+D7yE3i8fbgC/ckTWoLmQv53eM78VUppKW8IDO1lI+v
S2K+PWgZZ2MQl3WTw3szAwQN3T4rpk5ReQWs2FZ8vEdp7SYzBjUY04GETMuBaypq
IFJOYtFu9hxy4u6kppXcNQuTsuwFNHvOfS9QBQX8OuNzp5teyCRXtC76NeCNhgqa
OyID2V0ag7IU90j2lxBYQwPdbc0EGfaSkCxabMzSZN+TTrbi3V3LEnuSB+apuzwg
A8pYd5XlC74iRfyuT6fODu2AD0ptQavycUA6QtA969A8mONnQjCEe83Cqz49Uh1X
Z9pO8ewgLnU/kXvh0MvpXIamTblO42VDFfH1tOlZ/QsmUw3vw0CfMn/z3GCEfsoU
3Va/mqUz0LUFYMh2zmhpgL1WoqbgCRZLOMBPcayKBDRg4EsvPrrsSIa0E0hgzkzh
LPb6HriIydIsSB+xDDj8M2UnpxJAQSZjBjiqeblBP7CIHJjt8fPoMB1MDU9W2Kus
2RT0GNi9NhJ93aPgEMhMeI/rwhDGFquwD3XlHTufdExOqYFKXgTtBDItk/P2QvdN
1POzPIlmOYiYCuS62KkLetFo8q0CJlkoxdluOOaZAHv3RzBhaaWDaT3nkDRbT+og
uTFDex10zE6juGWVEXlWi8W6pehyqN9VGsc5edpPmdLFqkWshjkO+PtAsifY3GWy
s4ZADslmInoVedBbuCHv0jHa0P4tV0HrPZZTe+RrMH2CSkGmGcATlYfIsuVpHjBN
r0Ii5P6nmzZlJlHx9cDAsvyvndlsc8kD9/nWdgGCU/Z6bzDBTmwBlunQfPKj/i1Y
bBMzph2G0ZabX4mS4y6BS+5xmG1ygkgqE4BOSvjiAgCt7RKv6JLD6HUhv6ItiHBH
H1QCe0NwAC+lT54RDBi5Y39mgTCRECsUNLY86PsYLo1CfNwNwjWVeYQ34HRQCKja
6WxR9TOUgNsrzaSoOP2LASc3RzQ41hS2YKIhC7AEjSmj6bZ8u8LH7tD2BVR2M8lP
hoYaou8FdnGJwGIhl9J7mfBn8obkGHVtGtYbsjiq/NK7yApoT9qNwnnRxDdlRuwx
clVpdUNkKFJo9DHZKi2In7tOipWCwQwhHxJXSRjtVFPIToqMxgjm4zulPOvqaSJB
NYRdDFzJFlEPHll501/2ltsBZcot5rvX8sDjqmjEIYUIlxaCGKQuX7RK22WhI3yu
V0iNko/8tBorqv6dLtGe2lq0Znr14Hlpm7W7vrXCp/Pcu+O3pmdSr4+wmqdgihKa
qqfFTn/l7MUZIQ8CN1wAm/bbze4xVTtFB1rkHg4DDeSilFkKTpFut9it+oG7p1Gg
qlqc3yL24tOBdD1ykxO8/p3Yfod947GVWQ4DQmU3/7tXUJtm1tVzYJ+62zp2yoNk
wFhXA1O4UIdtDq6eztPIixnFHfzuXde+LGJXhAYh3v+w73CvfCPHdzXmNyQ9vO4G
i6RRmNeW5TUAYAbbHa5R+BsK+ytsLxREb1ZpDKk9HxJvyiSN6Bqe7Emw9+E8yGAX
xoW9R6NAj8Rkgwa8LxBq7ag78paDX/O4eSf3dt0aaYyserBI1ReL1+TTMK61Gjk4
+5y4wPJAH0I83XvlObUKz92Ql84oX/WBiQ8C9tK1U7EFVWGdDGrJmCeT/N4pwFUh
YuF6v5AL1u278DY8Y2BXzNN9loBH0MyF2mtLPt5ArdxT80NXsDDZVJIyuJF30yvW
5GLw87BJryVmESps+WLFEnWTK/XLljlMAwpUmR0OOvZZulhbvz+f2jDkRlRr5Y4n
n6Cvj7q34ihIjDhdVXLWEx1F8K8tZL1P7KlXeFaUKMlzsaK1SyLVwwr2I2047VUy
iG+CrD6uTn6UzSqZmHbpQhdcYp1ZtXmkLB8CwPG5NQzaHgFbyo9v14/svm/lvdq0
sFAm5FqC+zroiHDVbRP2K1Xi10U/dSOQK5glqXlz52lOP7v9vzq9Qisht4jwOkxz
PvcuEGM0TH+Yi/Iaubq6fQ1Am2wHxws4zVSt3HPYDEuEsuTgya+oe9q+qG6pjO58
Wcu5cc/mzEOeZEKr9gOANHl6m5eHbf2fQWX74TctdeTEZa/iOmG1clRQlG0Ra8gC
ZLUczz3uu9Q6MzQvNZdVcd5Q2WYMNYhE5Qd/TsaNVvTO6F7swqF7sDvBQbu2ZmmG
ga06mUjk/tWedsYWPOs4+BOMKIoc6E1IFiGS+6lA5RLWEZEnk4Rjc2uzrf8Wbsfh
UmcPRqVLoJeBJUS86geHLSHNeYdXO4W8aef2ShcIpofPqrvk08vKTYwbpEOD2Y6q
7y+Trqtfb9VxcyX6nmiQbXFzuTmMi1R9VMHKbHDeXGt9jg1Gw3B4TGmbF4oBFahs
wrkOJdj5Vn9z24S2TghF/qClgKam0m+TdEs3cAHCbVOKeTFmiS+gnmo++lL2lfOF
IL5AZqmUQX4uiFgNaj570cBc604JN0QQAk1s0EYUpUK3v0P5s7z0JOS9WYNKRevc
SqoOJWzt/cEmKYjpYhpT57YIMmwabqbQPqyzNea/585lNARCsohgJihYU86MFcnk
qK0nU49GhXXEVgvbAS4y//dgfMidZlqOHeRdpJGMZs12on8JZHp5lPiIxtDZYuDO
ayDG4+Jg4Vvx9QF9Fi06CmZGe2d67WOutsjajfX7dGZzxWl343hjbDWNAgnPp8fd
ZVvcw/IRgOr83w+kKIsSlQSG/pAJggpfGI9hTy9Jr9c02BTV4jmPq2iMvnuNnRS5
wbWW3R/CB+psxC6JfnxDzir/WemrLHyndYs0PErvq5u5l5lAwY1mOaufD5Fbjo7b
jDk+A7JZfQBioIERYsTj+Tt/C7wl5CCMS6niam2HiMiPgQEMrw0O0Ym+82gieAcA
wMsRkm42S2MeQIG2gGwMHBjoANGd7kiB/e4Mj1xkA+iEQznXoYAShEsabIN5+KVU
0bVTVwI6mFD0yehNu3mMbNKKNMQl+kxXNa8IOC9JODGs4U9XovdSichwfNZSPNGI
HnPAQXjTHGIiyQ5RQS9lwm8tKcA8xTfWCt0Y9ef78FR/9b4dZZxQ81QqC1jSrDrL
lJx+9tW1mogZg+9ltOnAFt3QaH2dhAGxXPBjAUXLAGKvNBQ/u+GUrvOxuC4j9so3
M7Xf5F4u9ovmxXCPGOz4IGsysc/Q17be4RWofgTQ+aYBD/rzfFkL9teJWrAVC7wN
aIGr2PZPNwgsvRQkHAufvQy5Xle48jMv5cVePy0Q/F1qJ134eZkCY24YPAKL90aw
AlfRxSND9IM+s+CZgdq1gXQIKxW4sdBAp63s7VYu2AIh+gr0aAjyWGemu/jHiPCN
yAKHKTzgeKdTSeIlmEHiELmtILZsEdD2IiNPiePETIuFWsAvxBY0KBS7xhqbLpkx
XHTkAYSAMg5Bidt8aJEkBAH8S63dYUiQS7NXGAZJ+eqA9HeeFBAUJBVyalBix6RQ
Zywi9Jn27N+K4CzBC1I1Lm6tBMvdVVVz+NoHXFOocEWhbytTuhfv0IbM4QHqe5Zj
SAb79p9njJAB3D6qeeUpD4+ZaBjXHoyDAdVojM3Dx/9pX1l412nKIQah1tWA8RzV
dl62ILJctvyI/fS+FFqtj6QsiK6/wZOwABRE6Q42o4HJPsuFjr3uvdqxU+SmpPnw
tVMIy+9j8C4Et035I699ISiXD7drvK0HFg8aq3gJDyD1zKD7x/UFkd5a7q1vbQ8S
jsW6toRXgJEeOHUCfuKILj5PMDpGnLyF9xaFxjGx3PXIeiRHa2xu1apyOa46CqXu
tRsgrzrsFPMspz5mcqnBa1DjFB3YkER4Qgjjc07W6tCYj6E6nnAHTpgzJJlONs4y
bQheDlsuTrqkh7NcjDTZFDuKxveST02zFgtkCXUw0FPsm9ytbdYA19GdgxoLLulr
823w9HltkXq1S8na+I1fVuc7Kvru3j0bbMurrnnX23nzRrB85K8BGNkDT2J47YnE
uJ8UgF3U5fvoLahXOjXSZpc7m+0ou/3eJwRpBlkm5TcGSG/1cNYeYuLqTl8Kvr4Y
y83Rh24uUXAZShgClfM3RwL16wn9YARO2mqwaZhcK1TsGusEpxdevB3y7/aFy/wC
bzTf4CyKZtfCEOsEX32UM+6PTMnB5ftjUZThLdUBiXigyPdyge3OaKLR5WgMBVnk
XQHZCGqxY0KyX18qaIFF2zKbO/8/FVf5RaKDHGBIgUYPH9QJ4Gj2m0ap81+0u1Be
aiuREmgVJFRIUH4AU8EzsdOHTU8lBdn9rxOuRdv7ztyWkw3l22//lFlr6uqGAn0P
MX33+qHunHL1IKSY8mNk1+9piZtQrc5sWrw0sVn/yzZdQ4dx8MLSrZ+IURikiSXC
F+vrm6f/Rrt5LRTa/JvxMdbDPO518l9HP68qrJCH+uf73S4WmMzr5QhRnarkKEzl
P9poqdcmt+0iT30U/53X9b6gzD/uym9DLyzQ3OvCO2VUQZtdfq245hl/d9L41+kE
skDwK4lZiQUR962wyGr+YUPUMCHvN/ZxLCpCfURGawzYi1ilS4HksY2mNj3+rP44
RFg+2QEY5giuCAUxwi5M0IYHz59q8ciwK365NnswXi2lwRG5i+j9pWhmWak1rVo7
GDvR/JRr64sqPupY6byDDlUY/M4Xz+IBnXXgWAqxnTrR7/UpHPCbDYJdH/sGcnaf
+gGy7h7Xx0vJJ29xbnPAV+wRmgIeS+svSwiY1IvdWnmh347m10EwnN9g8Or0wU5H
yaCSsi1ZIrcLfg5+iBObnH6j/lk2P/Nd/rNswBI7qwuW7qMrGRQgHh6hUHvzktCQ
g84PR4NF90Uxhq2tzpyNGxmbPB1GksRkKvVVNsYOpeYQ/hgT1nO15ybNEquJFk6f
Ghz9EeHnWNJkhcRnO3HeIsJiaN8bawQQ5h0K41EqDHODl2JxG+vfxpS8JkGpMyTN
4Xc1PXOFTRHDu1l6KhjM+Fmf+UoEWg6A6oPxUcWn4yBho122coMxAaCjhe+pE47r
9Jv9MwP+mVUiNds6ny1l1cGiprYhCpzL7LSRVU3Nc7x9dCqHqIKQXrqcTVc3HkKR
iEOrzJFd7iq9n2AACpkUbEKYtedLDm82lR/T4uczpM3gi579977/1cenv90fprp4
r2BK8LDWwefr1hlrebtz7t0jCWX6WsgswFmran4oeUakUW3gqyXMzuXCd07vGY7D
uvljNAqbrogyuXtfL4WNLkPrQ54JR9G+yUJp1TGXW2cGRpEZYiFzUVQ+ijdV9GZJ
DNStCCRcAq5fYaa9LJYEgO1GJIoxy0YcSYajXx7brJV+5dmCxp+1m0IACU3mnlEF
K57lEjREcyrOUm+Z1KAF7uTpJDFliVrM+qkZHlEhGiysTO8gqF3r/x5bKK95LITX
l/o25oYm0c28zG8OZLLjCHCQtBix+qskLgPvABObAtH+2tB88YleOMFkBwiv5Xvh
YLbDAEapCvAGo4hnZsLQDKIVAzO+sltGbEWnjXxfZp5UsaIdZ3i+uHU07vDt+e8q
7fDyzUrA7LuwsXdX2DF4Dgc1Vpr9DHYyVRYeGwDkBrGIcAZiNYOD3ODGRS9tUYXd
gfcNUKGU/+Sz1lZiLBOztiouENMQ5/7CBAfvN3oGDIE0K2Ypukq5fSt28LDNirYI
/ioAVZysMm2HJHMcj3qrZempOWmWIHKpcKkrFI8cDXCqPuVBZP4myR4+qDhxwAPV
o+NkoqaeUOqMeFEjFrf1Ry76TDX0G+UwYX6rJ3Idwyp97lELu4zEs+8UNbSftM8b
xZf3YScyx52B3PQm6MDtZygOw146M3cQS3OZ3gDvJOwuI6AeW0++CjPG5xOX/4fd
mk/I7uilBFVKKkgfk2dsKAME7PEr2rIgG7gPoEfuvdnpK8ks6NL7WWT2Jl04SOEd
pglbSgQ/SwtQVT9cC2ny6nI/U2DJ4jD0w4fcVUxaHyc5bCtZykTtCDrLPkvchGKQ
SSAwmYQy+9i6cEDljfAn9GVaZ3W9ySuVRcbelF7vKD/R/K+CkJ38vma6hPLIx6uy
rBmylfUyw8gBMrjDwwN/i6KUYcc+Z+owCJnB2+0KEkHcraR82ag5WiuAhb7Qk3we
CHUQ53UMgrmsPVhKXBjsOVBBmspZejh1NRV9pWUSAIyYPOs61HpDb23gEaYkeLzw
Vd2m4BOdct2xh977sjeuVjPHl2M+NBqJCZ9xPeZALuhDC6I69bnVYOYQ399B91Ha
GduHvykB5u93DXZ3JApTf5CiWsje2uK2MMxZwfSaLqnfR6kUWi28Bo8GfXnHBIVK
73X5BtyNy+bKOFPHp+6prT1/FB0bsysoOerlAyh8z+ZenTe+sA2kXS4eck1XP4SF
C8Hj+TIdG+jLMCEmF1OHNFri8kRhIOBKHg/O2TfdGc1pVk6r297Mj4tLmM/2f2v2
hWed1bu0vtzFRMtFkjiKHxC5iIntwf0Fdgfgi9wa/B6bFD4HKwAc0zVorcZ5zFeB
CL26Qhr3xRuKbPTUBkDfvbbjMLRmoBosfwn3t8hdopqWf4Yw4UWbzwRMq939oFyD
Qft8IIkafcpZzlWM35Brg6vD82MMgxtrSc3yAuHfZH1QYnIlaIw/6kGSXoWeYaKZ
8ozHaWkev+7xmuYP+7Oc27EeDKSI2OhijwVALu6OUH1ypKHAMfKvTsCoYPlL0eMl
6C44yHvDPfVWALPqmwA00zZV2XovdfU4jOHJq34PtTxE0b91OMvqjjCi6goz1h0g
66dhLMPSIItRcFDso4+3vhuOZqFHbLLbSgDRS3ig2vxDP3L2RdfMV5HR5XpJnJkx
jq1ca4+IHEC5B014mn53EJkMoXzp0iofA4kxyNWWKilexPhsxlhO/O4gcBp71kyz
t7RjGncWcMmTZcgdQZZngHhlmqd9V2p3+NsryGJ7ziJNtKMgrn6lsNUXRzjCQHlh
uPZIgNVpd6YHZmpdZYB9g+EbQNAVF3z1xkC2HCAWPuIJanrXeznZoI7YkBtMuH4T
4FcanGqfSEaroP0xYCCqLG08/QZgh2dX+jrEdvV4ZUAWCBmBN/mjId4WDiDsTLfh
kzOBXDERc+hAArfVFX5TvaNlHdFCRYZ5WEBTtlLWc3xnXAMqJGf1kw7lHyKCCUCu
PFcU6P6hdZPhwUd9iPa7T5mfDfAFRqQWCjpnvZjA1KaB7tC9DXMD031qIRdVZwO/
IXiGYi6YRpxiwASzugfAK/PNCLaHRyKcUYS9+L6aCx+0uZU5PX2Z/Mm4RYNPNfQL
PBwbpj8KZ14f5pnSWnN+PE8rjh+KNjXEaNoD93XOVK92F6gfq/Q/y2E899YFNvVx
KjSQbr/3+J7wLgM0n460xXeNmQsSSzyvlsCGTDOoskHvI45/RJ/PBCqconANgeL9
eyPPrt9QWOpjsU4EJR1+H5p6aMFmm+oWxXQfoFge3JRFfJAuE3IlND0rHTS5PDVZ
ts4hBAZAJl521T6YHZj6uya5NxSW5NkIwe15Sm+nEv4hN5FQ0KRUj/zrWZ6M+5aS
sDxhaXFIja7o3ML91cvf9VVFcf5Ej4obF9RxNIB4REDUHb1AVhWqk9yqbC3+tMDf
u+wMml6jwUlUMvBwLdLt0KazpVOUnWW3Epj/NO8yRGTfCHcPLb182WOl7/cAQo/O
uWwImIAuBzSc4h7ohuXyxTCosE0DBmTfo1ByqrdJX2d9qNQMIvfA+Zfy9+g8kxMp
E64CwWvS9n9Ip2mrgJ/s2ozrrSgTWzNoHXMTFQyn5Ze0LbtUeh0K5f9w0SFRNZDM
FMSWZXXUApg7ZQVP/g7O85vdsfXxf/bzldppI8NoOf1NMGQBiDo0Vut5T/xd1c8/
uBuLJP8uqiY/B5t7zw5pGJ+KAwlRrDWpTTe+WD3AaurcSAhb8MnsSf/25E0o9BZF
nBVkg9JWEY2O/AwZlKXO7XCRJgoVka4UbIl4mNpnHtwg2csGlea0b9m2Y89GA058
Yfc7vhxbqE8+oINR6N9wjTLr0iU0iOhOaY4d51s9N0cCR/b1v+3Hjh2n9QsqWVBe
/AXRGqmcmrFSczX10jB3MDDstx2r79RiLM+A2fDc2SxQik/dqvvat38qzA7KH4Ze
KJfc9WOQyQ6S7CCPXj4zr4VEza/SsuCkDqBViZcjYAqkrXTc/pMzbO8hgA2fqoPB
vLS1lIXv+MgS8F381Mw6gkVcHPCbk8SjSUSUab+OLWkRgwo0TOnz45abSMl5whs6
uiaHcFPY6zjIg55qNsY4Y3WHPQdhFpBS9FH9PQmzHnmy48KtJ/GJ3/vAeetd9aWa
NKbtrnVpYOdIHDFOsX3yCDSSNjK3hY51yHvvf8fPaiAEHmQjlHzgUCFef52FQCmo
uxKfvFEnuMo6tP/IoBSfnF1eC0P9uKB+21WvTl10HeZNtOiiDiHBcXnaTxm1PnhR
9W/tat7f1H3y+Gp2QvjY7cL2TcDwVUv9zf7aOh1tQfQjXeDuaoU5eH6uIoBW5h+r
oMQuP8pS4tC10dmDD8sSxoT4jFj5ONpo8slRE3VGFcWWx+28IW/Opd7S8Sq60B3g
dUNTk7hft9u8AWgMpCW/gW6aSZzg5N56GtFYMh1G8xuNipBV/ewQdgxmrx1a4Hg0
zB7pIFgb0WerJQF81ErQB4GgNTgvKhcLsBYQsfXJ6MQcdSHnXw18SDpBtDswx/L3
rcBKSQMwuRXqjUpVr/MTQ+ljOl9plmhWikgbKPOHSelA2bEFq3Fc6FSXNjqxab9F
LYiFr0e4SG1znMkV5B28fM1aMl+b1ETv7AXSFW78JZS54SCkPVhlcrxhTNnPGKGu
Lpk6WHq22IkYia30OQJIPvp8t3gvI1V8PQ/DI36PXBzGZucCFkmx5mB+au0gEJ2m
5TpD44D8cjKtxzjMuEkKBsAWI9V/2XKqDs3TKSEZSigNuXcrICnvVA858JxP3rkY
NsNmFxp3Eelw+mZ5fB6nb0rWddS8HiN1yvPqYdlUfsu8EnavTF2IWmpO6VFDA9iN
49V8l0DKL7ZS6BBj4XevDLHkkw3C+0LJ3TFzXbzC0kT6fQHyb7ZaryslPTHNPtIo
r5XKdbCjF+gYXCsBsNrb1hC3zH2ZGXC9oG9YHaOnlQM2abML7qXZRtHS+Q/ncTsy
RmmyT0vbxG28uEFtQ93C5+dyqaag+4Wg72aV4lM9SMoqXcdGeEN9hztEeD9fS8e/
/mWrNlL02h4U2VnHCZSQoZEOW3b0F6TGJJJUaTCfJAG6o9OEVLFRQlaiXgcMaY01
Zc9QJLM8D1akDz6+au6rvsgZgLaf47NZvK34x6dVyMXmahr2lqVJSmg8pqSupQRq
JSBSHyPX4SfD3aXQif2ELK67Qr3y55JzO29idZzyvUEa+G2+aeeG5Y7ZLPfBBC6J
EW/U8NwvdaD+M7TEoe6cokb7O+NOqoO2DZYiiOYI675wVpTYof8WdQax22FzWP8s
zhVhlR3A3QVW9B4vgkwM1rsgogsARn3yiev5HAM7TB+HGSntN8t6fMIKjJJxXc7a
BPx1O/pUMqhIX2FVsg+HgP4uR+qfP00jY+dRogM8UQX2qOawBiA0J3or1T2W3/vJ
KRtOz3JSPuLLv5nXG5WuNzfRlNzpYlvl31BeTd8tmfmz/9lCkpykCNx69/W7rmJb
9i982e1xtCq8UNy8mtd9MP6T+q3P3vQLEMdntBdNDE5Sb3P6VvXkSZKJJTBnkgnx
UnyuIJ2fyq/p/o79nzm03uF27jjolDJufAmh1oepvjdx6VP75GDUunIJf1bDU+dG
+UXk83SVJLy9LDqdP1a9WuVzCaPSHGwW5VqasLcM+MPYiUA6aOKsZoPDW+Nr0O0y
x+OxlgBQIS876ptWZA9scr/TbcfswI7q19v3RsB3wyaPPmdWvmRkq1e9R2OIKuRr
ArglOyTGy0sL7U5M3ByjjfOsyGILcQ9KCpKS4tDcN6OZXj3Tt0RiFlH5avhRiJIE
qcZxqe0yxRMnmbiENNATS+WmYrUM8F5qji1GZVRZJwmAam2cucirnzxdkSXe7D7l
60yaUetEu8hLt1FZNdQRTh7vb20//sNmsFI1BZoI2E4yZlOxGAg0N2q+Hg1JZldZ
pJC+7fv3hbeIGP8IzuaktZsv6Bae3evV1+ROxj2p8wJ6RVi/2xmr42w5GxxU/QwV
TgAC4gYCN4wUZNy6oZQsPY8id4LoayKKGvp6qHIMtpjDeP9WTlBXWmFutJv5bB5p
vJ21Cto4yXeaDuGEA1A97r1sd4XJnwzDQ/dh2rv4an/X/Cb9+ieAbJ3P5DixjPVS
QRK66kLRt3GNFeeYbQ961nkmv95kKltihHFMrJWkmFXKavv8/NUwwt/rJtq+LkVf
8z+jc7lcxqANG+WrX2HrtZemnvkxAygf7/f+G2ODW4ugVuo1NdO/ynQV/GQqvJi+
2aaXv/aXmgGIfE6NwfdeLVxyl7kfn19OI74+vMA/rtzYR/eFzqMi9fdAlHWOSzC9
bqrp1wzzPqLQEwmpX+yxfYcCDbCCMedc3I1VOUauPjxghQl0wuDPShCf2Po8rGqM
nlu89Xmko7vTB9meh9pZ+ZUVipTPAN4EqgF1xlW73v+Y3nIQyCStyUgh+g0BSgf2
vfKSvawiWJxrFdwL1BEc1yo5V1A+TIdvYX6GrRTjMsK0Y2Q5kviLQ2xD4NMfoqaB
L5519hWwb0juzQ8+pO0A3nlyLu8DGWiE1U0noXHoTv3Jtxs8rDKlLEqu7x1SUxfc
H5QIdFwCS7uAIDR18PerNK+cj63l4IqM5X3TQj7cOuwTKOFS6lqIrl3yCgS8R7im
Y/szQo/Ao6gx1+7h6MHiqqlHMsi7CojY50+MVvDeT3zQkNzvyuGs8xMWIfsWjrKi
zlOW84HGx174Z5vlRWHYqrETVjOkS5SkYUjF0P++nnMDnc2If8GiJdeoL7OI4Byd
Xw+oZarC6JaGaKMRfxVH+/hd2gL34NBqfcSRMhz09SRnNwrWl06D9J9SJIcXOJHq
PgShfMWRCiKzbgABgkW3N4FfQsMV63ZRR2Q/BfFEYnPq04oxRZgOEeQluqYH6g2J
iCvDGQYYCPuk/K3R4bCobUBXoCIOPgA2Gi2lOfo/hwg+8VELAl2dnphnm2iVQQEj
1/sEMHwcqHsQJJ4OpJQiHt2B1xDagezJbDmHEAWkKAqn1vRGHsKmGSn3Tbam+CFS
ypg50jvsKBSzYgqTzryZUjRn5JqSTzFATiOz1pwAPtObnQOaNBdVZzE5nsXgko0z
QrhTKhvPJRpjelw8iiH2ik1/Y2f/RaNd66GEsGbC6nwe2IgPSucsInEjypo/h0Ix
fUbNYyfc1TQKVKcc3jrbVrp4oQqgODhfNKzMkSjtmAiUota8ZBnN7fKDWsoUSf6w
z/CHTkg9MM+eUX/08SJ8HLcTT3Nr2kKDm22wNUZsLP9st2ACdtnn6IS/bb63Wxua
VtmuJ/WFEdg9FswYGGBm6ug32uYQN1LA6FTK0d7fKkcovS0mYuTwWWjKFTn+xjtC
Nd4/xKViLdXJ0EuH4vdwQZL/7QzSbAFjxdn3jvRKkyb2oHXrdnQO5qoI4DQq1ANM
MyyBBEOf0V/JfLhjAvVSi3d3pENB3rmpdqxiI20FspSZB/bMALFXFfyJ7yTE1hoX
F9U/I27wjZcu940GRGBH/UujsX5B5Me7L/5MYTEI7UQOv9jAWpEHMAfgDpoY8QBM
EAK5KFVxTbI3BOXjspu13z/v/2OCdUPvO8k7e463TLWvkTHWgtnkmSiNkuX2M5Po
VIoBqLr85kYOj2c3YPBC0GmePbdiuUsTaZGaMrklY3zTtE68ZcKOQyMMM6sz+WsS
OTahtZWuH3fP/e+bEVnpT5u+gdsnkJx5KGNNnw0DT792IH+oHBZmEIOM9lUzgi52
NiSF4wztn/5PZVuFXdFcK9Nt8u5dIbiwS4lBmyujq8pdKMEW6QltL1e20Ng0VehU
psVGkSLZxu48/3+66noTX5+IEvEm1TfXORjniTpXMxczgWDJlTEts5rt3l2RtR8Z
Koenps72RCyPb85s4vMto6lbutc0gbhBnF6tCrlL3lhZBQkFMI2W+TltOMXQ+5mk
AHFYGAAROLRtAl+bAjubQwgP7TQSAwsiDs1shivGJ42cdqJsKiQ091MsHEtw3BF2
8Tbgbw3gXOaClmJXLR1ZroGof7YaHm88HFvgLcdY7buFbfUwwbOitUTRmKm0a1x9
vQHKupcAjtz3b9E0JD/cpZrnY3sBw7tygci8sL42j1g44ASMXApDMe2vtgXRoH+W
lxzRyRxedTTIJpIFfjWwRSCSP5940u2qvRxnYcGZGUD7blKLpFSpNY1LD0yYQdys
EXvuvamQzS1Um2k9oujK1QLwS31a8IVoGMTnh02HoEVse39XCoFLdSz4nu/jiOiO
IO67iZE/vGGW6kyGv1hBbFwTUvSqhWjTOwoNPv9/ztajcv9h5ZMGJSF3elQGNrf2
t0vgsDSKemMMd9RZvxTdAXC85D3k4tvEggWBg507sZhyaFdqecHtF6BYBO4euTfS
gJGxzRJ6Fua3HP4URXqQiTUIMy8n3BFknb0mhD/4AM31zW6ILDeKZi+R85k2fcYI
tWZ8/9eynGU8iwZmLQa6Iuxh3vBUvkPuxqrJw01Aub/wqtVzYrY5jTlC55f6+pZU
Dk1yvr31H2pluw9MMfC4XcfqdbMqgIfcsvRazQ9mDKla5RmSHjPTvQ6T287kMZZ8
Pqv5pSFDbcuBMxQNiMzYwEzLjbqNPjBpNYUcWzZU9fJgTMJELmjZe81Y7hp/pRJI
TgyzftwismQHXeRINtE6CVBlWRTJI38BAY56FPOSG2vtfaghKSGbruuXNcQDDBnj
mIBbh6eE6QHQ0IvP2vpAzdVRB73rWrHo9N3bkNoziegYomlZlI6JNSI8sznFW6V5
0e7LGzZnU/hLdrWB+BwIadYd0WkjxLgbjMRGLRrS43+CMFBxe52k1s39z1n3kkzb
rnGJ+nSohKJMOCXBhfcqAu4c4fN1odIU3jt0stvGQkHJv84AmunSORz33j2L/Jau
0NXaxprOiviu5/YmU32X/vxx51/cX+BZPqN6BIK4WPvY27wIzVAU+Pa8mUTln5ZQ
vgOE1hRexY7qCDFG3FaeccSu06t83QGcVD222rf2j0Jv3B52DDfWwErCeuB2bYAG
c2nHHOtiNgDzw+I5TZRAIhNTl+6aLOyI/cZbFPfbyldEwi3eml0S00HOAC6tKaCy
+lHXaimPEq8JX4CbUFlxqawh6jUHbb3EkCh2fMqhBFKG5D1AfrrDGJIdbfcZcOLK
9XxaxiBjPSLhcnRytYkNBy+mLjlbSTK76ad29ocKOTv0/SoguF2/Ii9InbJXf7Yq
SRbvyDdHUD3Jcg2Zj9jfF6Lrd4LLY7Ha4+2QExpVQT/yT7F2PbwtuJzDNI0d5LUw
iereTz0sRqNPGeYPrb4YSQuVLxA8k6IUa/tWTuMYmjt2/x+rQzKUttx8ZmjlvaPP
OaeNFVtgDGmXbgyOLj9NsQ28pUprWMRqHJOQskpVvTLBpnWkKi1xb3Gck7xJWx/8
yy0zaXfWGs6dVssuXSkZp/K293cE86Y46KPn6ALrIr73+bGjTrDr/lqV9VrZDLKA
mqnzEvMTC6VmK14Zb/e8+sFJPTtmi2OE3Gb2ybprM76HwDpqjz6YkH+ImIvDoK4M
/Tu0/pmHi4LiMqgH8xn0uGFkkPSuEEBa9+4Jd11rKu4SDvkFenW54EWNWwSfm0vI
oLmLUPkTl2091QMVvYq7t48o8pkNKwVwG1CBD5JmtdeVv5vmzcMMTVKL1ufJ/CAv
hgAwQEY+w9G6lvRgczK6iANwo+w0Hraw5IWm8rBf2atZIo9I/TmPBUlcs1rgmWrt
Z+/Fxh2Fv4dEOPwYQ6Ov63xqjiLR86rJtMK5z/1obQHq9N4EKv/VFVIFjTke3cQb
B+KdYmeZ2/GO1ndgjlLIshwuQEcEAd0dQDwi8y69xTOIU+NNeO7Uq+r1iKfQQSU5
zaerviRbC932og6RxZC4wTQYkhVyQCCgB6PTATfl0XaHwKk52nYtLJdiRd/hL8EP
Z6caPFUrqqP9peYFCTjdRdnocazHrvt24qigH2WzftqNSuLwSDoT4SDBglD879et
t/nVOlTd4F5uQG4buJf4ogqFS5uoR5X+HlcQI7hT3OHi0FD5D/SGqEVDZAhpvBAk
XaLW9mq0vY2Z/DWs6MMOnuOQ8flkAphGoJ/8+rT/amGsOESzAxzxgN6wb8SCwNif
/fIpIGfOj2+bqYXkb2zOvcVLG6cOwIfCRh1bbNi/nLSM+LA5lc0YcCzlBM5TPl6t
PTjqXCmYuC3IYPXlb6qZ/h11WlugcfGUbYcoNs0HOCkbYYwTM6dzZNqSSgCFt9ul
3VgHDB5jiAHxU12qshI9UYmD0VBDcmxEBCnzeTEspr89cHYACZjA/tKPZyEFZ5rH
PR0KsmWX0zqDJ078HjgAfDyYEYmTrmqpUtb1pSRGhZB5ilp7IBbTPL+Hpw+QKrT7
QuNmpJnpV0Tv7nwl7MqpwS3Apb8KAktxG0a9MiV0Orb9Q9MXRMS2DzUJbnRjlrLa
nnhn1pqvMOakFz+AQceilZTGWePT4uh3XutG7fnl83811bNFeOEIW4rGe1ZBrKhR
xD+e4J9weoqt6isGOkzmU+xQwlJqMUnxLhvMxUDTJLu3uFCpMsZCR7wV/v81SvkR
JxW4YCKDovlwFj1t1rYBx3gk3W31fkbCjmb0BbaY5oHekTUQZtMaFYqUhc6HbN1l
Lm6V6oSbFzGfzHZJy3XdkbvZ3TmBx/krbxDEgzZtT4AM8fAVoC0lYu0lwoXyWWV8
Y2R4eLSEDL4RAGXFpom4SOWJ19t6D6/eI/wahTmA4EaVBtvOhkiERb1Q8MOK6TYc
FXFJY+inYv5qc2uiUNCqdvmazfxoR1g68V8GZAgKsg96iS8wQVEsfqOYbmLkDok5
20WvBUxtxC0NJZzd2ttLyr4BV68q8/LGIjMfkur8KJv4Pi4WiFCcv3+A0pOxBImk
IERJfW7x3+BZyG8tzGHlwpXld4PdBg2HfMiItTg31QSlOGKBpZ75dooTQVIS4uKW
l7j4PaRiP/Gtx4hnlvWH2M3N7/HJd1lCNVA+eEZ+SctimApD+FvKoK8NnGoAgEOY
gFtV3ML0A4MS2DYVTKDdlqAVjCmXDMAYveM3Jek0DMPSlr5dWij/4nZ8d28/PUR3
+AFaSHe/mMjIyWW1PLwu54KsKjtYlWCBRA1YkH21SolCX24HUdAbXLAt9+3Baq1p
9yLPTU89eAnbv4l/FSjoAcJpLd3ZnLHQYlfhkCcdVAEHiOWILyv7YMALzMHPDq5M
5GEGoh+xbYl1GZI31HTKJr83Q2IGjA2Xmbjtnb+68WVM1UVaFVMvuajgJlYjXYuE
dNiEAi3cA+/+bCIk8H/6g/rKgbGyl2cbqgNlzY5NuJ7eEEigXu++f2fgXI3HKFa7
t/LWRgG6gGSSYoHMh9kW2gs4HmQGCVPI9lKTju4qiRgm5AIPLUM3yFG138+CK+W0
BC/4ENUCuwTivhIXlBufecygxUATFSLU1uWbsTB08gslSami5+v6wwbZNpmWQA8N
vFXhKOqlzL3jebOPWRFg0wCx4zs8hihgJRTuSBMJzl1w4mOAH2zxdasdEq9MzQMr
9evCyYSsGiKCIizr2Kd7qc18xrSX5E2ON1e/aSuo1R1jstDqh+A246aKZCFVfMCY
y1yv5i+bCmAXQ6EEVUB/pe9/U+bkIaKAYg0oycdg0kCMuNVxs0Lu57Ix6HxCl7O8
aFruOesJZE38UGsYtrGyOiSsrHhjyL6Rxi0UZsx8hGtbkuszJ/vELgWVpt71wu4I
Rnz7LR6+uyB5RQ7pMmks8z6IAKNRkM1saGiqOczFlqpzOrvDSe0aiOA81Jf8EonA
SgnnLDyBz6VyIS6LEjhnqdvflIsbi/w26dYS41rP4xVR6lrr1KOw1lg4QRhS04xD
aCU1FmhMGN7CGjbJGMND5FqZMbfMIyzPS45fOoZaalr+dhEV9NX1kELMy5uB+DD6
h2u2sBKCLWHNhbCZPjWN6L1xukI5nvXek9L6EJGaTnIksXivri8oySNN+jEYGd28
XcwHGeE55IEhOOmhPUJM7nkZBR8hmxay2yCJjOx8RMq9N33WCabLs+BUfFsBWDTJ
+k6cpkKDe+YeSDBGeJmG763AJWbx+j0WvGQrVWwkWF4jMwKi0WsqloKj/tyL4HJx
72xXjhIweGPMAOfDqM3Dc142yj/S6x7Bjf1ohfOGRukMemGbxwzwxCoPQXEZMA93
1P+b6rFm2ZPUYO3CMcu22TEapDEAIifRf2vruWwSZn6z4/lD0BMnWV2J4QErnxEW
IsyBD4VqroI7GKrpPZuwX+KsweIMzlN2G551k+k8i0xpZvQ1rh6gAxXiuwzKTBEz
ABDYfomKZOHMJ3IaBjWydtYUYlsKuBLVGQ2ZhSNmbLYvh6SdipklrDE0jm2Rb322
lvqt5DCdklAINehJRkymuALVuRA4QFqJw9hUXY7ptzMgprzorESqKGAuGC48E6Wu
g7MfmKmM6Cpkvamhu238rMiEGo4sYzDEGJ1/2808s2U03KB+oQMipVTjikGIS+Xg
wBM7704Qt+iSfNINWidX5357wuUtWLxAstZeiiY52qoViWgkLx1dFVQfxY9EjXAF
i7PSzWab0g4FzX5fal5lJ37TYIMHu/tOjFJGpbNshgRkAXDrD5crC//7Z+xg2Pum
+cVmM5IFg1kz+1xybrbXoDyZWlOhm82WWaNzq/w25yp1O6k/4x00o/XaPJinhBX8
r0LLfn63vD/5OV1tBreiDEbl1dV4hvAyox15H70zJc4c0oNmGOab3gWVAJCKOoeK
YbOJdEhBbSMxGjlQ0qrsvvaLiO2N8BdSow9CGNqPS5pwrnulmCNOuQJGVpwQKkk/
lidmRSY8hfWewJPaISOVJK1S5b/TyXARiAKvOOuZy1ntPO+LDaFFMSQiSDGueMrY
jLeJzvJZQOK+9yJZ/QCAc9P0qTBMyvXeK8YCuWrAfy+f4U8xC/nmENxfNA2OOwnu
ebLdVS1ey0Hq641+1Lo74XkOQSQnPdoa74SiQpQgUEloDgT4Fu/MuWaLMWLqCqkj
8UBJFbDM/iMUr4sotHV7996wBmnCM2L5ZGCbPeoaKR5Cz7gKiOvu9dHXuY1AXnqG
W9MVb4W3oPR0MM5zVA4FtHXoTPHDhFM3SG40xj+AUKjS5tBMSkJW/KG2dAovjY3w
2rRgz/ITEbolBNhi8CAozRlSgsnKH3xwCrqT7puItqZ9SCR+XoJhzHMgKD9irNbf
kzgi2cGe/N4s1BHDCCoZo/uv5nQZUnBJoi4wFR2N94uWnizPIFTtez2z5EXnvLgm
guUCZZ4UOvgIsIho/4Kbw0fUwXvZPZas7zqLzGAn23jp09K8y8KVeietBM+NiZjO
ORH01ly2/5HNFTPqxouSFT3NK3KD9t9RG32SebU1afaGKszvPnEdJ9FYhgjzH/oE
wQ46olr6g3dd4+iSB1RfkDIrbA22y/zoUQajz9nQLWDsNNY4JumwKrZMQvV6F1rr
p0722MbuhENDzxbmMSpU6WKW29Qt5gB7qTQlEMSLTINPALqiHx3t5FPBeL/acWxg
XGdu//wXguzoqA3qFh1zstubdX4lSWW3ymV8t/D8vzq6Jw+LoL0bzWPUapZFA770
2IrFZ+BiwYD0nVXLWqQymt2yK97vbtV5el/UaTHUNJX5b6O9xTy918HdNEF2RxxE
0pYwv9TpOEhqrJMVkIYLF6kL3ScJIF+oapiZPFOxu5Q24DZ+eR+L5tLC2kAc1uBs
zN/chwkhPw06548i+FU3Y+LuYoNsqGPUGnCF5DEv0vKTdabeimjpEjQarUlDWh1/
nxJ3jpgT19x3ChEruqHD+q9vRN8NMhXtKLczRDOUPGLFj3MeC/5YWmN2eEG1ZMxG
ThwYW+oCKiVBoMtugaIktTRY4Hi3me+LwvEy+jovZry6PAcXpm3k/Q8qTFeOr118
ge4G9qw1IOYh1tGwnxoNZ6toIYB7yEevRR6T2hTHOOOlXWLpsjNV0lckjHpqcQIH
Qv75zRTr/LYZEJOPFs6d1WXsxemJTQshZTbwvx7039Ucq4iGuZZF0ZQ+SxnBskiS
dpul9iJ2tLayIeqPWzSOMnBp6rw6LJ8CDyMLLGpvz6iu+ZCWAhGGulFarLJbnueh
Am9tatq8U8/OdBMDaRDbhwSA0VUo6va1RDWWEHx4mcikWipwJTFTwPUXSaWNTO+t
jxPvJ4m60qrhEc7PTaZDNeS7dCtPAEnHCb+pw7GcYyuX67cT/XGT6LOTOJ25537h
HlgpFqqbYTqcdWkvFLJIPFY5jcKNCoNxCnipRBFbIKX0cOKoDo+vCT7Z14UBVfK3
8Im3QlaNrTa2lneE8oLIV9lW4qwtqCqv0sBZmVEs1CEt5M2Xn3oCfH2KXbbrH9Du
UQ0qcLOGj9z6fsoFYGhvJbL4KK4R3ZHvlUdAUAZYSs/s9VzpG1gfClPw0hxaQTsU
DxQMkMzANnsEt9zdZhQtbTvUa0BQ3475Z1/f6tLJCD73VJQWjcY0JBhZswG2bLnt
7hYG8vsUNrA2WW5hifUbSYUO/LP8uS0ty0dSAoPKWp51nhwuN20wfTNo9LbJvCHo
xpEvp204QpFqoPIHgd7+hOzHxYM2pPQu+PK9rzalVqkLTi67uLRcAOk6pbobejhc
X5g3mSnFGqlhPFcbRU9U4I+Hf856mS7Cl67RR6OnviGWeUpYWxfLSVWkzlYa68Tx
PGPnYY7C7V3zgrfeskmZ7Np8f1ymNGV+O3t2cJDOgLl1PPD5CXOsFdPCHpyWsHIM
azvMrpBXmyjVWewd8RpciEq+piR/1sv+rlTH1JzuLc98PT+TvGIrxwO7H7UYVq/5
vhLJCHi/CgsSlXO1IysmD59LhX2VFfp7C+qfsHbqGpshH2EQzIbPh4KIFKNHsjp7
6G9GWlmXgDuKBe+8rzLUTfQEQePqCkkR+eKJxFpFkkvaG7R3g4Vy1IGPRFtMq6UW
5+xNf8fqeXS2ZkyQvO8Ou2q1KBHDNaNBycUHg4w6hUIW2OrecxAsIo6G40kAWT5a
vtKZEVbOkP2xjnjXbtnRKL5aArH1VaAAK8ChBvELw2hMUwtLXOCPY92FHZ7vr14P
hzFz/HsjOeyBR7Ah4fw15ADd8JtSCJmRob2A/rmWRF2d7NIZp+3QcVTc8bcK88Ql
m+ePZLUwcRo4B7fS+cIG+WbtmRashPdrfZ6CEuXxd9M000wqPA4RPODCqiIOVs0J
mz1DTTJlZVVbGFunvoBPl88L+Hc1b05OgLX3XOHTZKOYn7f+CWZAsWLMrAM1W4D+
1spvPkmyxM4yshKTi5NEwAlO+R5N1tefh2429NsaVKVkrhFJcNEjMAdTAwJiRspZ
hSGi+7hr/8oq8Lyua3zhxjaJ88a8HlB8GMRFC3T7a9kF524cHqGWY2lSX6vPLx+J
NldSoyXhEmjomQBHUupYUzbMcLkaw7Be0zySgsi5BDT2hVSMCKAmf6g2ZNoMTGGF
si0FZe6lke3fMTVjEamxkOiCAMK+IFtirtLhBDirYC1CoeTRfDYj48m4cs4qRiDK
QjZn3Vsm/zzAMrKTgrMQw4jsmaLZLT8nzs5pOHprYI2wqvXe/apxlA4JDye+Chlm
jRZpHdJEr1R4GqiWdo2CaQej0Qo36xSSyw/iz9xb9UtN04O6Td2sbwOhgG3+xdLe
jrn1oRJRHaVHFF6D9SCkqt1CiwvvARCoxIRRggU1Ux4ZgXDOW52FVmMVuO4jHg1r
rf9Ek4lQOE0Glqprds9EWAao+ZCyRD8236WNAfsMdKpQhi/qCjkDsyez+G44IHGO
G88xIgruM7SuJdr8gLPVfl9hq+oSdx+IyQ2D1rEH9hRavkAiCDc6+05bybPIrcH/
1Xjo6G2yLvy0dEhIUkXBMXDHFRLdowgX+YGwtzAL7VGYauh6WMFsId5um3jyblG9
8AhWpldZCLqDyCtxs52zaOkkl5kjzQD9Cji6hgvqVOrce2v/ZA5m7ZDK5KofbDeu
zWBhoMi78NndS9KX8fJmwBv2R81DhZsvSsQky+V+04tA7f5W4b5DXdz7Ox2rwN5H
qUAk0SDIqrKxjbzpvbA95dvavTltXmCftxEXZKaK5GxsRGoc3ThLIwj0apIvu4K5
slwQrQSsCAd/TpOHl7Mb8RsYBTAxycmkSjCckxv4DrGTkwKA08YfzkIqGrOqD0ub
JWJqtXGM3g2GjOryprK/K83xeL5iPF8bOuKBunqB0NXsDPg2HXlRHHCshcXNkEm/
VfatanHXCiQJ8QqIUMglBVia9hdQFcekBcHHwXNGAb/LnvrNwsADaQt5WGweQiSg
wdVm1auIHaBBwuIJaJ9TeA7AhoVz7puTigNR4rRk0x7ssAN9ELRSvYQQU9AHSYaH
hfLNVYdcXMVOKUp7KW8e0Rs8F6mTVpOinXoeoERckL4Pa6B8lu/ypZwJioRjN5D+
xZ0zHTSkU2wXYkdeSgCVoSYEll/J0RqUEIUUIokeFPTctDlpzNFio3sj3UiJuQIb
DXp5u+K4Idar54f6yXZZDhkKX9LYSykDJJvbalqCcwXCd2eAbPEW5fv6YRywvwI/
j6qG+L62HZnHy6/iZH1Jm5GL5uYZqEUeCVsih2O4BEgU3F90WRuop0PxmVM79NYA
XpMrsQcHEnZAVLYLKit1v/+XHCwlLttBBYELI++KKcEFFV4HuopE/mA7Q4LEeKdl
UOXzQyBB/XTBygio8ifuwXpz63BetOB/Q5/PAyqqRIsV/La3s3L9Cev8ZyrQArie
7ClRY33ctI+EBFpIvdPtaacRTMpVf9IBy0hRUfYOCGMSlFkDtgiB0OElpqdU7eiV
wBep5TAlPKmtyOCTPA5T3aOddp4KF5guj6OoEFuXjPB77wqwWxvtYlnAP3xrgDwr
07PN2vVG7oeNGWml3M3P0nO2agHmXL6AiytzFySczDJY0/eLYD3NBE82Ie9Myx+Z
6g5JCW/GkQCZu/BB7mcf6wTuqpIdwwSc2yzbFOuOxIb3pElzqQysP7JsIUMueIsJ
O18xK0Uhf1MQJ2Z7SCJcvCPtLp27Gx66XNxE2BTc/Sre002T2cXfDTE4C1/QLRpZ
d/wBBlzCR2XtMD7rkBfNeSPUFL+kLVFKQ0ByrgpjtXA46rkCr3C1sc2LZ5LunFjN
y6HClnJNLwOXggJ8aCqx+RyJbltIDkGZ6y+EYueB2MBxnIIschy2nxZGyxee2cxa
phgILig9zrP0HwGNsLwkYCtF876yAt6hErtAdW8+vWjCYljplZAJt5t6JWCWNqXx
8WZUBmWyxX/giMwOWdCDhNhieKnc+FL12ROkPsqc/+em/NzR0cafDZ7ZtVBbImYu
ESQr8zUm+gW5UYtSBpZa/H0C+Bttc0lLmw5THx/vW3UUNxwu+gfPOudxUfL2eqVa
EYv6RX8Jm+LzWO2osG5+ipKmNh2ZLwGnzmL1hAfyBGq7+VeuL14Z99Bet9uDvBuY
hzN9Aydye8g7CaAxTEuQ8HdngDi+3uVWqZN7svx1N8ZH44gNKvzt9dlhddBPGfxe
MReC//Be41sR3xVJVRYoGs3+6rF9y74FjArmDDqafMpyZRg1nDK9vZ4q+eEya/PB
gcU7T0ygZZqUerO18rzVE6+QGCwNd9powgkmNZXY0oirSH+st+vQLvYOf8YO/Ptc
701BwIIyEqzAmAn551U+re6oj+WoKmv3IPhRPHqIMdLOclPdOCfo2L2IH+WhYejK
Oxnmi2D7ao0c1UX9HjQSFfGsSl7VrVlIZL33Cl9kS9y5i0+EQ+fTL0CK/MpoprVi
HkSu/t3MIKq1nemJ3xsd4lCtn0g6nlnnpvNwRlopvuiiYhm8AW5Pktx7x7d8Orqc
n8kConrgL4Dqd+fTX3Jw5Cv8k0XYthQRGfileT6GpQXDb4Fi5RfQ3S8f1juVvqMW
p+hY1Ldsez3WwgKaGE59qV3uEaBpn78pIu0dX0IqwedqVnAUYMbLGv/MllQCfPff
z+noyQUCI7kD0LpIC6Ff5lr9GKEErNoDuqmjw4dR3TO0ESKX+8Fk9/LRyAo5mrXQ
EF0PyD9UObUouzSvTmp1eOAS3YxvJO2pk9wR+NBvgvBoR0+CI663R8lQZHFFZ4dJ
J2RpydQcpDqnQU0CwNC9qT6mj/1aTIdIji7bs9oFp1NODJMSmI1kUfUNHTh2eI/v
iOv+UPd607QcPqClJIPv4woDiXP2sYEWNP1wm8Uoz7XUJTTokjvEZLluzOnWPVoL
YKJWVvflWeMTHtbp7Wshkm13xBhYh85p18Oj7T7u1azV/oXIrdphY/0c4ULv3KxG
Qy0pqHyeivQaSk63s+oOSwUuXmu3voYWblzHxoQ4Horzrx9WlZ8rkLDdmKPaKB1h
PcCFxAnM3PjPknAp38Jd79veuuvyr0wxM8o33LpgnF+ZW7jm2+dW5+w8S0BYV8NN
/ws+5N10e/JLIGyCkP18//vwEgr7yhsppvEtkPya/wT/99Z3TIxIXzo+EgejY/sN
6hSsuXQsJd/9ehaGfbWxBRDjtKryuuRmypoI96r31E+maO7vqvF9LzRTnXqaaYSy
zJTvn+RNnXGvTzjtAn+JevqlA/iWcbPDjOPdPKO9Xu2OxqbVdGrjYny7rAK7PcvM
fm6idkKqc4ydvluBCvZ7PjMPdfN7kZzf3Jn2x5boLhj0mvQsXDB99s/6WJjSY0b+
iWstr4fwMOkatzZMgDrb+gmBZCa4i6+EzfhXwxBThcsFCfHaVFQrAjisYAtVCRkQ
yEJJe50FKvfg5Rr9sr5aN5omFnND4NTEIuAUrYGzqHnM4NzeKj0CpBmXoJpRRX+p
KexGDaC/kk1yTdnnEcqmyQGBHPNCbRmHwoj5w7fsilpZkVltmhrDLxrCXbdmxmNF
J77ifbCnLl4dDMeRzWgMLmRDkliFtlCWpMPbHDd7s/K5axKSlsVaj6+OSPxz2FOv
vDYQw4z/yOdYJBQSIWx6QrxuZisEDYKMOqbGahPLLWlo3THgmjEG2x+RxtgEETxG
daE9shaH/1wW4mcIulH3toHYygYhfFsd8YwLNDoiiMniw7VK+pQH4LW/ouoI4pnj
063bdNuo+NKi967oyHUivbDEjUyOcWxxJX1GONxfmGLx/6BUXv5ioO2B07L+TWLj
mJnu4Hh79PBj8bbovGk7UPC5LjkGQ2nPN8gDrPsBo3SyGpruh1PfRreaqAtOWL0k
tCUvIaZIIFAGkt/H3mSP0X4fKEu5XzrKL5Z6MDViFnwsTmxj0Nf3w8Ux22VKWure
FkLTFUx/I5dWc9doPIv3IqhkrW4h7Ozk0oiwJtzcSU9z1tMp043Tqk6XaQh334y5
pIZTTEYLzNZk/+BW0g9Pr9oMckaw4iydtBvh9lT45MYSmUO5I41jmD3saYb3itKA
//PoWNBf7vvenCPsIIwSxQ3f7fX5NDHPy4Z1ASlA2mGzL9r3ksLsIse3QFG/TEFZ
2F4EQFc4yq/L3Q0yzv7cAiKTDEumXG2Us4G8mTy2FJZt8E9aWwgVAYyx8OFc2w+g
SUkpx3I5Q5+BYDoBT7C7RfNXxq6SdrOON9VLfyTlcVfVaTYGOwcM2iPJxAYMYttl
YnTbmqZxnen1tQG4e8n1wziQQ87X5Wvhp2ACLOv5nSD81nuXPGz7XTsq4B1MvcJU
lRMEtPH3FDAL+EW2AJTMBgjNkLF67c126uftCy84NruxK9UejUPpE3pb7hZvyWk8
zxQM7CE9G+8EX1t93Em0f5EnZtoR8lG3BW3LKzXVtkMHc8lTNRA1u/IaVZ+czbpB
62sLV4n7+VeKGNkxFsUBbOmNDs0lGYteXFZ9X92ZS162f7vV1Jm2cUuIy4fhZUBB
RmiClfWWGyTPZWJJVQUaCW3n1N9VHtgSuvtcMn4MVItdV8ZCjBA4KIMTGkeR3MkI
TdpqNOJzzQRnW8DSebWE20cGsOD1qub1Njka7y4XhnATUScovpoDETsrIK9aTk8J
uDtxVcnxWYYFnT+ccPQyQJFcM96/d7pO0aVFPbCUYqOBferOzjcsLSRlqRKrAwaw
i43clpXadQepkWBWWCq5H2ay4jwq8dpqidRDcWYHN8HYw2P9djb/wvfDw20zJpdE
a/u7INYS0dmtesXNVkk7EUfnFuVRhRDsvfFHGunPwJpsWT7DvFiBDx3GzGF91ala
VvRFt2qDB8pvYk6seze0wuFKh3yhsZz8QiW13o75DWFWpxXLjHuwxJpGyM2Il/10
Ns5HvC6dMi5eu7xxzWPOaxU5x3PX8kT72Jnxy6OfbcGOuk3b86r7Pd2q6yASvQfO
miUeJ/eJMyC+EP711/98rCMG/8e31xVUavsJSFvxxOGtAFPNolLGl9kzHXQb/itI
Q8lf7splT1rWLtv17WptqfEJ+WZf53CTBEDKziEnET0VqOenxDLUBLtwOahMGSiF
UZIamnSmHSqRNNDOMoX8Mr+zQmUZ/LhCyIg52JMklvApKm+ERwQ6gl0m999KwOkm
qhlDF8KsPeghusfej6yx8ZmQaBZmk/TjII8/sSmooCR0XaQ90FJXImAkzQqzfi80
Mn1x3/RAC9d0ElzSVa8dDPW7k4fkD16amiU2+lf9IgqbNnI+xoXID89WcoM31QtY
UPMh6/Ug4wETZTRCtvKndqMj44imH/nnt/ANdjQ0YhP0zB4H8wmOb3g86szSH2bA
iJqOw0ffhCyFxrkMzBnBRR93flw2QkhU9AGmE3V/gL7WfNwYrZwLaNx2vUvpHb7C
zDTWyEKze187LGati08UHOhjdGi5ssJtUjq60wOEVAPLX+RUA2xdmpMjnQT9jjFW
HEOfHuGD+INLt0FoPL0UCAq2EytQ/IRQvLOfudO05NmFD77yt2hap4PE6ZCU6sFu
pQsKd+FfZ/6PrFYKf/VyXrsg9CHzI+I28aR8dJoY1qI1xu8icwIxMiBYmYqoyctq
+VqmXilxlOP93LLp4AzkSN6Dqj/o82ij9oFLHfxHMeNDTQYLC27baOLYNyoYhk1+
l+IUPVlv/1JUgItiLlpef8O2oXk7t/A0vkcyZEB5gNg+9MdazIA0R4uSY3WMV1BE
r+OOpvUlKWtXw/YX5g29TQFHGjSDtsMUudBj2xiHtL9NiLrV/PBD1ZvznXSIOcMS
58XwhzkdcAqfssiHF+NPb31cg5litx8OwL3H4hPEqvigH4g/I8LXkPrVPCzdZCLv
69AHYF9rc5iEPGRBUXPUqiUBy0/15c6RisVXjNReAsvMo3hWgbttQ+SjUskiA2XT
yVbwqfCFd+q66aXXWakHQUNoP3tKbBGHYJW8jXD+ln9cWwDSLCtVr5q3xo8ALJi1
kBb4RCiEzc+Xt8MC3JFpzgLsPa+8hun1syhF362afMq/8HkWj7ZXb38LmUKu/vDW
Gi9x/dgTVLV9y7J318Q7o7kvncMeVgvgFe1mbmr0iUcYlCyBVhtAEZDHQQeZybLN
b54kV1rY9EwOLY1nEu/UIthAuE9XuygV6fVyP7DSr0eCXUm8DV8U4J9w2bA3TbbM
PBjKZdYuWtws5dBy/vJx16bj/MEvpJI3Ul8pULvi0C84uO5/yn+nPHY/YWZh5psj
uECqUUfFh2X07BDCOqAJaKK/BkdKvCL+d0NRI8ex0gx2kIsQHFqKKqqHFPwLbrEj
udCiQqOVdvDf6QERL7+11vQyBPNgtwGpRRUTL6pNPaKHf8J8zxke9c71viEQdA2h
OAK2aAMX272nulzZ/1ls6cDuvGZbb037s3NNGDyzcwEmBs+kfDOKXX5h2R4LasOx
Tr4ScUnXnKIVg8uVmvRKogZiIE7pnYJNdJHnHk8UL/ZA14fH2BeFm8UeOu2a1hVM
LRV+jQCwkwkbioArvyzsOXMo0oU4TdKJZ/bixq4DaXTuo+ZnKew9CkqLsjWumwz5
PKvL4V8T6zL0IH4DhL/NRyj+vKGMPM2nQ9ketcZBlV3PUxOwQtys4IMjY9i06yfE
+tyojLG9wD3g7bhzhCrQVaaig8ds8EBhZeuKKh1/c9jR7Wxzs9cfNVHBNdAi2taJ
tVN/8mU1uABwcUAg/ciOhWhbjsJEjzNBPBNGJ04VJJhZfDpUYksTdb3GYgFM8rtU
gJmzbFjtdtiCfTypFS2VR053x/gBRA+DC7ivqv+s0rV1turs5i7IdPq5U/Kf6c+O
LGbeUg49xOvGCKbGMB3NwdqGW0Jo/9QvAYXzKIp9ki1QXUDzp0JN1HymL1q6h4ET
Mac8/RK/oIdEseFMs6tH2V61+japdHa8hhI58IZAqHFC9roRh+8XU1sI85y5w5sa
9H3LyY+VkCf3aOwN3ZzFLlA7LVSn39XMSVkc7eIECXTaA/+LhK2J6wd06jy/gyTH
8bhup8w9uoXRGyKJa0qun/ZlBwMlyuscBmDDThfTYPDUSZBw/QNnhPJziHCnqzEN
aq2l6E2RUAx+FF+s0B2XiWhFOBAnqNs/HLTzcGaodpud15WDGYwQcYMnnJq811/k
xSZfQ3db3PjrbUrlDYtQ3uhLb1PWxq4tGh+9Ytj7ObjFCIhNWIaDGy7CEEdMG8l1
OiqJ16z/hoFRjxa+4qb/OyMOdSceoHyCvgIrCuR0F2M/pDKWhOqbDt+/KjM5rukH
EcDi8ja8Gktjo2gtrggFm3OrGoW/k+R7BZCD7YJ7rhR2aFeNToZ1JP96E0pxRDmN
6SOZ39IEoC21lugFwhuH9F6q0k5zQ1N/x1gJdcJPW5tJXRKjm6+/ON7JhV4h0Ze7
SWc7Otpht40+KvlsUaKOEv2fT5Hh8/sG022FwsnnYRPtu3VvftO6+X0v6iEhg6/6
dQbgVdVsGkXOQRA7UapHH6fCwbHJ2Dv4kgRvEtyvhjtqvnQSGEc9ryljEqhrYOIt
augnv6rPhp5e0OyvTHUqfMKyw1GVvBAmqeixfBZH7reyyKWipHKFiKdfzvDO/cEt
068WUGPCM2Mnpav9JFAuPFgcxXIi+mr89cCJj4DMZPV8NQ0miBrwoZz7SBFjqDfo
XLfW0keHcjM5uTO9MR6N0YFDXLS62xEkgYuLH+rFxhSxQDJiAom8ikYhFB4zRozc
Ws1mxZEbq0dbpVS3AwlyY94T3Wg/T+3rKWsGyCPuZOhLWtq3ybPrJghR1itOxgKF
pj3NjBDmPcfaldTI90AyYgvKTD9QIlPTAqT32Q8/bcCZ/A+y2/Ysrgw+8w0wOa7z
vkrF5avnqR/Kj2Chg5pEhT79kgPkfo9WtD5SX5igIE+ZuI5g9mEO+CYdU433wPNg
TNvbEILrKj0NhM0htjLZlvyNkSdtxE3BXnAttskWqCLCywBgkEqKUpVkgwrpwZd+
v/P8tQRCcUcc8Dh8HdlFdG5L2pLVbRE7hG8+zBVdFvXAk7QOAgUrenjAST9u4b/c
yxlLqL3het8jvjL5Cqfq/dqOCh6eLQFAY7F9f58LNFbGjspLSZntEvaoVUsdD6zx
OWHsMOAB8ntXTj5l+7/AvbXPNUGY7wsko8tl2GL6S8Hi8HaeIo17GBqGXSKRGPgq
uYpd+6hHYtN3LeMTURoYl190kLBdBWje5jybYuL9m/J+LcQgvo1Cmmq7CovdknpC
axBJy2AcpWUBuYB1E0hPJZPTaRSquMBBbm/+zvKKOO2QWQIaMtWlzXm10K0RXSem
RaLJKT9476R+yqXS54JE4JPplJ6Wt1UYzBVtAIr7ULuY41alG23LnwtV5cURP/CK
6S+rgXLuALfVSC5XMrHPfCA+65NFwHQ7XDnyA/Qn/9IIUIR//rqm3unDHKpwYtTh
x3CVGsqV+Y4KVj1fnG7+Shvn0tVOsJRPrrQpEzAFsk5sUSUFXek6BpGOTs4JFt73
l4Topvue81IPWID14jn85B0E+zxpV6tGXYaGXpdisyaLyLR6bcNycBF+yHueUbVI
2hxjK8lCKRh7mSC2yZy/+gMccg4oghNFD+LSyDQcVqPaZOMjWIUBv433rHy6c2DA
gQL8ipzpOUPFw5upDMaZJjdIEJ+NiWaQ9zMQm0JbTaZRZ8visgUSckcCUi/W/Ypb
1ITTAv/gPrNcF0NisRqcBVFfWl7cuG4zYxt8cZj3dhPt4ogcIWVr+j7z7zRirwHR
1tJSpOyDIeXj5JEzG3e98UXyT1jV70/nVy85xlm8rQoYw3K4fQLZmGaZbe6FXq8s
WYWwhCdaS/4aHzpdi4pC0UHnD9R8bujr12VGk1qMYyEkJF7EKWQf+VUBF6JyAwPP
EUwuGcS4OSBK00e9O4MlxVdds+z98pBPsjltGtrlxp3Wr6TjjZb4tOoYBiSIcxTN
W5Dm0CYCy5au6V8cINTWOIo8vuj6nevyqlxzTxBwuCJ3AcykWAH/oosjcpoKZzmN
qdCVx7xmrl1UiUv9orqDWwroLQA7t6IDEAlENZwSInLsFf7hp/gcGQvoU5coWeSN
XOkZg44aptBi9KPSAqKlgOTAXRGenf4HilOPHl9Ai+4qFtQAKTaYko8UAfc1m2NM
vFXeDybUKuhxw1h1Mbu4ega87Cr1C/0PaybMs7xeK7dian5RjqhZOIXE0r0EJH84
vC+2wX/hZB+yI/F87H9IqC/hbwWdlHZmDY8L18qGXgurRWOJY1eO+EitKQLgZgGk
xatav5hnvRke25JeWQ4H3HZ4yohfIb01J8TieJGQTHvLrX9hgsq+BVBNipsjlA4B
P5J/YTVQ5CUCIF4/lMxu8CT2Y0UqT1gumFeS+NdQWrmhlGzmpPhsCaJnQZZfyAYG
ott4n71tad5bkghtQ80p20aru6gPBAC/McXkYTx5hWhVPGbVZQPwdJKkaEBK0IQ7
uFQNqOMGrPTDkziXcX90xYJK2x2e7tAAOGyMcTlY6rSK8wEC5C8xRCIjQIxDoSmg
ptUbnyA2ubnRlrYzqdn+djpUoYeQGJeSKu1yNOWCqc9e8lR0qyjepsDsWkscpUd7
sdgIgWoNgXrbqGUihn3DxH7ohhLPvYFj1TMKHQIxnCw++HXMzwAR6ZyTfIe+zcDH
9OFuj9I8sgBaQo3UdFNoLZbG/jyzKpALI7HdfAHAXrlWVUCwWsIIokCTOTkR/Drf
utEEUZARPQryVrSvTWekryUPax2c4GrUbOeg3pmKTaFVhGFi4yLyE11Bb0G0I2ea
MCSl8hLz/UksHWzHFvrBuMwvSN/utTIzbuYRTaDp5TdO68WIrfN7Ah8e4gWaRC5f
FD7gwjrtHvoCj+jaogsgkIpghdCaB2IhJGLmGGm12UZUPW5qInp22dNyjYZKp/Rl
4EVpw5rbwwzq7zBsbhX+cg8JiE9chTLoDxAjOdkBecQdz3jCKJWglHEXFveTU2cd
aBqufEAfYxPK3Sd70XlfUb0luA6Z3OGk8ONbUA1W8sDW6DzaU61FHuJbWggpM9xN
NzrCWGnY8MWTi1Kn8bACUnQ1l6VCxfhov7c19aCPMEcdyUANMSvxSTFHAuQPw9qF
XNZ4Q1gyoJK8EOa+QFLTgZC2AVnsC6MorlT4zzyo5J3Bpcz9xi7xJKLyKndSPuBJ
j10BDYjfeTM0KUevqykcdMSbDfWgeqT1hnjgWfTr8E9Ll8d1LUyeP0iVd1akezHO
ucfyP55nXF7uxjxsIW8qY5yxd5O7t7ZIifD6JxzwtQt1rW4FvPh5goQRYjE1UH1I
LJZzzWGAcIjAWSBYRoy1q7T8/ST63nr9tY0TTmzj0f+pzy4qPwIWmCI0xfF6J9Sz
5XTPAMLPc+Q0EtpTnDkuFV15qBbupzd6zP/86VuLG7ZQzET5qt2QINmRABluB6p0
lGpPBB4DLg2ASICEfSMUbhi2xrqCPlSJlFRPkxQvCy9BNzuGasQYiJC5M7Pmj30h
lE4s42La7YAte2Pz1wjj13yvac9c/Jxgh2OUK4iAroVlw4FOCo/XQPdt04FrA9RX
Z8a8Kv1Mdj/o807Bupot3qYcZDw0Mmph3+379uWOWiilZ0Q/4DzoZxr9fw013khT
WmbBuLTqIkD+FekWDrtymv29oJhpQVdoZJNV1MSpz3wULdbs8pOunygAbURs1f2P
nJ0vhzxdF7yCDSSdlxs/KfDsn2d2IR3AdgwgWXc0ZkHt2YUndyHkjV0E2WArQxtl
ZRyAST14aYMi5wZrmga2FEG4cQ45Z2CKKTvZU1YEiVPy9jMNzXpwr3M+9bSuwrWa
C0JwzpqL0YcOx6E1HSE3oePHgpFAGP2E0UOAcCSU0TNRmhOipmwGF1No41XKnH2W
Oz1r4COKK4Qm5MUrH2847Dqg37uFp3YGl0pcBWi19qHHXtPV7kPrtcE+SOmwtW0G
oAmz1+TD46mKb0i9uG2WNtIAiwGarXRncrstq+rQBWgcifKYumT8dPbs566FkTUr
rNryT8LOXh4W0XsyZpbDmOBd3JssXC1Y/F8S0dUpAFq41QgV9lmadTcO2Rpe17V2
fFFrNh8SjMj/M0A+eqWsfDdk3mXs6SVqzP/+cBzRjXg+Bb0Cl1AG6XxedaMYRJo1
0uUBpPhf1ANrfzEuuUJvzSQ8RMQJesq4cDgl5BqNqSiBYCQGTTZuPqjjosQlsy2e
LqD4UnNLFs+3chHs4dWIZcjo2EMCPKcySWFG1aDGVYzHxvhnj9dk+vSX7pemyaFr
KRQKtYubXkaB529wtk/Mi+JS5IYaEbIIuCQhQgcEhjDsSbLvbH+dK5iq7PfhL9Ok
O7SHsg6MTFakWmaEUTe/ILElmHqXBCHdapqxyMIkVkZdbdn4hu6IpEVmIU8Ou0zV
3LJSgcPYjFd1yuHxTPgZUHXy+vY58UKwieykXFj+e9p1ombW1+c/FcupaLqY0RDO
muL5XiFg0Oho+a1L4xDVfhXR+aXe7LcRnuKuAqg8CEvAQR0v3F7pbvvdeBqmqc31
mNjERfusDI3cEPek+jtZSbE84aLZAQ+AjqyWpQ5i7dAS6gM01zEephn+hBlJZhhS
MPvAwNRADE+5lMK89U6K2Esz4jjN6kGL5erHoneMtHTZw94WpF9QZo60Ep0mOV1e
4zoMgyIRL5939ca709HH8H72qpiyaTCSUsp4ZiPDhTFlrDLw1jfnqUX8G7v9m/AR
5NfD1OO2kLfR6gEvJU7hWmFyP4yoxJI43GFAxVmWhC6uNnieapF73mDthfy/FmF2
NNziu2+qd4rx9o0dX/63eSxsfQ1AUTstAuP1p9W2HY/FkR5QPQlDywzr5ys2eMXm
gO60xPX53hN2hDbiISzExO0sfgFWmR/kWD+u0fAkiH6gYA9qSlGkFMKc04AZB0mn
IUphtC7DrRN3REBOVUYk/8xofXX3dtme2fDIMQAsoJc3GZ0l3x/dj6OHXHm5kWau
JQpmFwS7N/6id9zYcxBhC/MXXiLncEn4n5WZc0XnNRCF0pbv8rPbvldjSxX9CAJ7
8NtwI45RipeaH89RcayHIvx9eOoXdIyt7zF9kutBY/RlbCV1Qu82wtDxvcPb4BDN
W61wkyQQG72b3bh4qwTBxRUUF9ghGOXg+CF5NJWZ51sJwErRq/p6tc3USzsN+HeE
rKCqo+2u3/Ph9hf/rd72AdHbAEbBiLF/4XHLccEw/Onso18eLE93tAoS8W55PavO
yVMu5BQvZeUlTtb5crvO2NjcgO0SEQ4M1nLVPlKybWlJZxsR2quAoPs0vqmMoLQW
gofSQA7+IdMhnJle9GYyD+Orn/EZ+zP3M0uGKo6nxxu7Gos2mUjafKzEx9p4hIxe
hlOv20IAbsM2iyrL398p8gIIbrfGKLlxh8aeDTB49q4XQXpM3l2kKIKuOkUD/Osx
fQegWPUStHDnycMBxpsEsluPUeRmh5aOqgXDq89cF1kKJaranuwHuPa0kjiuFAL3
XDrWlgfe+UrzPttHjEEi64Utp+1xj/rtSqouCfVMYRX5p3BHulRAISLRvEjDeNw7
Zs+AjGyB+xRNVqdsvGHmcxoACKBE2rzEngv9w8REu/GvzxgdBQR8K5UpvjNyZ8Mv
NbgNXaHB2Tk5oslelMwwcHwXJ5H0gJhkZ2gqJgRuHREgXKYm3eI3LMQyJnmABGjc
fWN/Mww4Sy/t4LJz1H53SR2Wwm3xCB6EQXDRqxC44ICBt3f+AN4il1b9yjBII/km
snii06dFhoAJZ9c/wRazTcCrjxbehzZUFdnnWxBXSJLK1u/csAFvFJxhbLFWNUDA
JQ+5LsYW5dweimDBpN9qPYksLU/F79WakD4UygHUu2t/H/GLLqoI6XwaNOZZN/cD
d/u44nUXDopX31xPCSWDtiIiaSMDAr//00NqZz086LMt0NImONO30yJcNkYyE/ei
/tIJujn5h1iMBuMaeFHxp5nCaoPaDbcajbDiI9ZFpI34FHb5Q6O5VYzjluV4dg7e
4BLyRmIU4I38rUj6pia7o+yZ38N9Wq8OC7wrLxpmtK3SzhiskX+Xdv4IOj+vusR4
u8VscEiAldpBtS0hTfnVDnZAHxFnSNWKwMweGyaOwlvSD8VblnW4nelac0Yc00i2
HCsbfM0zBqyiL/vWTXCrBtUXb3kcLUbTv/HzA4s3wibVoGT9L5Qo+g4BZq70CKdY
bDw8cXr23Ue11LR+51C3x6611KE/18NVsizIawjDzxibf4lEE8r/E2tDLDLwQdOF
ADG9xKEH7DiOG6/EVSVzLbE6hJiOZaoNxnmwPYaYw+AkIga2vo5vU+OvzW6I3XQF
Pha+U58F4fEgaYIVwAcv12RXw8BSuz6PPokEcaRzKgHb8CqNxg3LDfdFt2FQ+Tej
Jp8K1WzBn8HOPzD/g/EYCrAGeBncrsnh/tB2e348H9Rglh8GgnVhFR9IZPFXWqPu
F0zJLBtg/KNeKVJO6lDiye10qhoDM876Uqf4iFwP0Gy3NC/lrDulda1Qrowm/9GV
3FnnZ5oGvfFWbxGCsbfqrN5mX9i4kQ2oxBBtYzuh3vE1JFQItpQkMYSNIBQrOKGq
nRkBjMiEpZOJJOH5oQHVEjDfS/hJWqsnS1Mt/jkcxJJDCcE7yGHeIA9abZ4TobBE
s8pJmcOEx9rt8yaHPeRuVluP7kDiOg3K+AflJK9YMp5iCokM5iCdxuRPRPKla8ZC
NIFJD2jCq173GpqEA5jsUStabZgFSh6DaZtnapywbL/PyvfNTvlBMeQnK5d5Q806
sO696DJRCOMGLxRCYsh99PfNhDmhp+5s1yx8c16e14P7Z895FV+tpi7bQasLWYDi
r9MA1rZZhhcAqi1r63gB8or9kptCJ4NoxZ6P+ZGE/J3ciEJAN+erRoMf0yVjcUEM
9QR6QaGwqfxpQYfPyV2O752kQ3buDnkMvAR3fRt1VMBEOo8MKg+HarhbPUwGGU4B
Z7Q519NIoylmJd0H3J0E2PMiaidxWNpif2VPxGEVVHV4zgUNAiFHBPG59ZjzU61M
QBNL4BGSHUG1bQnuvvZmuFjV1scKZu7mEYJ1aW4RjrbYfi9kiTYtDFBpgyiZ0Rjh
1BwHIn2DcipHHcbOqSIc5m5ur53Z6nZ6rdgjwkipXxK54x+/MGk3Kok7HiMQr74t
51UzuOQQQ7S0i98vgUnDwUkr18SagSXjitojyUq5xaGwjlPQAM+SJ7vU/dsrKPTQ
v1BCXRzrYcoRo6N5RmayeermnA9i4AUCKffVP3f5cxxX3AZdE5F4GjjJtWQHhivM
M5WYouxgdYtJjQ4qbf8gKZ47xqdwDlWQfQI3LyDpXTTGNHNrP2/D1tQ0iwRAKuaa
j7xSEH7moxVXVpvM1+q7ZUun9LZQ9dFUlt2kCyYAOurWiwL4F4fx7SvXoF+apPDz
BAxeVkIiQFd1YoHBifdpV3ybnqFUV73pku6dZGAJHRb/vk3jGWQuQvJisF8eA0kt
egOgHkT+NqJkaz1FWDbUA9J0QkmOHbsI1d37h6s9o1INSxWzVog4BJo72RWBTRFC
0/f6LjN8w7NWQJXG5y94ViwUFFGmCXCxcFt0D5fs/IM0+j5HrfyrKSkMCGy3Mic1
iM8ERU0D5sZuRdp5x2QwWctGvnOiJrF/E+By5v2ZqeSJBLt02wg8mEvK16RwUSI8
GHjrJjxaQA+wqvor2CrDc9eM/+OmX9AXZHzURWov3zjcx90doKn3NC05bpYc56WS
uzDjYHdsV39aPRrJpwBrE1uTxRr6SASvIzY1Q0qPoljMoD1MRgqA7hkeuyzIdCQy
0+fTQmIThn8FF5/o8Z/3FoHgqPMJSxAmHB7QHxSEch4ATJaOzch65+QxD2SmJ7Hx
hLxYPiNdJUddfDuvohJNV5QaycekDsuoRL5CfcJX9Bhw3XODQQpG/Umu5joBXs8F
W6+2h4IX7+nit154/B1jz0hL/7Uiz5jVZrT2S24pNLRNI9O4FG5teryzCzjKnSp2
w5nVYqOAqAy4CzqVyItFp9a1bnEfuPJ2DWDrHGmTp2ajEGA4DJO3XTcx3i0LdF1o
B9SkWKOUJOUg7T2k2imZJ9rm4LvJEj81GP6ACDB91e1U5ZdZ2PVF2mB/1oO2iiX3
m2h+nhESap4ozDTarLCCjIxKRPMlHd8g9AqsZJybPdnJyPoHdPt8xc3WQRHAuicL
nh+m3EQMpKukE74tBayRwYZjvUz50M9sBTOKDfDyOTCLSE4ytK8YpC2crskgxvjn
sYONqW7hzGRBlOwcEDYpopHfrSgKKixWgm8meM+1hwTh+HEbaxxBnpBlI6u/3OUB
+q9CUJhdrY3bxwAUwLvkEvzQPXbJPep2qOv3xKasXFb5CQv8enKLEbws0JPbAxaY
W9e1b44kR/wwED6Y2J5FL/IpY64gU5QergvsDnTIIqOE3LwXxyX5C99Kru2e/Xjx
wSU03ScZ9JKT4h1tnEI+LY0KvocgwXuS5WLs860iLH+54U2UgvDVUvymE3GniiLn
AtoTCXzQjY7EtIoqGukSj4G9yZDpaHLmARZMsGiIYi3kagM0PzuKPMp/LGn2su8S
gBNQns9KzdCNewyfY6Lp84LF4PgmFKBLeVVVQdkbIxmGQzz39ItdK1CeTyVMjTmO
LljkWw4anZ0d9L1LPa9zkIAz7Gfwio72daDTU7SkEd8T7kEbb60bZz/82KlHasmL
bOOzPGuuWy0HLrOzY39VXh7Dlf2Sf9uw4sPOq6PO264K4TsuReEWakP0o1vjDy+l
4PJBnaoegMmo7ZVvfZpHpGePxpGSz7PdkSSsOiB9GVUUwBwCSn2BxeBADXoQZ/Yd
/xfIzdoinPJF1mmh1qc7xyQhCVX+kuYJe428Geb5d8TaUXHQqhhsRTIYG1QpR7/w
ZAATl0BXACDCAhEBPAYENd08Vaqe6uT6DGtwsq4kEPj9sJPudMA9FXxHpy8DCLhQ
C5WHIF4wJrS2bkbPelmDRHv32P88n8/xRbhLpjh4VudwV9FVQUe/tGEOFp2ipD7L
H09S4u8RHuMzkK34HmP2Q6HOGam1xcS+7ZQ81unawMq7UoQO2yzbhLnItsOHU+Fc
KwoJWEVQIsbRxH2uhU+Kqz6yNrSNDQoR+jQP0Tn+GeI643okgKW8V5CaWUs5HR4q
UEw8zZtbOpatBkGxIJo43b5PwnwHJ7hgqjKP6cKl9G3DgvAL+hYtzv0pb2JAWwxe
hl3nfGqWjiWI/RaL+JjJOh5e4hqJpiYFa+69N3LrNRn3XdYjx6bdwxdSSsX375Xv
u25/ivUZb+TZ/dBRJbUD1Il2OG+1Jkt7OxI5cCrXau9ZNzZaRxJ7vk2cNfXjn5eu
qyjGin1koSmZyCXCy3T0UjR+985uvIHYt761dMGtMfV4MbTGEI9bovAI8X5ELVWt
Y/g08yejZSK1WtkMOdH03TfjPO0Mp4l+7GI83pcGC2vft5TayAb46StGPa5umO6E
pI5YBiWKIAB27ttapjh+vtEvH8Meikzyyi1nKTcIxSRXneGs1nJqf6dIBKxS8INr
K/rRO5c+HXyVVc6rebXk98Eo5Ap710svdZ8og8rSl/90g3i6CapMiVnCua7M/5PZ
vAv/a3+9U38x4wwK9Ki49Uwt5/dPRSln17NKipwpikl+3QDQAJZOBNhPCgvEb8Qh
DxRPTiQDTEOQ83bGRucg+OjmDOJlBcBH2hvn2g6w+kbL3+qD77zSPRX4Vn/PSMFu
zTBmOm31um+8ih+lmnHSAM71dEJwTavevZxf/0ORDwIUoL01qzEOjCHJHYiaYVJ1
FEWMNhxPFqSZHqCS1eTOHbMFn2S/g6Aqu0Hlj3TefHOR7as/e8Ds6qu7zcYAjXmQ
hva03N53vtjXlP4s/d33ty/Z7SwGUPXZ1W3y2fl1litD1EkzpwXwLdEwOBE1SaWn
FJqVNoV5xbnlkKZsEztFSOWUPPzq7Q5WKrhbv57ekNtAjtjSoY6Dgi8Bzr0w9qdX
ZYFPqAj/V+oUcsnVHqPevAsPRdWSE+GlzrKzG0XMiJtY0h4TyGvQiB7qQIvYCYdG
GRvSpnDjposdYVpma3lGJvsmuIlmOQaOiJiDQgasauuF7IsZuxcOLv9CkMKPsvwf
vMvN+5OCb1W430ZGaMQv6O71n6LKfJxV4DHG7D/tSoRMapgj/kww+R1127gQz5s4
A8IKypigvuaa+kboLGKeg5+FqhgGkLQ9nv3TgIEfaXDNAH8wswE/IgS3eWdHbh66
ruQgmCsb2XG2BlqgXIrpJaggaLgGtgh3BZbNg1aHgOwfEspzLghobXt9JmYUgch3
+Icda6UEXvE4bMYpR3a1TP74bnNwTb0z9jOtdxAJvc3ecnjTFYsebwVbqgdaf5sh
y0dUmwHXVXeIzSzEYFAQkeMn4+3IY9YfcPf+Ww1YBNvqCICvrOA9Dsv1nYxpuUPp
BRUKepVTfRGlqPmlpsownRjNqtFrRBH0hrAexvuwEWAhlPXL16woAgXJ5CDXoxpH
l9/IuxwBitSv08W2PMWchT1Ebqs5gINtXFZXkeIV2urPHQnkJezAIQcGAY/uQEx3
b8YPqvceN5kIrjKjOKTEbBdXawShAYddUBuYZ7Ay9MTqzhq6bEz6GglaSf54J5ta
+8fkrpP+i/+e5cm5LD9tGiPxDTHIYYIXW7mYa23a1oWuNjFKc2XOsc/nTuE4cJs4
gK8Uxca7jrhTK2nGzyhWf0TP8w8zPDhWqEmvHwZ9rgS9Ltz9o4eg2cfJMvaowPKG
e/p9MRNXfyyBzwCWYCYPYcA89bXvumMnbQzrkBrTXX00yZugv245uGlcoyX+btoD
KvPYNlZaAifZiuN5Xtf54+AhtoaxC184tE31TWONO4p4ZUbC/QAthytOnb3D1ouQ
ZyPhWKrjDwiqaBQC7J9y5GBd6QxF0pjZo3RM8quGpS2kmBdgUV3XF8n8ybwsmlTM
jr7dkneaiaNc16sHDNfJMpNfwmbg5VAioxlk1fsi3ceyuCSBGVWV6Uf59O+LXXwr
mPOxP0Zlimiu4BeKpk//kpMrCbx1NxBr+UfoKcSgwdMUA55ySVlIaj57lGl5sVry
CUKTG5+eWH+HB+ll2hLHkCGCZTwOVhrAL4p2qY5Ef3/rf50Pjpa1ppFT/hXNsSrL
Ul8soWp5ksYx87Lh8emIfbA3LpXrKp2e5bErU0uHnA8RUK7Az1EwSxc5GoYO4tIQ
LQHnGutONOQrBuOiE5cBnZOKFQavRUMlLpw9DVf1aS8zt2auLo8jPvnmml2Ifdjl
UROPRwDux+DU6MHW6xPgxJqdd+4kgYBHfKp4LLXCi0OIof+9emn4TWnqwyelWPF/
w7GA04p2LR7NUXdQydMvJ8D65w6ak++wG9vixsGNQ+FNYjTkPqdQjpT8+0V8UQ1u
FRngCUafRVADAVKRudkI5+3AQyvBSsyfYXWjb7zqbhXXuXtzzVkIEW+BlB8uI2mc
CA7zjgSkyzUkcyN9YxH/91w6JXsZM4Socq8whcfHbKGHJmFgGi99nrkfGGsoVckb
hcTgH7Lc1U4vJSeMtJTTMypGT3oDG8g0buhN3SW57tMAom0J2wptfjlAk+upLhML
MJebHiEYgtsmpm8YRITRje8treWWKKaGU5ilO7MCB+kj6DCqYf6lM5hIal3dH3sF
LKJN1zgeSvIME9TUWyxzV/9EMa+WxNIfKt953gDtUNHqzMkuIp9Qfv9/aroXP2G3
UHSA/NVFyT6+bWZuPfzpuCXwOY0psBP3ioqGIp2be6UVQ1pZKEpMoxjq+l+vWwGI
uqfwJdXTIOJGzgZvrhHYtd+JbXuLRaHA39oqOtwrvLTqNJsopsn4OaKpvKyDipOl
NXpQtVGOJR/SyygulHw5GjRyUTUDETBgLABKiCCD6IY+31ljKMhNJnu69wRiPfki
t4wg/nj6/DVPGnbltnGsG1OGgmDn5BzcBg+hWimNlKQWazerfEqVmfvVfTPS0OPL
0v9kkQlfb5+rWfqkw7QuiKy01voZcmn5P+ugn8WCp1Ls5h6kKG6ywxH7u8sP45IT
y26cydYPuaFqulnXZT57TG4PdQZLY3z7PN0O2ky5R5rSkm4j1hc2jflMWxx4NIVB
QjxmYQH0UEnKdw3icvOQyFYSyq/axcEpYUts4n+aSS81iQ4ky0ZJrmaNkAGH9kSF
GTlPOKwffFRwoOhq7L2bQOrDo63WijD8DQMXOhJenw9OzPfGmY1mjxCFOKb0IaqD
7oyeOLUC3+J8fSs5IRBXU8lu0BGCgamLymEto2x/IADdc+mu56oCsytJptAdNK87
sASkiDhUOzs5j4dLN5Rnu6H69tyacFQTuojVmHgn8z1BcIwSU4d7rKY2iM5eBiGn
qkaqoyUo7zexGo2HPpY+ylDsmUVrQZhmbg3Fy0hUt/h0MlA1Rn2rYc/6IaPt/4wg
J26FGWNhaZvX8VyVC8TyOQJVp0beN/coO4IHdP20HcCypCK2RAF4Q8HfTrTRc7AM
e2sMT+kisAxeC14nhmlrVSZfeaXYFOU46h38xspzfSSNtUG2GSf5LIonMKbiixOt
EHBtwYDcCjnhfzunYZ2FiE1P79SG757Q89hi6RqVn2AYWsR3g8OXT07zHA0AOtje
M3Pql0pr19DyKpVDdN63QmcKEWJs16ZwNzFYSnzgw9VOfa7tW9v2E/nrVTnSbUhw
B0XaZciwT7bc+GFxYtfirioIY5s08GveiOHotloJOl7tseGJOMHV3rDzeBzRGfHr
jMTBVoHvWh+Gu0f0f1bymOnR2EU642UgVjKhBBxcpoRMwdn8AxcDGZIehJk7fONw
XedExeqU5oPKRQnYqcxdD3dci/hY0+g1qx1ZIZENqkVUCk5BdiuDrEL2uGD0/LBU
Bez8b8HP0SCuDRaEO9MqrfXBtQyKQZWyf3MVY9CjIPl+6X7b5Yb8u5Wcp1BYNiOF
af+3N87Kd2hujuL09T0ZYuDRqGZKXPEZHQevw5VDL72e/IFUB0FrPbMctdvZ22X1
PFmP+KYQTanl9KDlNs9A1HELZE/05CWCnkyPGdPo0+awUruKanIVlWT8HDx+UTif
xJrMBikMCqocI/LPZnPIEDbEaJphwRgURn/BVxWQb6BDPMavirXUuLhh0niBO7yZ
MiRZ+FjpB4/NXwyysYhZFuWnlsTpeA8pptddG47133rk6RZhUWYcW7Eflp06OH/y
mVItnWr2b25dV7eZCED67XDFlZe85hWVCm3gpyuXx0ThxamqhR3ZCe/JM8xicwDb
kggqzFw5JbZbRU+2oH+YD6P9xf0QQtjl99Ijj4Tm3V+rTWMuGO/c1k0HqI3WbXiC
Gn8OepiAP5raem747hXReIiyIbsBN0vaxvya/ZNlfZ4mZ39qI2KJC89Me6mKFo5B
y0Ts3BMS2C+8jPD3zZngmvubJSpq23tt2AeHBVaNfirjTVSbCbOGYVd/AnOcNTWG
iMP28PQJPwjj8GLcuJIjzTWu9VXcVgMRNzb9EZNFgPYqGH/tITnOMF3HgLEcuh8I
PmDmgMERGdy2KgSMV2GPxA4CrsTiOCKmB+oKDzpV9yKkwmPoHrYeXaGOoqgRDrKV
WoLXgpERvajAp07US/CGDNdlAmA28c18b6Ec7AbHK67tqjgBZZYMwuTCM9C/kmrT
8WngHRbSFLE94+LFtmpef4L9mCKOmRiMXq82n52dtEVzT0UPOOtGBQ6fWC1PF03L
y4nKyojsC+EfB59HTq1neP4PRJHXzIQvy6iDgZarqD/JFjkQOl7OVV6+UOma/T36
HRRHeGwvTP8r9J7L8dG5oO6va8z6uHXUatjp7H+HdJg4mKEFArJkXl7Ih3PZAv/Y
aTGZSvMxYcVxZsdYK3MCaFkAf+QOnkG8G1dC4v07AhmFvJZlMYINpizhcGLRfoms
5GbtDmXwgq1D3LiIzs9neiIGnaYci6LZgNNVakYgv4hB9+66RK4irULiqoC7Ywtv
PKFWvP8a0jMNcxNlVNi4xmBZKQv10cxw6uWmeZY2DaafdQC8vU9pcU6a9+5zJB6a
ohlZGMmArKGfMAUXEIMvXsPmP4AmSAGGKiqQPQ4EaKjuOmHQ1YKsfcEgOwFibZjh
SmDPJdjuLj6s68oQUyBjEQMHJLjWwVX9aceztwZ8lp4ViUAJNiAX8torkRSXCWhG
1QiUE7WZfasdtPWXk2cUYP7CpkHLZ1UH+y71eo2DhSyxrD/8gEOuS4ct8DUuhq7f
N6eVxc5SZObV0Dajz+qj4BZPKakls/IKWjwalMtxk9OVBwdXduKnHKjOqBqUCqpQ
o0bupIXfVzDtMr6kvpBmRMIFcjAUreXX6x4wOAPgfO1D7F5B67y7mGP6kM8qxOSb
r3Gpv+1sAj7VpC2TnuntXHMskAP4ZrLMlyYZtTUjU2lLzaq+98KGK9ad5GB4NWeS
MyAAmTaFKP+lBllqqePME9WaBUmMclCEsgyF3QRzOGdhCi1X0PpXgF3jBvRpKvPJ
EoZ7Qe6sgfiJdgfhq6Vc9aBFOxIQRznZnbwdbA3f2DayhZTGqDqZ6kQPIZ/piazy
ANOVJ494nkW6r4YdQYdYn7DufiTWtr8ldhkpWNraHBT6C3/DTNpXEj8ssVqdNc3F
0KPJTX5YFg7kofUn0z1G15jLqM6oWwrpMrX/Ysnvnysy1RFeeAxDaUDunch/zhQu
xcaja5yt2NVfXrvU0x7HzQHMqU/aPNZYs3nnA6yWBFpGuZrWHZdxHoDaHP0Q3XRW
oMLXScLfCba3Xh0hKzR+RSr52ADJKlmNV/kTN1Ux5sb0PV04RJq07Pbf8rm/HJOq
y5+fOp8ZEYHzUn/meeV7pVHctCRO+IwGyh5Teh3Gd2dEWxtVXW8fAd9zM/TAByhH
bay6iMkHcIn/JE2zVAqAQv9+1aBLpBM4QtgVGETQmhhkM01TRUaCReoejU/Z8G7Q
7c9GfcON62JFOBhFFTfPjX0CFORjz6pYx+ZsOVw75ghez32kPzZCAJlIoQKxnha7
DCaHpfFPecgdH6f55+4jpFzseFNhrZuvCLqWJ1J4WIiBpGcDBc642BJOH0wWl820
9iV0MsFVFfId8FcTLTAIVHbmguaV1vZgJXOVlKHcgEOioITHblYyiYUM0As9TFbL
C2pgK/NWlBfStxOZUjH0LEeQuKagZdeFK28bFIPLNuKAeeyPuDfPGNH1Ny/yrnUw
SVHk74gUnfHBKP85oEdvqzrB6SjuhHVA5zYqqBoODg8cWbzRDXaUVm/BG/JUCwB/
xOAvvElnwsziq3hpdMEpHJEiKCkSDaz1yAPfla5hWyb6de7p+8wTOpuKuwnvivvd
2a3YxlXBgPanUoPAsUgPHtS0s2RuDycL9IJp/EeF0okfaHUBiO8ZIPzo7b12PFl3
0bMWtU2wIislHhXLgxCLspheVXmWODLIq8Iy8dnq7MbhQNYuBS2Znf4kWtY51o60
9XDuOSO6olkADxXjcRzbsWsTZmyiCshJmn1i0t1RaOJBetYojvRBe43cxKQBH3Mt
nC+EbLx/ulQiAGNI3NQG3emvZLrbz99CEEAosa4eH0Mx8uVyfuSBmIVMe0cRPz5N
qkAWCFC1CZda7SxAsftFLMGpXcjxDVxiF6ATu+x6KyNXzcX5nX2BbCvKq1UkY/Pe
++B5pRL5R8hHCqa73DwYM1EyAPpIIWTCRfql00InGAAImK6hBmjyoZ8Dfr0WlvIE
AITcOcUBFe8OMYI+rVuhynHtoHEDezKgV6aTqPeCgQ9S0Xue04j7SqQmtdIIyUuc
cAG23i952YLQW140b7HxAkNraWZ8CkWpA7WwTDEYs2MXnmvbnkpJweI5JuY64V7+
57D8POtygUtzz9VeUIxmQdfM+CFTIosJEPmkw7RgHk/MRGZPmbdy1qTmmAsKQ8QY
Xg72/3/mke+tU+o3xtGrlatR11P+S2qhYiKu57Vv7XvFL3WdcIiWLC7iiZd5Avls
wGLCaPewDAHBGCdvgPG5bAkpvHbso06B0AlPVnSnSLhVQ4cMl05bxYDJL7/8Urts
acVG+45slkfPxk6bzadXQ8d9AsaLn0LpVIjX1cwGkVLSePaiZp8WllzIbD3G8Dra
EQVB+L7StBZ9aAEwYxSMAe5+RX7hV85arY+Bani4qVomvrOz32zrnaal26zVN7Pr
xmgoVhtsn54NEJRxG9sFGAYEvSjs630a1RtEMUokAABRrjxdshn6RxAZTARMnNMs
ujApqS59b8INjEB+DW6Y6JkYkeWYYwj+Ktrog2lYHtDUo198BBWL2L56mfY5Sldk
MrRkX5Kj9bNqjBkIyeyMNE3YAikF6iTR0I9d8r7N8nCIWfWBauMUP+zSF6D9/CSa
GMmmMgoIk4ldVcvtNN+PswtJzHokqYfNizzwf3ZhEjxwzqusDzB/evmGIW3arMKM
QBfLhbI3qULh4kc87qBa74//QDXR357fG6S2lnJ8XfuJe+/QYeEpe5Y+JRwks3Hn
XNCYUMqRQiDXWItPzVZtXRWxuWZeZZwwAx8VYBNHF7weF053CgbfyvM/WHs9qhzF
odKD5sQ6uHNp+A96TTlOeP7FbaTPtjH1YVWogafxTkvmZS8tDZm+EU+E4GymSqI8
RH2Vp++h9KNjnxb9p9pPZNVis2FiwbLI1uaqmyFpNXUa4Z115pr5+zKCalU3mkvK
0BDLDM3z0Jlq0gPKvwQKkJUZGDDGQ4cPimC5QN38yCo3VfpMF3YiQXztPBOKjb+p
ayoJ3+f4DmtdQtqeh/z6hxEkotue285y3eIP4frrYuMoE0nSoZudnyNH3TrS2S8Q
TmjLtOMXmhxVCC4hrX8zU+ZBT0faj5+VnQOHB+WGvNtQ4psrFZPP857jff/fv19v
artxpIw2dUe+Leu8hXOCWB8JJOqjFigR08RTsyDrsxQ34iEDFASF4E2/sgRWeyw8
/uQ/mZk2sLFNWTEvCuPG6nVgMXk8bQfTVHjtDbbsK63WnIkmM3FOtHs4rjy1jZkn
D2UgqEdwKj2PkVQNsWNWWmbIez7RlaFD+Rw5f18oeNwlueCgBXdLr6Yjmfix6/9E
8vIA5TOJ5oJ0iXeRTkJSnDJ3aLoIhrTNsoGhkPSjpbRNQCuItuJ8AfSCrkM3lUSU
DjYbYU7Iv0iZ+s44DS+z7XmS+oM1ZkF+i/7oB7Fdn1OHgZ1F+7z9/H0jQ2JVlJdN
dAQ8GxBtw14F5o67BVDFQDjKjvB8pJazwBER3ZbmMYaQXFZtpU9igEBC4cXqLx03
yW66PMx8SKa9jGYmLpEqpKUxM6Q0UcNncDXo2DvOJ4lQbFPhEeu0svZd2IjXLjGA
RCnyShGTpSx8D1ezkRPji7i2gx4WyyGAXF/Ezho/gtCkjdWaoDha4BdzTvlT54OE
HPHJmPM/TEDYtFeQn3Hp2cJwwWGm+gj/8hqBRVZVK+CAAiwnAisqaoDBPXXQZSh2
Ti1XowixLL4ZrxOQzA5Ocws1SN5No/Koqgh/taj6ShEnkSR+iuGmlDGbbq3g9tU7
p+mPxL9nMaDN8dRwV9fSAndLvBpRqHtt8yMKxmXP3xX9bHRuA9a926EYYcuqeGLC
JbWEgEaIsoi7d3tSf0/hu5hGYx7H21JWyRoLEWGT5Thyj7HF8quXpRQ7KMsKe/8z
jKqNL2bKijUSVffu9c8HncSWh5H11rfQA7oSIpylmn/UoOhEwnOE01q5PudWULGm
3w5Ej+mFAo0SuSeT76PNpdv0oG9PialZsA/iKiMsb3uPlGU+zzwH2gAUpzQt7uGt
pZfH/rUbQSe3jjfR/XLC8KQbkewn4dxxfhtJaOXv8oCTOhmPYoZeuY1pfeW/Ykzj
JhcFKXbtN+hHHcDHUU6OZoNWr3Ns0VAiWiRrcK/BY7fDaAEHJET8Apik1H7bB0wf
oS8TbxNZNj+miWJnXZMTVCfoC+X/eVZ/1COXmSHhrEwTuYkAp2TL0til0duWVcqb
l2nI1ElBcb08BPpoOH7DzFZXU/HaA6C0iCOw8Zifb0P9TA+CrBBXqG3ztdoRSABb
tE+efuWKcgVWcuITAwQJw69GgKHv5fIifm9S2yRZGvAEcN6Nb0G7UlS3O42F37j/
D2VwzBiUBUqZ3oqB2maaOEgyS7BqbSapM5dDq5prAhEvL4TA4Oa5GSSXB4YpbSqA
NP//VA3GpQfe2QvFdJDT0r4jCtAhJw0qb/hTnIQCy/75RCHIeBO+jBArtgf7viKc
ATEaZP5W9CzTjYkcPr1CzkZKnwo9v4YgOsFsFfOd3DQ4u4YnEozVFn1xeHJKXwf5
SzCBKjhYjLXcsy0Yv8/7W1+4bc4EE07p0cx74AVULRBslHNCw9BaW7LHo21FNTVv
XtTmN/NioqlqVAwwlVSDPXZ4P0/Ht6eSyyoHcA0LLDRiL41VT/rghsCw0M9dgB93
qNRkLsgP6tovPI4HdbDLpOEQc1o0NlV2pUzOIVTvYjOP1NebGcsTeU6kbPqhOwzg
7FDV62lQSPz/D7I7gNlluzMJrEeHW7Iy5q8U0pbhSgdT0czifsiYwns2nDGoW3He
UqCSmieiKYECMuLT7XutvmvCBqlCskOdTD5FqhhH/syN09xKsgT5UHF98m/rHF34
xehNPCzlvan0xINehyZyJ5XPRUxzxthaJF2P/Xn9sUSNEK2Q5P3C7tbOJh6go9Ie
7F5Jna2afCYzpGuY6aWgubhqJKyBpRDKrgVj7fdwDOn5uRV6xwXVolhDcRn/8xvG
pDvhcYckiBRBkX34qPWNqk2wd32mCHHW+volzEBke9qwtB3dXgkw55TmOhNPbfOQ
sf1djESXXHIr9A+lzZqLmxPXdwtcwWatjS2z7/XfbCVEkbSaU4zLHQZ++FnrAHlK
91VQga0pNgjAPweabqYmBSM0hZO9CuedxevqMvIC7UZP306tR0/qm9dBHHK50ug+
o4TAuWZpbj8sBdGwIoJ8lJu4pNZZpRPo71qG9nLzU4xqhB9BFD4XJB8rLO4JxkUd
matZTC4dbbFr9EfhY41kiMS9NBhLGaQg00yQ+ZKdQDM2ULXM86hCboEkporFoQT8
Y36hVWwncA4m5xkOv5d7jjWh2hbdG916Crc0triDBA6FxHDJL1sfpJ/ZIR1+tEIp
B/Xbzq1X0GFMaaAEnkUEJUUKMvfPLqF+IrlXUR+17OZl7HYbWEI8tA9BjkSAkycY
5rS4BFZl7qiF2BGhAzuHWdqTWFp8gTuwABb//BPfIDF6rJBpW9FKG3+JA6dF4Sey
sJhTADD7nKcQAdSSbyrFX1v+X8LFJtTviJVXUBQQpVsclaSrHu5Vz99vmKXQkYP7
hhnr8YaAVBQDfcB9nFEGdgqiLtaYuLbZS1DW1yjD72ZzB5mQvY88+y9D4SUglhQD
NQ7ZoWLeS86nXgSBReThzC/Pb+hIzPdk3+HaKe791f2RvQGSBSeYiL3rrN+dkj/g
ioQ9FIrliW2yCuqsNHLnfxY5jz4TWoNm41IW9S+zKHELeSH89vinCMrR+iLizLyB
YKjHobSSPT1ZPNHBY0u8IMgMhKZNCyp26XaoY0oU5dmdwOAliXbqNHYRU4xAueu+
Ha472pmLGrkLP73cBHb1vzbnL+NHoE4I09RoYCJ/vk/NODcDYoIfR/ERtnnG44j8
pC5hjUuIHdSuiR7tUu13n9dLR5O5bzmjm91TlWR1fFaXubSiOm8WmcxnXirljxpF
DtBTJf9CB3P5yJydxDaNMdEEJcp/umBrfD1Z9S2BvrNw0o4g/AFg3BYA20Eo+6PH
PJlAaZp6xniNThE+9n/vc1f6pBjrA7RpKkO5a/k8M5esXUXWcBmVS/SQBD/evsyU
mtovMLhzrq+0obzxRPauE+ZokFHJguA53FJwBKv5XFB0ub8pD1PDfCktvr2XBomj
bip0FSEiE23mz766DDBcu4MsbhOcML7vtsxnZfkk6Z21sr/WRU1vzQSjJVU0/wy6
bHKnotyL8sMW0NErx5jxKr38iS32UUSl5w021mW8Aes51by5yt/sM+r0eYmHdYtT
O/6lm9OWnVruT/9VmgnQwy0zbCTRprjS8/miPogNxAJbu8/obXzF6W2fqz736Lqr
hR/LhTxFm/zw+TKJiQrQkEzAdxyWn48ozvJXZ1u+LZ1sWC8z72e4wPwxV2/qwRSh
R7IPjd7TE8RQh7CgMlTPARtQKiAiqwokEGzyDRdq49BT/SyuBJbIkDjZMq/3B3Kc
DgO5BXMtEw0G8HK8lKS6cnp/uqTAczuH3HX98MhOOsAH8gzdPw02Oip2k+Z8Xfzc
bGha7as47kCwuIp+jtJfFvqA5auDAjxOGig+0K5SYVYiP4xVlxVrvyoHMLK5FPJj
ME3nH3Rt5E9Vv1qgWsGnj3w/cJPzsF1FzRPZkFyszFovT4uAS1+SfszcR8Yd6gxY
WxBaM7vuly6kRBZDbW+tYiu9w/e+xylhyNMzGeDvHPn14Ra0P4Kki+WyR+UJ8Ynk
fc3X4AdQM3f7Yjp0CWhuhZSi0HBihm1Qd8GcD4FuKjKyRAWOgPoXEENZ5JA3ryRJ
IUAi63OkzdTvOgibLAUU5rnQBcoGhfEFJMhrx+I1YUGLBpHpORfHsVkQFXc6T82E
nr7DiKrS+6M6WQWXc9YnWEfJiFVgHjwXpXOy6iKFQTIy5JI5ewusnjFTB7BANspA
espmD9TmDrgVg8PPZpZcdS5ICTD665RUoYKAOWC56vmgiYsF1CURhAyels80oMgg
HHljLUHyHt0pX/Og8JdqgG7qYNtteISnyilpil2a3Tq1fzD47pe4AzZ3PImuKPb5
6P9hhFg7yCukt86961fWUyx//OxRWf7uzUSMQG/lmoBPsn0ONuyTB0tkD5Dy1M7R
7W68tpi+FA9c+qnaM0GzQ2LaE3D9SSyLGSVEnvjjxulxYqfJTvDdV1SXNjorEGBX
5Xtr4leGM01toaRMcOPyQ5DKVISLCmtBr39f3xPbpRUASIaR0ykemoTzhI9nt6pw
Of8RH9QeQq9eoVsl+maa+kxd78NPjdcVLmvjudlDghmzMf+xqnZUj5dL7lIVD2q0
difkWsR4JaXyKGAy9OT1xkZ8wdQqJ1jq/Yf42aeM+Ygl1YR5uzUewSloDvOLB5ht
aypZjFJ+obOK6SzSK6KMqvDdQKIyDknIPhGTAZA+LNF1BZdbT/5tHoz3n/UWZnF8
3POkH5WOlpM1u2wpEbuG47ZyWA7YSJVttuCukYDTVL3NN9sTV6dL0IIFTFXHIAgj
TGo0ye3FCjxkhanItZZdzm2dlk6fjm9byIh2gWVFxuU1zx4xV1UDHzpIJ9G+bYGv
cOnk+REwfjiV2yi/NGSCzhf8/i+ikQoaT0zgKyqjWoEpgHp8JSxwlC2W3OGg6RE6
EGDDmNwaJvPatFUPTngIoipdvGp17nLzLnBowTTjJoaZPtXfA4HZxr5WIbiPCmbk
WmDfvouO/n+rstD1Xu3c6kMLYnirJCeX0d3t5n85XBqdSAbRAOv/Z14g/XsvvjCF
FFNTwlPg3QVaW0DDBcdp75x1B76u1T1vE92n5+NIgChuCsgrrhKyaQedF59nvg5r
Ks/Mv+oSGj/ggPRd35iFpXRgs3ILFjcE6W4j2GfRuxv72OWquYlc40pYYzlrLTDm
Ooq9Muqc/iFosp2JQ9eHLX4whIl5pMFCXJj+xw2Wot62m9Ttw7BFMHju6c5+WeTd
Oeka5N5GOpg3Fo2C3etj272vhlZ5dtenJzF5w4JSGKn7Jw/oYL71239i+pTtG+0Q
Hy8tMNxgXnBVWlFSOdzWZkE2z6yZSqVuSS+yR/k0ekRD16KHcabBUcvurlfSJxMu
1ArOBvluQBs/JOZGlEJBa/pR8kjOfCZl2juRnM72fYXC/Mb8rbp6B2v3YDKd73Nw
WCFHloupZ4VCFmbFd7RZcWxChcmX5SCKcW1DPw4aqKbQSPwNJTbGekYJUS9Q5Fi7
7aWkaIeJQUN7U4enimSKgbZo05PxrUKasmSUZXM3dPIycAzA13q3jDSN0+1WjuNm
2sTEcjwDJx8s/Pym7Fq/4Z54GJhUrZbligAGZzYBhyJbDOn3O7+kORa0gpJH2DYM
YH/JSaXe9eLhScIpyO2RhaySUztY39/1RTd8TVVMtHAfqBJGRTxF/gnJTVpykFCY
Sp+57HbYm78wEyVSrIKoJDhB4NouvPh0+r5/jFUvfT1F7fkSUZQlOTA4vjUR3cJS
niEXpHDaUwobj9OXMNtyObYZqdHvNbNhD3Ykn/8rTDH+0j1bw1re7HnyzG4eFenW
eJx4+UBXf4zdZri8fe+xHE7tZVcxX44ps1Xs3To3sKV1IwZhNrDy4YPG8Vpt9VvG
To16KmP7PT8oxGRbgurUKNuGIyMDwlMGcUwf2Dncr781ZsPtnncmvzQWivUkgUp6
cYYhWPjJSumiftC2fXC25Oy6RiaIfGpjfUHf/1OhmhbEvGp9D71tDgvKD8MDF1n+
D6MFYKpIOMMpPw8K1+novS/BLDxbN84GD/KcfHyltIf2G+RixMaS9zfHcaFaIl5V
W5RNcQSTC85L7xrKUR7uedRAvuR+bHISgV/T1keeVrnZNsxuRadCFtJ6bmOY7gBp
yNo2YEBMJ7w36IGIJvWb2jc/L6ZFYqspOTOIJabX1tstjXTz3xOdIKzgHgqSGd7E
qiSmUXN2uurHGCQUYaWgyc19R1IgrCPu3ZHrtuWyEnGkRsjZ5b1wgxYlIT5dybnu
w91TiPRLRS1+BW02LJhOBnbZ9lKlE6cD/bJpgx6qCWhcc4J6VefC3jcYhM7ZzeKa
5WBlWmnGSVxwn73IiOoNlxU2u966Cmw1eWInFZovbFoc9Vzpsx1y9WYLZMvB7cQ9
68QTBGaNYqFPupmZhb34tnboROvja6e1qZx+WxLz8WEx5emK4MopsBBdnra7bShV
F/eLFo3zpywQK+1wJXS2kKTg+3L9qiNNhqjSxMCvZb39MKIrWLXThFyY/uEz6LW7
gNWH4epfzm1axXJ8PNvcD5dF9Qnqef45R+6hDvABOToN4IphbIDXBrK6vdxzpNr1
ZCr6+//gAzu6uUVyNsdY1nic31cMleol+BxVhaeXvFW2MnzZVgu4xgc52Dy4AUg1
rq3/RTxQ7tnOCmxlXdl8LlNOqpyOZ/p+3nzEiQGEhK+j5Gp7YLnXNxR9MbR/g2au
rmM3zcwKikMPgOhL3iA2NmXfaYTOlfDaAWlOuGF0EWjLWJhAsfKwR1bbHhBFMZ2p
SoX4dwUOLNewqGvAkLpOuXJCquHvPE4ZTl0BpsO47ND7ABnxlrZIcwyoN/UMaXnX
Yj66TV2GYhLzhqMwu2YglPXJHotJebf+USe4RgGG8n6qnUIj5rz0/EfnAGBDP3zL
T0j38EXVgWfbkW7sAir0dX44gw4h5JK89yAqooHlmpntimIQRCv6PKzcSGiS0iau
8fYZ3Y3uhLpIQN6r9BOXoDCjXDg7ElWJdst4MjurwwE+a42Fk8ZDTFHTvYklMK4z
kGayasdTNYKoR2QTO9ooMDf3fhKh/y0RFV5sF1L9rvPapb7Y9o0RMe/bpd1zZeEq
2qQS3AWSlpiCZmCf/apAk4NrvPlueH7l/l3k+gFNvZ60lVuQ71Aq740olCq6z1XF
4qb3ofaIH0x9bDIr06AC3rFhTKDft9bM1pH/2DwM/mZcnvuHRXBJHG4nCkPdRsOp
f5F8a7MHDn17SFr2NGI7uCbPu4jY0Lhooj5o98Bu8VmyMBeC7+sRxeotg81YYDsC
zGb/FaAMtN1FF9cI8ulQJKBd70JbhJxoHN+4EbCBTkLn/7ET36KPeAIaNO79V4tQ
iXOUERpCstbmq6zmnvFoVC60+4ufK8q9wIw/vTpG2GliuDv2QdvlExzNHd2oY0df
f0WoMN7uNzNko7cm/EV/ZDjP7t5MDAyxyM3alnUSkNReloQLezUt6DxiR7ffUF4z
6aRTSw2H+bRqnNKCuIbl8ealLZj5/nw/2FNH5XqyBpSoLyrWN5w2U3rmLZFU9UaJ
abhvkAAeY52dIQDrZpoOt4GVAPVLexuTg3eahVoz0afH9jCf4wlEZIhHftqlWj5R
QnhnkhPDmfE0iiinqCZRcsyZBh2gdM6xmqIlsYBUFOEiDy3WvqptByEF6g55esx8
a+AZNdJ8IMfdv60VOoecVTpinezsQ0nNynIzfh6kP1KFdTD14NPBOqoJUfccR8GY
9yC1j80CqojUQdA4wib1yskMdbgK3uuHa8aKUKgtu1lm/Cx1QyUQx0cRWQUNrIqy
A8ZlnTuWeXPiY7eoC+2zM8ySVnAY6fUfl07iv3wzVmTu7W5c64Chl1g/X1iFz7Ez
bUtCKlZHahoCtQnnktRPKOzcuycGNBWT+X5eKRNwBagD3cQ+XQJNM0+Vx/m2E27t
YPMXl8xKrRx+gTlz0mRVPhzU5X2uzxr2meeIJcbl8bzYqS5WNt0yumU+aVo5tX4V
6YZVPLAMgZEeTJnyF4T8nmUBXw4T/uBCT2aAuF00Kyx2V1v0M+e6u4G+3auw7v+I
+BKf6UkkqQPXkZmEtK6p0XdOxSQnGcC/WtS3fLPy5SPjcS+CkBXwCx4RMNdhfSFK
IOpfEqu/3gqgdWIRwaZbh5HfvC2R/DNVlUF9LE/B4VR6l/Ls47q8kwUEEmafifKZ
1CGyEj6Ua2CDbYx7GY7RJRhjxFUAMzt6muvtmejWjvH7ZZkybaoSzw8y9Bhl/u4p
nLaqlzurF9xvKfniFp18YLPZeDepJG48owANuXKZpV+nB1QXzNNWn+OWTwtayJAY
yetAQhgB4aLCia0WW5iK6WY8TW1VgYGLQm+gpcd3dMCxXhDdXIAY2qmP9JZQlZGO
986A53NDEvsCivd+LThyD7zUjh1zCjiLyfvPIfhFZdvNsKEPFoYi+WIGlVepuoVx
hsMbizZMj4RxXqjataldxzwHsKF8FlX/hudPHFlvJWI567naGztpX1Olj8Qu6Cma
UbA+fKwABPhIl25jD/rsESUcQew9dzdPrqPOA1ltAelNOXXaSe+OCYyIvnjQ+y6P
pf+LLFjz8ATPNSzxyxLromVCJl/bvL+M7maK+khVQLOsay/33cyEM0hfGo6QOknI
b1+MAW6D/5St1SkXx2POlWRNmILa1TsrF1TvvLxOcDzBPja2tvCOajJbfKAowpZt
1ZQeaMZitT52m+HoxTKaEuWB/aO5C9aZIdxaDII1SaIJULgURVtkA6vrDJ9OuYiZ
PyCwo4jJ/HtSJ2AmuC8H8zbwH3vGCNRtRTCsdTwrn82WG7lVjAsImziisiLNFW3X
sETHgMl/Y3N/pvy4lP3bZSFsP3dS5IqolXTEWaxTrC/bsmQEqtBm+BpZxdbSJ7tf
pzFXkkH4AK3cM6pcql8r7FcEhWLDkGL+JCaF5OOkwM7db0/VZwnDIVkDO1RehL0r
KdmPjUqE6YOoThOL0K3U93znq2G4GC9Sh5LfcDgAED0jgZV0ga5OdqElqgDtAre5
+1OmKHdI4UGLwFu0GJ+7GUEQVuDYdzg4vfsKzRl1Q3VA0119jWojDhOLu9QK0tLY
RPs9mdTDLcZZRR2zZxPvPTcnDNmQMoZyVzBP6S6Rzui6RxPC8wl8eDqdB68CSgvM
MqwoFrlSI6gFH9fXdYeCHGr2nXjC1D5ddCzliMHI5O3TFRLbc1RrpB/+B9VZVJQd
Rls/3ibodaB/Ejwh0YTEOuVeuGX/9JLiN54bU9O/uAtC3zsslFj6KMIyhTBYdYGM
KzWhpWb4xRiWwQSQW+SnuXvPOItKyOPs1SoYwUIFkwUMDPKZTWKNZP/LvRic2y4y
EXF9ipt23sddevIEX6k4pVyPS0X7Rj0deonwwg4iVIRmCTp6EE3ezPGwHkmF4DZ7
JL+XS6n1oea874uuzhsuZ4G9qHmF5BzfUTWESSkkAnkA+ZEzwPnuFswoDJy7Rn8Q
SkTrnTFxMzMERDcnRKjs3X5ut1jv2hfPrhfxPgT6xdZU5X4rEOXG+CiZM5x6DVZU
mRo2yH8RnCOiTA3HN5338R04kNyghROohgxzYezkXCunmos3x0Rjt3y6eyrGZXFK
UpznTT+xjFOLnfIbRblj9e/905drcYHto6CcevH4vaF+zZL4G2yKTfOpfdOdsgkg
C68jTpvXo/amEAsMioCJprY+lYukzo+zkLFpHXv7HRa2lGpU0jDB2uapw1JKRXfZ
Ix2EcbRvLUIxjYJCYAV5wJt3JYzIU1LaFFuSDj/wXq4LxoSfQPMVqqFWQ8p91l+y
5VCN4DGSnjoqb4dBNDIy5cS2QygtR9hiUSxgJu6B0OijtrQABS+2/dGdYbU2wxHk
60jZ5s6mi1M6jmSeNUjdRcxqGmmoCHIAXAoCsFiHyPvKVV+RBdg5IWB0HuDf127y
AcI0E6rl+pt2VGmuINUXmtjyBAkj1Aj1siXSTnFdKzeDWlIHCki4xHQSC0/LBHCo
O6rp1keo1GWy5q7DTGrnSki/ATni65jMMTR9cq3RcJS+x1LT2qk6pWan8o10Z1GO
zHnCHvyYM0a4RhWQelKsIA8F4UmlwiAqfIwgRoQMp0B0yilJHDfehyt9HrMMydMz
k4QGzE6wsmjxFwSGCcwmizvaNtdT3zacz53HP+cpco/0lOnAYdYUYYMw5Ho4XsEK
mguzq0oHsqT0ut0SUCdgG5D9DqHZxamCAapas9i1DmdeRb3qCsKsftGhQeaYe/vW
ys/wkbVntvypRLIvF/Udh7GwXWySZdsNNHCFPGrIy4orh3RQLGv3TheEgjg/hYvZ
39x+UknILWShNd8s+aeUT/GAedXgQpdAU8BlgGitjK6LP1o/xBAiL1cCx7XDD+Ea
6kGY9jO/N40udWuvZsXKuzeqeV6wEsoPgJuDzMpscZZFEldV9fM6IAk4QGBdXBSk
KrEv/FeMtJ8//RN5ztoR8dS0eLbMvgZ6QSvrPC9+EbZgxXKTluwDxhrUASUHQp+N
9Vp83Ookj+7ntRx5PdVx29JyYFln7tkcT4R618wIcJ3b3qdhew7lO97ZWHzIQusc
8kSx+3D3ZiQpMgRKqfrIx8d/n1Ia0LmW4P2LRNgL6sBF3ws7qORn5pEWL7Avzz/6
lwRU+EdIj23pvhx21xEjyUpFZZL/r2r4lbgqENnWx40Q8SseQr0EI9PC6xZGvqp0
nLnhIIR7IkJ1YOIOzVsDzQxrVpSfzRprlmiFdx5KcqiYKd6CxkffknObkOctFrtf
l9CoaMxTyIZMLk1UXsbNurikiikcd3vhiniX+16BNUi4F0Gw31CNuu4A1NNXyiy6
n7774Erdxbn5VBvxI6B4dcLv+LvSlnZkZ+NgR8PRMQpzS52Ppbh1dvyKQp+rPQrF
9F2mlBnF9n7bYy5cUAmoHED9/HUQOUbumY4kFCaeQd8ap6t8JIiYicElSccopUY2
e+Sxim2Cy69vdm84JbcZYg9zg32XhXuoEit3XzorjAQZE9V00YLGjN92bowyqdgq
R0JM+8T8ey0/EsTFbNkI5n9I13CI8NJJFM4uTAGPPCM1PQEChHHk2WyH4DGqlI0Q
1RmDcv3MVOV1bmt0JqL+ZmEr5K2GfXtptYcqJSadeezGq8aRwzp4fqN9U0IYHm8O
LWGXpb8rVwbj2YBfHDeUv0Zo1QqVOxJlJHZ9MqGghUp/jIPr4ZirnkVezjj7Z1AL
xUu/snCziY1Od9QkMUuske+kuyLHa5rzBtkP8CEhCJnJ8DMbLuA/hLi70RL8FEwe
Oxge8qH34Ducrpz3/uKGDDMmH8lvvVZrnLbvJBn+xFzlXn/WeOCVH671DkTJVn0/
lyKfIYgkriGOmrf8lZi6j2C/TYQ7MyeqTVTP2qVdIMiraFxrtyP3hp9HLqhLyxW1
8KCDCcjWzngw/PeD67zLyXQmfnt8xATnJDGhE90a26NBS77pdb7ehNGccfzO+ufN
SFIhzlq2P4DmTRUO52OAJHaeSK3HprQ+7fCGSBCk2hUg7P0krWTKGYJjJArKtzyC
8zfTOlgnkiamoMlmt2AE0zVi+QwidlzwjexbSaBgSWegxsT5SkIWnyZGBjM6CcVT
6dZT0BZiZpj8aoRGlez2YFGM5JJ/B0yYMDhEYX7U5kP2u5JHqVB6glWVVsICsPKE
VLMkdpRX+Qa1OPKUiAKK7HQYWsr3npBZi9KhrFyy8+2jyl+/iXbLdurAw5/Nmu8c
rnYdVsQ1ZbTKGFk+QcGCbMrheJ44UeEc3aZXUJ87uUTwrAcYShkX6AYp2hqDazvt
2ReA1m4feI4Zl7TG0W4C+OXVUKKzzDd/MCq+espktcmoL//79vnvGmxfFUT22eW7
WdlkHFx1OIhvtjv30ZJmTufvDBH77x65mnuq46msPvXjIlNP9phPgaJYgAp8rify
4q/F2OuI6meGDENlDH7EtltA4pSmfqV6gFbzDiJzn4JX3LC3qx7I/8m35EW7eZSQ
AkYNsuPTgZgVdVCf1TXXCsR/P6373kGxGSD+QrrT2wLiQlVzczw4QTwUGNRr6Rqz
Xbbl6kAsN8bH17WbaSOXundwMHQfZgDayZSfAhXeRtuzc/TwBFYcxZrvAf11aG+3
u3/00Wx0eC2l6rYx5DxDvUlGdAT7RqNKnasnObKG5eU+i+8JUCp+NwVEdFeV2FFr
9RhcPUub5WU8Wn13diT4D78H60ZoDk+aoyAZxc61IvDGhXZD97p2+lVWj0+Pl0C+
wDxZQVjU4vrZabogfg75t0FMHLc/ypP4MIM/JkcfWhMILqWKcvo/CT05hkIlU8jM
Sre7bZEyBFOQ2Le4yETshidJ/IkWeTigleSkxXDvma7HZMbDvDdXQWYqvBsOdA3j
eKMUVe/8Tir3udfAO8bvxqHerfFUWLspwvOR8A3kFQNukU00N1H3JVMrv33XDAwp
vveudtTEO7GSuc7ZJjhK4Npinzop0XZdmmHt/SA8iUmGnSHkINdwkhWAOgnpu6p4
2n36+PLnSEC3XVEPovyFD4TujaynzI3wMtUNOnUA4JjgLoFzhfKsVroMLmA4Wl7x
xI6quQ/SLO2CdQ2/54+B+Kz/j82heb++9FYMxPqNVBopFxNUSKfXVMpNy9+QhxI/
uvSldXeQxOX0DjNmADqRcmZz3kmPpkffwdGoTywA9sECrVSaIFsRFZqcq1TcciO8
L8IjCM+swLjCupY9KhdHwZio5BIy/Y5Lr2Q1MPw50Cr1GPtl2LSr0CrW+H/kkZtF
GFZPtlonTWp5JhbGRrIAYya/jqPDlHE4+96S5lz8R+wWzx0xzz08uhA7R9KMzcnS
lFH+AWNpyBQBTlr3TgpIqm0fMxkkVihY+JVPJfhpfLmjQ8WQP4q49PDX0C7RwFnF
djs8QLms+az/vn2kou6fdBb7zDIJ+uF0OR+khnCah4EDri0Z/dP0sbqnf3VB4Pl1
xR4y3kqfnq1mlVK0+zNO+ro3g/g2nYKPVdG+SGSCwx7OInVyFGDgh4yu8Mpv43q6
yWcg0x5DcmIiGFXXPilAymD383qq7O/xddCQPgr1eWUAHTa5KCiBfwySrl3rtslg
zhNXSmosNac5QKwAaxWPXZRjFEznT8mSMk95OW5wjO9hYgU8ykiAzb8/6XKzX5hS
wiE/F7WwlDCGWJsxsgq0RjOTngTPebD0gWdbuFKoFfVhM27mAea85D/kaMAQ3Wd4
Z7w36i9aqVtFF5f6JJ45puCShCqbqrmDxMX5IMCt/EAMfnqwtvfUikS+Ap8rW7sH
Lt2tltlvpFu6d/le4yKz5kCvMpVe2MXMzMPbabfULAtPqqLEO8DdeqN9l/3y3dW9
ePRYLQpi/GK3orFo+RLobHcZa/oRBd+WZ/E+ZAc0L+jkL9ViW/svxww9c3AfJL5D
rEZkimmWicp1SxgEaoT1EJvs0ysZdOk2AmK0Hf/m4FutRHDNYvWXYkIZ3DEEHIiF
Ip1iLdllcVbkVFzJj7e0Zm4A3ZzJk0O6v9dc2KTM2EVT4QaNeDLM4eQjOjJeNslf
cVRSTSWQbSOUKrWETZtIp7S1Gybn/5GXjULWld6gCELVvwGKX8oIi0SoJF1//E+H
IztTRpltg5vajwsRJLxcVgLYh3yLavJMjTNqPUW3XNm8hNM1g3g6n4mL88D9njbP
5nBbHeUTntoIf9OCCRCWHD1cSQkvHOiE1YUeGqCjM6SO/SlkHquE9JbeivUMCSOB
b26QvzNVRIL8N9pB80c8/3BeJcemzG8GvicJtU1wps2U+SljPuGlRq7KHRgJZGaO
YeMD3AYWFPjZ+y9vSb1NkKabGHFFxLk7soyCaaeNQMlo4SpvkqdFeG0T5r8JxJSG
ZS3GbfhzR/Ptn0yW3ZSBgIYRoKJul77XF58x3FqhMRpIoAXBUv926F7J6l7hloVC
Ilqy7B/by0Wa2BOUaa/2IROR9UO0SdM/0u/6Q3W6W+W67m2cgE7Ckwu8wFuRpoyl
PHuuL6MObCjFgJFwTb29LN8usqH+JdvYuWBgpwUeqE5EpCM8Rq4o/grY/44VBHjl
zpGEO47zlFYPPFP1GSYbz1iLp2d7vqZmJmu3S5p2WQq43qE2MCmXtsZppEC/TYyJ
A6cRRKYtn7LvSl6pkJjkRzFHA6h3yWom9/YiaZMqHc8Nud1AD4tA2TBWmFFC30Am
5bBXn19JdxbMq4x+Ty6VU3/C5xEGwYLbFl7z8R1+OTMax4qwuHeRLDCl3pmbWeuu
gS3cM5a4DJePe6qbk+p4RsNzLjLSB3EoR7rWH+q5lYSEHykl3EbaKAWAmJIB25dW
F1cqwEujP2oGe3l/JuI6EdJWwhCiWweBmRFm/uRNK8p1f7q9BeH1pkq/spzA1g+b
/26N5401OlPfQOCPx3J7rBOMWiQ+AeVlWidznXjhLUzQ91Ws/QJfykg6CdBiFlJy
Pd9OjN4vO53RLbS2vFQrAJUykgiGsju7NEWxIbiQIqBPfkh1js0E57GSJ4hROarr
GfRN2exz78DidyPrR3it4s41l2601FG8qJw+sR2D1qJVb+hTWYvi0nPx7QQOP0l5
kn24aUKVsOBMBn88krhMXWfE7LTRpJSuL4ehxrisU1KlmAT6o6LNsnMQCKRsVXCa
J6zLz0rY4gnSqja+3A+9D0Lfac2fhmcrBF5cBuRc9XWmZEHX12JDh7g5dYzw1shH
85z4R4hUdrPb/xHAEwtKJpRkvTaLCwqxQU+eqEYV+glTrUSrdaIqwazVOhJreTIT
rODSd8TgIuKaeuCwmuoQZGN1IBJzeyruPbeNZbT3RcxuQxkr6ZkHzW+KzSZ7bjGS
heXVvowEKsRSWsPXlkIWAlbunwHd2pHMK0OByoKiwyIuf7IT+YixzRdeG2xViU20
2Pd7dSlhF1NShHJefAQ/TfzRjMcFUMbkNfip26rBM+ByeDxzDgNjjfBjK/FUAVP6
c1FLvpk7W5aUaH/vxjPxI367SWK5EMJkrp2yJRhuFT6Hn9iv9npTVnkrhfx6FhQB
Xs4WFo5JOd8K769kEdGTkwdLFCgNif/8j/vqBIKKqngr7L3/I6i10701ShXX1UaF
NHTuH6eyTMbNI+Rzc/ReM8/afZUtWWeiCisZLwjg4dTBYrm93+Iwds0nysW86pzV
GE3ocaQjiwcRgl32mK68ek5nWKwEgrY94IUiMzB21gQ0BWay6TPWC5tzIzvtOazA
JuvU+O3QKf+b/yR6NyOea12FFUWg+L9jfhZaj0lpxYEpQLOgAP471Rsy8wZyp/aX
ppP0337dfZvlEw3rbXtRnFaNT7tjs2708O31aFIJ/6CIw2HLUY80vSonRdL5GqND
O7GH2VJZNzH3YlE0KHOZphRKKwTRuiJFnjR545/BDtPiZB01Nqg3EdAvY4s/uCta
HfbRdy8weKGWPiLLY5HROjzT6z8FGO48VFlsuGCnbK1yvzjBTfVUVaUJM6XReyV/
BsvC5xJZgkKzo41bfPgJNNihzDyo8Q9m2iZpdDWvAlDjqA3EDtq12W+rPD+N09a0
ABGUv2gJMSu/CWcibMNvg+mvACXBdwWuWXtLapXV4ivbGPJGJ3ge/U+LD9SGgQIT
OLZTaD7OPLhr8moqi4W/sHvUcNwcXxnRnWwiGXyuzgPahevXHMusyUQseaj6Btmi
675AVKioeawDGZ4DrwyLAmsZt3ZBavBM0FMa65MRRznZJqq5yW/t3CZu8DyYR3TN
pPXYPGw+qunBbTaDtn0HJ8L/PGoqBUqw+SsGS0esKo6iqKxJay8bW7mqlVH7z3yk
peW55yLqMrGvLoKJilr22gc0oUEgYDmqBoU6Sa4iJVJ1f8NNRcRuf9hpz/Tjg5Mv
dpcSyj6chqjfEMmSpx9U1T9vvhdgf4i793rELKtT2rXxKPt+7r2yYdp47H54dd2E
j8jzwvX210qHgHiTzC4s96/zQTs/LPbIO30m2joreDftE1/PAcbyjmXCUJjKZZj4
pPDYXcU4BaKk4oybAAxCtRcYYurw3S9dKkjtOIKW9B8zBO0wXtmdjVFTp4mrzZ52
08QMQ+1Z2t4v+um2C73fKJ9xzXYMyODGWZ4DKtznesZzimeAqJBSNoY8P4vRo+oH
VUD8rWiZBe+fUggCgfE7ilrANKknP3Mv7K/Z/MErBBQWwYi6CkVV/sXshmittkYw
ds+SU3v8y+hwDhqqDJP98TvpxdnvAGgV7hDr5Fv4Lfgudp9OZs6toZ0sSn33iKgd
fUAalH/l2ZkZTvOZYUrANPUTab4ovB9jZS3E7P5kzyMtSHN5p+FhOTlNcxy/Buo5
IAGyWaFCdLw8w7EcoSjevlPYev2PE19IaLDuDcCuwNITMybmWxhypRLywk+jpw6+
VErwJv0X6+AL5aDEB5PA2xt0IWUCSgQgG8srsvoVF8Zh9/GacqtF7VcOYVeG0fcc
N+ABECrFmeTwg+WmrhaKTHpWAjPLj8RIxMwSKbmc/r77aGP2jStBzzIBcppzCpZt
xIll9l1CECjjMEYy+0ap2o+638lWsFaCrVjFqzUVDX3qrKgB62V1k4aKAzBAC/eC
ScSARvzCsvz4A71tvVnyNIf37/bwhaOE3SCj8eTGB+PR1Lg/Q+qGGGK2lZIrzcz4
8qS9DW5D7gIkLA1Su6M3+zb7FNFrrJeHr+efkJPq0dBnIhTdCt98bIgrUGwW+Iuq
QHJvy9Ts9x05qs9IOU22oU+rnxoC+U7kycFp1yhps/hJrtNoaD10NqUr+1VSVT0i
Q9IHUbMFQ5dKn8NVSEoRFA6igrUjuCvtmabCyklZifAnY1zbVNqNH17aa+WkbWjm
qX4XRkB10Kdmk0PjLNEM7gb92SU5rGJx/zctacB2e79NkFaRcf0vWdiVBMFCYm5R
i96zRBxlampN07m69CKLK6Er43dXZ5aVhumt+vuSro3VuP1at75Yl8/h/Ta4Pzan
txCLOpFPrXNBnl/NJTU8droAcR0zM2C0Z2bxEEypudD+of2bU65Y36p9B0G1M+cv
8JZT6XObxY104JS8uVDv+1RiujXApQfdS33ZLVjcFdq961U857itsV3IjwVkR7Om
mCzo6v29yKww1HUoCDdfgOq2mkk+PN2xfQZKmvdfyEBSt4l1JQ7JtuKg8b/MpUit
wSwE6S1mQhdSSIElvpU25NJH/JiNYkYS4XmXbLb5szAquP/xLknWbYK+L+pezqZ2
sLOaOdXbl6GrSViFdssmEVhERu6u4+ajbWAdDmJcjAtQ3EAASz0fRe3NFOQGfZG8
oeelS0O+Rw0yxtowAKqaUSU6BVbTXOiWZDGJkLrZbGenRoIKO0jjyEEO8O8LcwF0
a7B7uGjHG4PaRkQC+EPzPQOHc9dndqjuEolrGNiegvqTi0FX5g6mIGP5w3aiQp43
l5iY6/Geuf7O6RJk5QPogwlllP7016topaK6vJBJ80O/lWCXyxl48zao3UZBSDC8
J8umEXxcr/nA3iMOu2fWT8+lOfPGN/BkrYlZbpJV7/mMPeuGCX3CZw3xCfatm/Xk
peGNwQeJTbLYnsF6T5S84apgEeE1dnmtzfdZCyzCixzgGnkuOdDq9uZSacX9cyx2
MBvUi1t89IzFPh0Tg+/bPzmlPKxdedvfdY8UCqxg4NuYMMaHH460M2rw+fB80tOI
yQ745dB4bUh3cClWl8NF9EZsYmQdUCsM0VVJ8TRdvls3h3RY8x5JvxmAqA2VD4ed
pg5KgxJE6M3+3mgY79iP8EKfHdiK6jvP/l1EFbDeKko7tqM8QLqwQkdj8+3Z63rQ
+ixD+MW6iT12EmMCgmjSBQkTJ4IzNJjUFNmpVXRaDniDZZFQOmDYqUsSa5uiUO2z
vXzxOAmosr+a58m3hrjfOBchCap2zG/LL8YkmjHecA25bDYeBbAJskTSKcyBnkoX
YE1hYBYxrY8yrIb3u6RBmCL6wo2rmoAm2bJm3djBqxt1oBWEi8uriNuGRIqYOSRz
HbNUh99dSHEnCFjG84U3aCflcy9EkQPNUsyLga/xdnJIvBQULw5KnrYSW6+K3jav
dlpgblyfTiKdtxnH5C5EoPoawyVUYbTDB0ch20i+RmKWEuOVGncneoqYoqGADncr
OX4THT7S1FVhgYpn2I5K8fN/p5cm7EOP+bFlw9Ejcojcjtt5j7hyT+pUSBPmwPJc
RW1xyGrOQQ3gti8e09Xakqmx3fZevwduCLbkAdxuyK9/K5PzxkUXXp3dwWNDg4e5
BxpV6pUTRntaE/V2+tM78jxby8m3GALSV3uIsptDe8bwIdfN0DabRcEXh8N5j/XR
lKzj4nVdt1X1vkvsmv2Iwt9z5IRWCmdBIoKg1wzd/xbghep/j3ZQaZewEZpkxUEV
AYvJpywQjrB6NxolpEYoPoeq3JUl9MjVYBeO9FwDS3gfy7CHSzhAPVrT6bQzHQdc
yxuuzMjXf9oj+sJx0PtDuTiQj5ZLFH0pg9RZ32Bsv2eUpOxfpr79+tEpDwuGPrVd
mTZgF9qLc7NzUppXy3z8tx7jUuUVcvY/xbJWNRN8HpnUOWW9z2CzOicMcGCZpTrB
ckbDpd71NXiaEjJ3OCYUF2v05eks4zcngbFHzPRerkEQpKClQN4WX5x5Itjcaxj2
teksN+4Qm4EuzII3O5ZW3kxnTgZ4+aq5YwosfU/HYuNyyNu7onxQVcoPXoW9nByY
5pnvWBnaO3O4iGWSEFNi2RMGvJmU1fZjG0hd/Lbx6sltAl8i2erqsMl22pDfBSFQ
C53zCCaVXThrdjtEJHqF3Pzgx/Kvm1ekFYzfNFeuNbtmgxyXuce4j4tmRMoJKBU6
3hW4dNNVbigGOICF3pXCIQ3NgzoqBxPedl7DIY+rZoUFHhKOknNdU3bUfi70hF3d
GbWqbffzOb1/qWpB1+Nl2nPbZXOidGbOqSR7osWXCEsK3aVpl236zlZ2Q1Oi/ciz
4CXv4kOsO94s4YfsSGwDbKiPQRG+dfKXD6fFNIcNbcmAZ1un2sSeZAQcF+HBQ04S
Uy85iWG+JmLuXvT758+J/hYOOoIUIJIQjOQWsC6SdTArV+gjLR2Xr1gZWPjDO7Yy
WoalT560MgjH9uF0+kvJgJr13DLS4waikWh/8+7RWuggabhdMFXZOyw8ADcTnHD5
OvhRd5+5VEsBHqHbsD3R+hgz1u6nNO7CjoHc9bA5V6VO2rzMJM/VHktlHMU/HWDo
5GrWZggGklso+jmREZN9FaLefEdFkTC9A+//tUiul5JbsoE960OmHeVxtJ109bP9
HnQGQpfxh4yP7q29+QkXNIZMr7ZGlou8gr5r8zjYZhqYI5pMrenNg9cTw1ldeJfP
SD3paiGvaG78tDu03mjnBbdMpOL50zNVOZQdjS7Jtu/jrjlxRvPfyTTiAnV1aPN9
l3AT+ylXdGGp77AJvsoiEs/rdt2OOBqHvU931PiQ5Dg3Oz09nDmNxpvnphyVsWFR
umDvL9kg/thN8EvfKodbCiS0PfDy/2Fb4Yr5IMVENhUkJOPmRCTM+TDAREpr1XNf
hcm3dDjD9dX8ffOF0xGYVLf2Q6PlzTA9MvfEXLWDWG4y1hBhO3HjvLhdmW6qDb6I
sq9LwXqggNrFPEZ8jzQOupN7bHlbHj0sKPZKLLtzuNOsZj7VBBzB34bwEdwqJQb7
9hXyyw2bWMrLXgxUphXwhV8eefh3kwW27EQoAFtJR3iJ6v1mb4PsW5ikwqGI87UV
GzxgxOrs5Ebf2tPYfwoQR3CtLUQB1vrxptExFlMdzWdcKrAVCl5qxGhk3+Yk7d4F
FkXDRwRgmpbP6TG+NzSiJP3gdu6jfdHYNhWlCh60D86jiHagg6ziqYvtoxG+s4M4
KnZeAAO8vQ7Na1bkz3SAaxusgMuw8Fb8cjtRzbVpkMXA4jgEnhWU1nZyKTroRLer
+heNjVXAbmfehelTocutCfSnEHs/wxJhji2S3SV4+HKu4RWOhdQrolpnN2hVciB/
FGPirRAOvTSIoES0/5CwA3qnWv4u0eWlJBIMJ471Mh5dqVBeNHWI2zKyQclHrLzn
Xbdf00N6EUDFaLYAOaGbA9Gk2JQXpLIUhU1nQBqgvDovLWS3BAxEjwLirX0xo/pE
zpwdzDe7VQAKAAOY/xNMMwjqu4FT/UOVKjWKp3FIhiAkqZZkpURnl2V1xTt63yvw
u9Off+Kvx7Fc8TZzFmgMcbHkM8pjGipd3SSGak+nuYHyMCDlzNBHzpaifdA8BTeO
Kie2Yjby6/c8PEqkYGXKscHCqmtroiXK6Ak5rUfaQnx7lWTJju0WmQa4TMB6FgNk
EAE2J8pLwfgg81w24FBPHVjljwI1glVyZ72296iB/IJOfVz5BcTD/NY5uE8CQvpV
z6ui/lMWeEvxJMjfXqnHSL81lzYxDfxPe2cOeIyPS1WWcoKy42uDxX6193pYUYR1
lBboMj33wdKeDGeYmO82v45TP+bcZ+HFCUHOxsJE3RgVnWPJp0QfTvF760NOWkDF
UhY51uWQcSb/goNGHZu5vI6hg8SDAuPOsUtDSRFI5VxnJBhaf9yHBVruDWJ96kCZ
Rwa8wOD7S1FjGU9VA0MviFFMTvIMrEnGyOIuDD1H5npVju+IGWcuHE+w5b+fYaJz
4lNuYJ6uciz4SrvTSzauCWIoAhMJLBxoGvFTGMePa74DNQX4BMCHtf2evg3Ba3+T
PCIo0a+sXQK8clvtaX2pa6JtKt/onMixI4vt/adlQfNx5y2VAVs5dy4tw+b1R9Kg
sF7ETVqtNMWgarIsyHrZJL9w0DtJd18MuKUrBf7KTtOKC+ohWPDD0IJskZgnyywl
O76QjQwYn8Nm44uPyS8HbAEQ8PzFIWrnk+mWWYpB8S/Y3tjvXUXo98gq08GR7C7q
25i4V7ExUITE9ouKGsx4T7w1puUpn70jNwxOoFcx1+j9m57V6+OMhrUU0n4soZ6c
YyjL0UQcddEXT4tfJuO4x7Eaep0sXui8EtkU3dO5npCIboLBx+dAn0JaDRavdxr2
WxWv30BMJeH78gyrT9gOGBzmJn4esDXJ/ZOkU1SHtv2qK6i/MDlW7oxoSsxRyvu2
B2orCSXBgK4EDULBKTNzUGdp4WmXkTiUKIemQl7YXxorq3sPcW9Zan9Vs6qSmpsG
t41RCpn6pp/r0FtWgdJydnvZt8ZXarmiChq9zVy7FFqK+OFXbrD9JLAZPyBDTXOZ
ZtbfVbrMJhUKAhNNQJZXqjfChbNR/6nfYFypdBxaAWtHy2qkABMmTjkZw56Kk9A3
6FwtJxxII46uIaBkqRIw2oQhsDH5PvGBAMX8OuZM7gtYGiuvbRfpDxwLRPJMszyt
JD8TFlBLj+GpytHmvwQRn8GFz5Y4x0YPLNXdyrXcy7AaeTaWaBioRgINSpNJ3+uY
cY0ozYvSUg6Vq221XrCDJKpldUzA15eOKmgjAsbNfaxsNN2Y2MmkcubsqyN5ZI7Q
HJz4/RbVzX1PVp5razPytcbx4W5PfvkQUb5grBTbeNE4MhlFlJrM/SwepnrzhMLL
nh3h3hdxAy3IuOwFgJSuC32mZUxTXFtyKasVir+jBbT+YAsTC1ZdumW9z32ilXcp
BrkQqc7j44FdwW3xqQsyFrr7/16NWgsxauxCFPRagjXpct2m0qjQy6l7JLNw/DtB
D5qvaAF8mnYne9cByoWHeEImsserZXJwOmOC778S2zhNHcJHv2YkD5bflHFM1wpy
6KoKxtATpqONBun+3jnliyhACVO9m7KdhfDBI0jDdMlYSEiZyL39BYDF6h+V0chh
iBMgs4qOKIokWdtvLBxEz8wDbu46OJWRhaWadyfkuwpuFdgdm0ezIi0tM2L1INiO
0XDR5dOHCNh0eMEusWlBJrkZDGPHMCFUzHGJTBghtBg3BKusyq6Czjy8IFIru/g3
e8zaj3iE6PNgUzENdcRj7q3bZlX3uwO96BzqqL2Ww9/mgcSQJyQhI5nDOIluUkCB
EI3cs+/LeUi3UXnirmopnl44t0asvDl9/U9RV4FIKPNRhd32YbvwS0myBUZ6qQ/6
s2k0Ksico/UuT8Jd9Qw0k/FTKrqj0cSzdqbCQrGkj6eaNdd3ta3l1+htJM4AIGvK
XPIFQJhg8vFKB5Ut4aixl0CRp6Ylr1CbpKzz5OyKgWNEUu4C5VC9uV6hpVmDh4Sh
kV2C4duirbRgzumKkz9uejjb4Irx6HY5uf+G9++0xrraBYlt3+JxKiBHsgdOd5Uj
i6CbdaaaubaxdKVA/FnsLCex5UOlyp+OV6pYdpoqzR9UWcFxD/5ICRHIczXblr58
Y7VliLK/Kxf0jm+XDzEmo7zQSowe5sjLGWQU1MpA/mdLccxSEGNBNvNmp978qvHV
fwB4SSWrXmmHpVrjho42d3JZBSnhTQ/xpfb8caxIZGz+irLEvPnpgeze6wk+KfOL
swo21HrGndX/wlpROrrZuynUkQB3waAas7tST3oTBiAwAvBsexrnjvMOlfnlF9tg
C/mlHl6x31/TRQNNH9cGUqs7M8qC/mzpinzMTfEalBDUshQF/u+6RiEgwpteNcUp
5CB2TbeDFOhZYV1I+j53oZB6lEKXPoZJOgkXHI5lcE71BrN/DTIVHjz7huK3hU5m
/ZlehBB/+zUO6tiHs6LQXMUVF0HbMRmRSDTDZMfxkZEfHZPrkb+XEihmced6pVoP
i5XgV9wySpFt15G74nGRm9leUcsx+vaWL6NLEi/95dRhxwzqtV6Jc+Ecb4qdOP0Z
pf8nwEv2IwXvl6TL4OuIZvzh9/FvwyYugtHpOILo66IgfWztTLA57EUrAZsT+znG
Sqj3+aQe4bYzjBP29xn1UfVAxyRYZ68gDSIrpoJicZ2+rHgJp2nQiZDF/st2cg3B
G0COEiet/sxlwUuMCiEtlH1ZDl8dLWMmhTSeS/3JY4+flK+qJFCXtGXdEFtsm7C5
yBSDWGR1+n+s2V1hJ6RhDzFTv2CrD/kYl4SLpKo0Ysj12MvCF1aMWvkPtnDYEcQB
eJCAS+aTyRghlB6iGQq5vFM8DY6J3daQLwIa1z1x5FzXLQ62TNxWJcHo4V/ZePft
5OUq+HTiylAmiCddCKRyCXV4GaNOIjsXxSH7FGg6lbJ+kXHRmTiqpYYrq+74bsc3
iRui09vq0c2vnvioX8xy8Av8LWyXRgeu5YjONEXVb2vzzTPShyg9TgvkIST9taci
o7zXKQKh5UY9B+bXllH2W5FI49Olr2oheb6DtfguuCGpe+YBjNOUHhR6de3qvtE/
U2L/aVGslLX2CAzLj7FhYY29aZ2Sw2YV8mocVNSbXErU8TBHMsFusLXrj0j8wJr7
Vic6JLG5PH+ZvX4OXso7vI5ZtSMgrgqvfrHLb+NlrTKKwjM0cmN9ckc1d4FLp+7X
tKxWTD9vIgOvkHfZPcAHBSiNNl8nfimEkhry0/OSUWUZb/W7Ze5Rc+fSItUwGL2C
7uwcBEW0T/XPxEr9W+4LKdUv0XZR5lI8S+29u8F0rWf0wvFV6nLsiNqTvY3+EeZQ
N+rw0bmMIkJCwhgunwxiUwYiv2kWrwTJUNkeY0ZYeJle1OPC+EJpK2DXb3+uHHM7
hA9zxoMUsAxuU6VFFAV0V0fV+M850go0rcr4/YKmIvcsUw0Gig0FCP+K9CbaDYwh
KNTPuiJBWgmzFXFpfoo7zjEQwT/6aobMMsG9MF6t3G43T48AnmJ5FsCfOYeiz2A3
voLqIeFKfW3SRbQ6A/Oyd7vnw75Wo8T8xv2dbjvOM/O2c0jw17u1XWte+hRKIJkN
rqVnne99RTaH3/O0OMsUyk9cJWgJ5cGNYX8JDKnvmghlXYl2hdEm2ZtiBOe9eR8I
Wc+FvL/OgbW3yIbUwIHSWWdTjWj0D7ZH7LPO8exZf0tRXJheBZ86kQrYmlXv4WzO
0QkgLqsmVkhm+OoZzlveWEvTzNzU/J0oW/5VvhGp4lli8YTwg8kR5/TTDfBcNt8W
3VIsIZZN62Z++vWVKxEu2x8eac4cdkuog4bHeIw6b3+VRF9ynddEqSRKDBVlQZz8
PN8TgO+6J1ID1epFNcLk0dfK46g53G38tYXj1qianiRQd4IhZrQqPhvyiWNjxCcr
eoUWWftTPVqO1JI8Muqg1740Otd5hHS/+qnZeAzH/rDUm4PpKR0u0U8NYZsb6iF3
Wj/Qm612Pc+UPqUpyAcRByAC9k5ipycFqr2sq+c0aJU+SBx9kMUVZZBOjhLGVkC/
LSmjeJMFwKWtJzLlsUfotHVogI2v8L+LqwGwpUprulNXl/zuwb8blFdYVNI4SXvU
hr/nBBmL5sHaVqUdAPjFm14JjrP/C1YdxysNTolZc3b/JbjD9vGoSpDgd4iitij0
oahKquYAzWSP35Gv06zlmYWYA++Ch7HfmASkPvgcGR99G1BsS/Qm7HwAFYaA8VyY
LgDBocdrrXMSY1gEU9+pK7EJ6a4AH0DtS0lSDcMP3FlSi+TOBs0D615JXUCKvsns
TxG2BDED1omAvm4QhoyzHiLIfj0dQIeADjuzmWwpZHmqS4mMEJRXeP6Uo4wtTHAM
P/y25OfDXRC/29NdIIrHr+U6CNjrbjBhJtlmZIGBZfySiINC3pRVkERaKfzp9j+W
+UxjznxeAgSoriaqIRT74h75HPTCjCarcotqfo9CZ3PqujQstvbn7ASobQDViYba
WLeqk/P5etcfGekZN8sB/BlUWPORxRwob5Ll10tixKLi8p64ajNVBjl0kxu5j6QW
rXs8fCwLxyCzxEiMwHNxoTwpqt4f5gaPvAFygq5/WRDLb/QGWpQCpcfFKAnXV7Hc
A1S/vlr0NdpIe5cUa1/nCABruGSuAy9PM290thM4M8q+Sqga8zlcCzXgpvc0EaQo
dWC8oMUHWbOeit1tQMKxXgfekFIwwspL0TjI11SkG+xRMnhKsKHN9EczybMaF762
cl+beT0zNI+CmX8+YrtBCgqMbjgxo2mT68rLiUFDrHNhxB9PJIrTXboQSnjLMWGm
LQwusUgAqxwv1Rf95EJLfRUAcrVxuLhh8QymDizF6zpnb+Q62aG5Rstr0gy8NM0l
GCsMYIScqADmkDkULppgwFhRrZ5cQAwKsPAYbeNyIuxRi+sRqO9vGbTzqIa1k8En
2vIjraDjxrXcocc9cKBFU7dfd5gMv67KU3Ax8hotg8zyHuyO3GKmPqAO59RZJjdk
3Qg0WoOm/r/RaJsSOV4lYhuhkqymPeQQWMA+CaL4eLqrZCQIkbpVlPOPJPlajpFy
kaokVEzEFfIHyzDsVviMrqFWIpbOQeZULZ2e2ByOqPUFhQ4ZVIuwMollN5yu2EQa
aYhs7scNkIKqY3GUdBT/51j4kI5nA/5i2p67/vN4X6hWchIORgZ91aVTysipAYhX
v/+zKO4KMtIjvScvh/9G7lfVVa6xQBG6ap4Jkkx9rBhwzWT1iojgR1t3QFP5sSMP
WMk0WJObeuefnq3ccY+ps3hwUtPYQ60mgKjE6PwovKrmJV9Ok77oz8evKqbfo/AJ
BK/PR8lJeVQ61ACF0VqwqxJm1KBQzqhTMSdGnhdf9VG3qPwcGGwdTzCxZo6LvT/z
5X9OKhOYd6jlzLeoRYwNyQyyvVf4XyA+UsZjO7ICxxwgOYLaaL4X31+tl16Rk6L4
osfoTaWkLjTSzrXWT+IWKwzvAz1NrQNrDdIq9THrNNH7EyDkshJWzPiHz4hzO/Vp
S6VIdL/WsEc8L3eyV75d7mO5PNI4VBJtTPUFiaYLqlTdMt5tEyC9yqKT2YDsell+
RK9sX41itxEp6hs0qaWVHFiQgBz2chehrUHCqHI9UP5Em9QUaRtLQ+vKb3U2WU5i
eTuWf+gthMVduNXpP8RvcF+O2bWFZPnU9Bq6UtqaKwOekDvbrdeypatSsZgjJMpJ
1TO5I3oOxfmyhgdJgFXjHlZFsODXu5depmBmL+zfyzrIwW1YL+JZjTkqyGyCC7cY
HvcFdN5CGYSeNV6W22OsrI4Ejtp51743lN7sJNPQliiO1GgfktW7keiZPXy0EbBL
8P3UaoOSj+ysPeEbx8Ts6/raskXtTXBOo75kM9MQLpNwu21kPsSlSa5zt3DYDqDf
WnqV/GQsmdER/PQNvCVLmZwY855z6xL/04ovg8m9ryEDoVJCKmk9w0DPi5G/0eNL
hMN1hB6Egw60bn7fXJ5vko0MZgxQ2jENeQ19xcunaCRGcMxb4+EUPmi3SSgudAoz
5JjVcKD3WIHOy1vCebIakAZs1Btm19G4xkeI5vbUYudK1dRDAcIC0nFZAO1yQN1X
8i5/Uakrmgv/a84YMAzmCgr3g7PvDOiSy3VQySGwFXwyzmZnxHW0TSfe8+BJ2rKa
yokeLN2UboXUG2uUBhAWDgzfB35DPzoncVMtAf2EDipcoKwlRBPxbIg3vjqPLvd3
6OXRau+mch1prEzf3DpoCRuEhcwu+lVnvyEFNntDGGWPRUlOleu/p2rDcwPQkswH
iWoavh0U9T9JQMVS/hrUWjf+hDs31Kjj651ee7WjBKiknGZNAT72KcJD4xVMz4fm
4iRTW+SYt1OtIEhHKDrvw5yD02Rq4oySz/Qad+QdhQRw6baU92kQ7gxgbLznh6zu
vOnBZ4539zb1+AsDhhurSS8RsLhYvHT72zy3XmQbKDGDwLwrmK9SfcjWrCGElMx7
DfY6aFUPkEDGbGCghblIOlv9y0DRg+03WvuI+4pneLLAVW0VRjNP0Aw5tJoOSQHR
rQ+19Cq8f9YXrTaVF2blLljmLhAD8uMbZdRahZyIEObMHK+67yONTUOQPJjRd5B8
k45oH/Y7Pv5KkaI4/9t+gEYTAG2k1mT81EqOVkRybt6w3f12UMMmqVJA9di7nRCx
B09zzyyNRC4Vqrl7JKfn01SHOL6blVgqyCxKD/m+qQe8S5wNhXQFPIt/xSUKEC7x
AGOdB54KJ9jNRQBTE4laZCZNEECvY+iUwXycUfgJuqthz8ap5DXTYNf9vmZsSBmd
4RVazlFaO+N3+7mBB8vdgE6X85uAE12dTCVwMbPHEz8TqGx8S8rmBSP3kac0J0iw
FdnUbLHRNcgbcJ0MaiZBV+VeWw/V4cwzHtx0BDw3u4OdTQ0RoFKKSTGzoT7p6P23
8IP5KcJf9TotUwDVzo9mZB05BbAFolvPUedAHXlIDNvd5COQpzOfEponSQPrvvsB
Ed6ByIXxgL+dukhK+n9ur/K+27KHK24bvVn8yW7mi5Q6R816P0KbBzBPwVczSgRR
MgnSnZt21omufNy40f7HBuMCBFlSDqQkBeGtt3g+bWHDroeusTi4FP98jzKs2gaz
L+QtGxbx3tu5qJR0Vzw80BHhgURTJXYUQe4/9et060UudigrxhRgk8tOa4nrhRx/
aTWzuNtUSD28NlrLNrNltmIKDELzaeROpabRdUgC/Tsl6HlprE2pvI5Dh56CSitJ
D20FhDzEWLp3sI6xqRkPD2yBMwH8O1h8C79a2PtukN9KtFPSdv7HHC4aIur0zlO5
6+HfOUbWd1OrHjtFjP7OSjxzVqaEwAYQgBHvZ+J4oOQVI0BWD65nOM4o+8mjFOJz
L0hTlVdT5+rF2U5E2gB9AGOgnyTAzUI04FeEwX178HwtXf3EZkApTKa+6Z8nat+p
yScrOAEFzfehzgzg37Yzgb/YQhWUKXndOjXmuT77CNwUdKdvW2tVjbaawHVqBBJd
JiJS46dS/eykIEXYqaVY5ffDWCPJVl8rw0Ffc3X5k342oTSr6wYEL1qnrJBG777u
1UBm6pDHMkHVasjBLU9J7hR35yB9X8ZliSzTzKoajPzkl/vtPtBtxCTHauRgz/3B
S+lAzaXjJFo1e9+6e5saRmNojiNyQ545HeAoTUoirrSHbsqI7yEDxt/H1ZPEo3Nw
MvNSI6T5yIjQxBujsfuo8hjn8x3hBLtk0y5MfwHRrljx83ubvBfke3Lg4JcwmyjI
uJWCN8n5jjjmk21urDbBytsmVNftGzm7Ix+lFQzOcMu3f4uPMRLuRG1o6cxTsqsd
4PEodz7swH6/HYutaIjzYwExAsa82dS/5rYBfEBHCN6KzY67YYXP2V64NgKmp0+S
3dtGJ5qtjUZE0Om7x6X6N6ca28lS3TLW06bCYYqYi+MvTlyjumJoajFU40ePl7mR
Y4GhIvgZxciW2oiWJCP3aGPFEPMxRlADHJxnhSiBvxAhySfbdBJ24H2nXUekGyTG
tQQcSUf88tgJi8s2dHmVWRUYIQBVnP0LlX7qcSQRebQOY6fk4p/NHiFraE1APvlg
vp1wq/VTGVDtgPnChKPHdWx6c20zQdemXbyyXoOmZcapLkLxz3Xl1KWzZj48B073
kL9Y3QhMSVxMnM2+gCcwuuqB0LRKpEw9X6wH8+pIrIGkuuxYCF6YJmhRjGYEWBVi
NoouRhZT9MJHD77WDnMoIImf6OhBPK6+m416HxtOtYwYbGX/R32vZ27ciz8Ola5t
72Q/YVL5c1s7Yu4ogNvCuwkQa8/s0FHzZjvxMgL+vdieMIxpBZnOMIgMoIJtFhWh
tjYv1vwN/lJyXBhgkcp8oECdanK899Yg1kSfK0fFtPa1e267Bl/o0qg0EPFGSKoG
UhzmKVYCb9/2NuFV5kTdmFMv2ZwGg5wmuKe6PToDlyDWiTCEiRlDVju1Hyb+iVvd
GKWpkE7mMtt0Jr5rhTTcRxVVswITcRgpr4fcr1xi1Lf+QWIp1643IOkRayvxLeKV
muMAiWnGynthLxliV0LobNwyFgMBl+PcfRDp022NHEOpe03169iUbdEGNzFI+U1o
ifXwonpXQ+A6arToM8RnPUZ2sPB0S39EhORheIpuypFCdot1+TIugLz/stwZ7mPv
au+y9Ci/FCM1CCOZC5/lOd52FxkbsQVpxo+6EkJZigS1EEE1FkE1FQNy15NTVhLJ
xENSLUYYC2lE+Cn91anF5WBuyEpc/w/+cR9+M2X7rxFVHz1+8q8ZQ1DondrE2i48
F9aeactopuOY5MNwSoLY3uJkkzwaM6H9D9I6vPj4HlVyrb6MXvILyVGK6GmKFsgc
4MDBJ0m/HfSYkSL4ZIIfsoWZJaIMAeBj6BsI0hqKbxeNiQ6xAuNMCV0/Qd4M/tJJ
FROt6wz+HllFqB5pn3E4h6PAQBh6sEr9mKEK9uy+XcOplHhvkQ4XBZf9lLTwSMeW
x6ibCh9cHHUxYzSeS5sLPsXM437JOPE90jNrk8CvSzkAyrWa/HwIsmzSAuv3+Mfc
SulsDAJLnh4nqjl40Dyz8TESyL04JQ4Twnu6eLGq/6rKTaWvDAmytQpLFP4MhPpN
FZ06c/zqy3otyFiF5FiwTR1R5FBp/dM/BQ9amhYBDfvxuxObnmyevpRIGRjOEBJK
yNXDq+JKNjIKl//WyXVuLeAC8WjBLS3dPAngU/29ozhUjyuSt3jYQCCbuExcIPcl
OrjI1u1gFwbWzZU7DsE3nnKntwcvESP1sr5qANspToS/LiT2xqSr25Sl3F5B6eCJ
EdFKblmsRl92K3ASNpj7j2ye0UCSFg0SS6Kq5stQELvkgk537ak0i4jwZI84CliJ
Qq69I5zz1MAL2b882e0vcEqaQ9Zjv2vgsEA0aTHukrJz/L3s1kA0/FdXjLgmYsTB
pFLWF9DvY2dB/9SP+PX0R3MUPbHcjFkpRPPS+GPJSepHiT1mORWo0Eh2E3p2s1qh
FdKxFAaBw47TuEIKAYY4hIcr+uAFXBMw3Zy9Mhsjh3MvDtfMb8WWuxOEJBSQ5nPs
ytV56QpXow8kVzHiuBdrO3d+UxTVNb7naER8sy+LJ0zOflBd/8b4nvlYldZvf2IV
UHOjvXNp+gI3BnfkoBFK0ln/ZaaZpEvxufPUqFv+R/f0Qj/2XFwzUoQQF/n5Jh+K
428tCLDJG6qIWHelR4h0YbU6/+XZUUFaqRTGYKD9OzMdXQMwosfryr8JsDAb1d7x
vVhNpyM74KUs0cmZ94TRGOW4EiefYG/qz91olRgZejv6ieAsOcH+093slzJ2PiYJ
hcDhu8d1lx1p1x2baS63BQiFUOlnFmqUlTlyM9WoAiD4ZEBPWDLz2SVypEG95m3s
Jveg4YXvhLmI88T3UgT3rsxLQ84E6OHYdgRbeWisfd2dhoymomJ5KNG9yUtKqD3w
6sQ9SuIf2LYXhYhdh29TLRhOhE4v4l9Lpf5MU+2QW8j+Yq8RJEVNFVFH5aN5j0Tx
U4fzv0hALv0YGYm7O1j3Ze++eAnD/YYype4Qguj7NsiUMHaeHMA+MMQLsdSuKnls
p9jFT6b6qmBXjhm3Ow142j9nHDnlskgfhm6pzJeuZ/KKNx2V1jPX0yG/A+ZHR25V
wJsvbwFgjXNU7jJyMCB166sLlqmWw+dQjCD6xH+VVDtVuXtUfJD1KDYiDitC+hmj
NaxhajFSsrV5AappscWwzq+9AKlUE6D2kJwHDofDqtWmISWIjfmZGeNT7GT9KwAm
9CByBzYgUMtY178590Mxi5uP9ykBp/9+idA+I2z4bu8uqNPsSHOJ68jMX0ENm8t7
S/fw4kXIdMMgYZGeKuiJrqfeJkghCn1BbrX8StfoAxd8mtoZ0MdRq7bjCU39w71J
WID4+7fdi8yxwHIS4cnEP9STF5HCaijmyP1SUHPmrC9AjLnQTvQmE+NymUEaTwSD
mGZWfHZ5OQsAFVfH5L/3bhKRfBfnAY7dPSzgnmDkH2d2mX0bmZAIVUnAnuPtXu3l
yqEcgqBI+eMbCWsoso9qL6i8mXqpKtpPoMdhPv2sSTVbLE1f2KKnurcvf/Ph+Koj
3G+sBpQ5URQAjdslJ0Q3KLvzVznlqeJIUeHbNjRv54irexAuLU/WYPQ1Y9sBX/ll
UGb7g8KqwuoruH+5X1xoKy3CsXIQYfxsgX0FOh2Yl1QsPt88HnFbWNSeeXpTTPGn
AxkmOXPDl4v7RJckCKbbHW14MkIgfD3anO2Gp5FZKLJxSO6RYfHLa/tmZgs9GlyC
i7fO41iWkbslifhpkk3F8QYC+GH6Anj9zJHNdffQk9C+p/hHoLdEn+sypguwTjE2
P3lbmeCR5Oh5jl1mN7l+X9wXfa+ltbYvRmCtk0gbTAyMiyLbUNlP4SwoW80Hculn
b8Wg2/RmYl4NZw/oVoo3ZcFsc8xh5nEwZPB08K7qBkQZIAsZhPeUguyg93nI/Oo+
b8UGTbgAlF6V54JWfAJLwCf+1WZYhPmgIZL5/1fXRBZKAlo69oznG7Kkg6fbV0rx
D5CImC1cwIV89p7N4b8NW0bopypwcVUzlCnVIJPnoGUOLFL2FJHD60JpPUSpTtLG
NTHiPTb8+f/dE4EQAxElum47pWBIqLaORt4qzYA4btPb6hJtG/qaVmNtcKhhYGxw
xEmz+y7QDK3UFytVo/kA6rirLBsakDuYXPKUN+5fSOp3YhijvHVMsPb8zzjyT6Tb
/Yd/5OvB0V6vucNzaGbrcrMgRfjqueV4e1m2Egz9p5MdcYNUcz14+YJdldKAaKFp
iwX8z9M/KSsxlSqhdq20twmqHUJRnLVZ7rasRlG2kAvkTkmGq2n3Iky8d+aG0VVT
iThVYIjv9VZKuAQTyXxr9EX/wfvvSNxWMcUQvjwe3eD224FJWr0/7ZmrBA4dCI4i
wc24HEMz2LpvajMSqXrkDjgDynn1SPQe9n6Qt265hbAoCDcsi73GyxJy9I01ebtF
FmvMlOYeWGbGUS9OeFKWWto+jmQViS4aYPHrkSVjRCusNS7wh/Ua9RzGABLWA4IQ
j1kk4PzRzuvX581McR33ks+ft7xttSHnlyFndf0f14sT9QwJiLDs/+lKapmrRg5J
u403Y1/3Qjs1fxZdZi+SCM4xZjE5hxx6Xu5xq4yYQokajk/HSDzPP/ouhI2YOTsu
ecUjP9xyDMv5bLbrNzV5x08eApc74pA/KElB9MZgFw8XrDpn7znEwIYs/OgV++U0
IfaF7Vd63w9kibjnk77OEJclBzF1ghveNtoBMobxp2X8JZshn8q1zyFgqYy6uBxd
MQPrwqpXmBx16UTpqZTR/7UMLVNFqC65Zz9c2lHAMY/uvWH0RIQAOO+XaSYdUtC5
XH2osRW428FNhhaMcyiLvFqJFyAMPZrx/Q2d0FlBBPT45Dt/r0JHL4VYuz8YUjCY
Oxh4T1vfNsUklvxSsu64fR2PX6dh0QX8HpD11ifiiLZ5IFO1PaX+RDvOszMCpVcz
OZESQnK37nWPKnVVCTG50KaHrKm1iyUWyr+P62XmEXbUfCuO3DHXd0E+DLmx879e
SaDDUjqw3w7AgnIt7iL3UhbNyOMFySLah+h55JHmP6WSnWNfPEjbTSlJ+Yh6uSgw
T0gLVzLG4+K94M7wt1E2sMZSpYc0CHuxyceLA+2vMEMLGDDcKurPOIxIp7C8WkJo
Cb1iv5U76yAsF9F5+kybnBkGBGfuJc+wM9DgCsT3f9hT4hOoFrIAh2ZhmVI37yvG
PoJrIGw0lGxDNOLY2JZOOqavIkQRHypjwEw+7s1BEYikFX6l4S2y1quwz39pY02O
ZknApedOyS7QhF4ouFr5az/dmrFuUSpqBfFMacthzKxcCJA8ZKdh4pSLgw7Mgkxr
aJg4XCA9mVdhdGqBSy7UymomafMau/CIoqSR0sqGD1UaBpRkFae6Rw7K+YC/FHMN
hOMeVEjY/eGKhsteh4ku2Anl7ljdmQIRLGfg4CZjdtd6hOgSGvbUBmRHktHbRN21
dPxp0TqAo21JGh7zeQvKjwohIOwIQlWBTGcGlkYrVdDTrQsvx0idztkB6FMVGmkL
mvNlFD2YHr98XVpGv5hbB7WW6fNzVYcqOnrSic5QZQtHD13zqRXLdybvwjPAs3c8
i9TzQ5MmiBf/cZEAPX99u2EyW5wn5gUR+Tbh7ArGuBm1KrgtvS81q/9z0qXSFYXL
OgB4vvFleaLVyHxISZa+JzbUSyLUaklBO5x5S26oQ0f23I01kCQc6W2Q67bz7nl/
W1l52QS+sVclx14dojSCkNCpaRXYzdXLSdkOSr/OpZK0/H+1YPfn9G/Lisi24GJZ
p6YrHVCOv+jhbraBc5X0gjTOWSJtzG7QbNgysFexi3bS7cWss1dkWyLEfjA/ImS1
1fczMdTO49tLPWwozo2SKokwf6BLuDqBSKq6eR2wWTg5rmnqn1MGsrycWBZTZ2qZ
+ljXgun/QfTgyP+z7E6aMVt99sKyzeV0g7foh6NqyK7UftfTm7YRErG1D3bDrxwX
ZVuogV+SzBVV57et2/3FvhMo57lToN8IINHZ6/Q62OV7jitpDCKSv2djbdQgP+XS
1uHJ7B9/zd+WZDaNLw2LXbcJmP+rAoaomNMjrjF3+sr8mg48+j75F2qf5aWSpT+8
sNm0IlhYoT8Dd7VwFiHu4xZa9JWnAXfBmYE0KwpQ56q7F4tUc+Nvf8WblFh7wJAt
dxonimclNhQ45vRvIhw2/etm7A6cwX3HNYdwPdrzPMaNgY6Rj7S8XfcUqTlWE7Pv
O1j+G443WBfLNrSPiVHthqj86/sHCXif5dEgtNKZIgakGNJ6kSdOdau9LqEQAVQZ
kKXJR/h1DbqLsK/tWof+5nJq91CYun7oX6vTEUVyrcwhuXpEqQP/HqtBiuoXXs7w
KSFJkmpR/AVeC0Efp1qKrtsEvjcFXSw8QUWZp5j9ktwNtsj1I61G9KjtKsng5Uv0
A8aegRHTQ9hijT4h2WTRDWYgS+sygYG/AZcKRwnxeESz/cvhYrFGGtSkoJjpcytv
A7C88Y2KxxYIXVZJmXtY4LRx3JjcVqhm9Dhn5baaKQ/GpWxzh5yhpul+gY1Ex4IN
Af2c2e750MU3Bz4T7YQpxTPST1v+ZVQgQjHFmPvi8c8jv2bTG3S/Vjb1PMQXxkI3
XxhKrBqXFiXh3Rit1OXFAPVCeaMC9QAU/T701ESOBmyrSw0KjvsW5I1XwI2UO/LY
sC1miLpG4QDK22h6BiokgykgwwXLhM3YO9Af6UCDJz3f+Cplrd884FvAMNqk0JhG
vDKPTbY6anOdPefoOY7y/gtWrLzfp6reTMls0YJw/TYxeGyF9LnzN4mDeG+s+ZvW
/E5lMyR10v5pFOA0bxo1Wbi+tCnPreKCek7SwjOn79fZgeyML1UQdAS3mYUPTkKB
7eTyK3u5gClXpQTLpha/UoA8YyEENpb2UWlyeo44oQfCRq2nkUj4dkGyIXwAYCoL
y89oMaZuVbaS39sjRqaMovui0oj68h27XJZChg7NzaNCJxwdcVGEo15DYnNIT5Cz
HGRz3R/YPcbn3CZm5i1JvkupSSfdogPbFdGyuew01rFE0z6N5fCZoBsO/gR8syVa
GfHx7oR8OVUySDOU4wolkxteTVRrkeAJJz++mdGuP7pjXSpXdA5CJAfDqZ88iU03
/uwdMBr1vtTZVm0Z5LC3Tg8IfuJ0cTKQSe653zq/yBTVDrYV5kuLkWVKFXF71u9X
OONLOswujYX7XtYYXVLEBH9HJSLGe1pcoqA24MXEAjjqfKiSDXZY5ufrC+0WQvHi
RjQ+fw3lg4eZzmowXEDdTkfbfj2fZBXZBwPYqnlmbJMZsO5ok+pGgfvRSiY8bzTt
foNFm62cbjUes3ONgS8whsNZNU/cbV6jVDk6sIEK/xV1TCuAwzwA9cQL6ZFgCpFt
GQm6iBON+c0clulcPUP3NRsYt/LrZu+e1X9CHFAdNFDl/qfptkKx78RbatIl7KWH
jj0gU3H4V6W/I4Z2D8FuQh2xoZe7XpejKurK922W5Yu0KOY5ih0Lu06uuGc/+Zcw
vJcivdlJsTO6RavQH1z2Pi2DOCltyaukS296jDviekA8MavGuP/y+UecZHu8Exaf
/LgfcqbgAS+PzXdQ0ZyRYTAe+DsXxIcNaIG8vrHhBri52JJ0c6hhPe3KyhQ8tcKJ
hmam/1KbyeTL1Ud1r0ZZ1q/JwJjPwZiHSBt2Ts+1/cii0v3sZad5233fAC+qF52F
YqBq3uga/CyFIECccGxLcW0FpZ07rUuMneroSLlMVFlaeJOVVjCV+gsuc+3R42cw
S+NzepxFagCLw0fOJJBPu9EasBGu2p4igqy+P9haJzA9U747dCrDTBhx5emX0R35
a785TQaWpxY/LNOQC5DsQOjCKQj/bX5dcPZcgJUa7xUn3JAOapGHhK4sOVL313hp
6eNJB4yREOhVcxhHA8K97JysWB8XX0dZKwji0t8cujeaQswfxnkJoUP/8oe49mxp
hssei4lWvfUGhNeNopvTXeZaZypQWKOE0tGPhINyfvA6HBhIWmBbunk6oNCDmJxy
iztR0hK2KlPgLD6XcZE4T2lV70nYByGfTSJwtBPpZW68+lLNmvQp1GIaGckpVS/S
PbLDBxvJfb+se6XpY3VfWi5KwL3+mjdEalhT/y3mtqHOuiojR8p0uAL9s1mX9uF3
WDZQATSiKjhQxOeXk1YxrqeriAo4Baj/74N9abcE1zbEU/GhwJ8SKjU8TyCykKeh
AsKruDqJM09A7OgC5YORpQPt7ifBPlUukEFZsEdfUmlwAgws2fFFOdHSMwRFGq1R
K9f1xVPYNJlCFoHArr1QbXxvMUkw1AzGRwJfSw2NuwhOqtUBzJMQstrZhvjoNDbY
ps500ifm6jW3X77/STEi/hxuOK7rBxSvdJ1tKmOMfac83VIYfiaI763o30U9hg6K
MgplSgNnxJu1p0TZSMajsUMmyB/k9QznYecTrY8MGWy69ILkU01D8Jj7Seivyp94
gETASspF40X4BIScWhm8kLBrGyhGBVpjpsseCbxmGV18qkcQWbrfdGX39VI48cZv
MCyok6P+23aPjdTSLtPTplIfhAbfz2Q9XTBw6bRFUxGMxD9EArMAUQ9CV0RIojT1
1TweHdMUV0/azOA+IDSmK49r2ZaXaJs+1pLrlUKpW/NQSJYcONS7ODaa7x2IZ3mI
10sFbC1wLhoavtYaK9TGg/hFN/OqBZWvtEXOeYmumPIuJigM31uN/Ugr8PConrPP
t/h61wpZdZ2H951u6nSTyFid93UmZx1mMldMQZ3SpF7LwuGqfO9EKxDz9k03TQBl
BU/JwC0m0iY6X3PRa/YFZSpIYsbXZprmOnseyj9tswZpWGswBKlTtQ6ij09yKFLM
6SSj3QfVCQ7ioSYM6448t9RRb/ZVrruatyt8lyHaQsjw3nHBNZFeQ2/P5Uai/reR
PEE3qFKBChA9Or6sJknqQHpUetRUR0eFwub0gFsQiCrSMDNkNjKfVwIT7kTWKqiu
dWjCM42VIkby4NSFxHr/0fVTaLn0Be8Irj/wHBskf/sTwVLR2u+Qu4/3XtLea2Vj
FiL30L9PQeO87iNHJ22mISEHRU8XDmBkzqJ30WeAHmk6WpYXKrAnP6YUvSzpoevX
g5vmp0YfxWv97MaX8dk6r3C+9TgbkXaPM6jNf3CGTIFW9wqIk7a+VaxhN6Hx0fMD
ptjwqFlQjCqyaXUyXFm5+DTrJGzodDrvSbsq8IMMq550Dif1WrP6G9OysekMILCO
p0o2h03eBKE1K5xGwVupmky2UqOKC6c1luVEX0j96HD1+Bo8avivl0OTKK/BKur/
iNFxQny5E4Gu2bFYtoDKoIhLAHrpL6lSCGWdr1tC+u6gOYmK7u9JXYx176HbWYw9
BwpTyQqje2kvXuAtOV4LGYyE9T7lgB9gm9lzLyCxuOFymwwqiNZipW7I1HHYKMKg
KoqDwoyHWIRrmrgNKpgfQBti13rgiIsFtiypq8eUiIrIjeBdsSyhhGJtnYm3XfML
DvoJbaoy2frV1g+ibhuKV41A1fVTzdYXmnxd6NInbDV7arYBA6W8xtUKBlxStpRh
quAvemZNFjwXNAwD7cGdWM+QPGbbdoOmdasmcnC97WhBCiOdN2mBnn0+Vfrv+rTv
coRWYc1BRMtwO+D1/CD1sUhB+oGPjyiHSH+4x0EKvdmUULYMfsqKSZ7fr9nLU0Zm
ORp6Q4Y/NihX+kopHK6DNbSVj1pEuK/JfKeqjunqW04XoxBMS8b1gQy0r3ySDxvz
zL5X2NGXkayaTHPJWiZDkkv+r5VtaHfISsUJhAlowXDXaMeTd7YmaQ9RBsbeRfsU
mepLWu3ynD+07iU/oCAGh3IJoUH2WIv6lCIcsQwj4W9DSbUhVCRJK1neOQ7yOIS+
20odyK6Bq4kn/PGqA4wU0sYh3NvUcjLHgfug9LsFqkR/BcsYJvVGeOc7yTaiMDRF
LtycsA8bvhG42Z09eFX9sS/OG9Xm8rSog88Ky033STmpQXsVDNF2L+IOWcNn4y9c
Bd9SP/503CuPIdxa44QhGFrdPWyf7uf53zdgYgPriCI3fS/doLPXsi6FmGDiJJLy
PmoJrXkoBh3zHtsWVOUHLeWhLSY1JoU7PWMmjrjocTDNPcR5K58ejcOrecnGwtrY
kEYwe9nCjyttaVC1f22HrufavNBaSNOQqcDyLyiaoR+6fpUMjPwhUgt7sSFeNfDF
QSERHxeiMiZR6GpBCvfgSpVn72VzuWi2GGT+uvrHb6kpCFbnhQ2uCcLzRdBocuk0
gtHNFpPo3IkapqCC34zF0ujNpA6GoifGs5q/VJvDbBOOEAnVUT/ru+M0Q4i2MkjW
Jov6uvu8EG9cNw8sHlv3xUR+1X3pT97yqB7cXLg0RWJRmWeDfyMi77+RS2P9zPUV
fip65HzLSXtbG3EXpixT8xy/MWBqckSXwrCXD5zd1bhcpcNlpDpgoaXtKd3MH+tg
E+mVGEYnx0WRYBYgJ5ScdxwENArRyAaV0sdjulbKRoundBCPsWuLfa3m5p/HtII6
Ufb/OkuD0LckF13zHCKnIcN2T/gujYkBARpKqM9mLufyIT/DE/eB69mJHxNcZKwK
/6Ozb7jkWtHk3wUy/r4t2Rzp2SNgadhWhg+wVvYUQcGQPszoh0b6J+MPTgcpFpcn
Z2XA/4aGB4Ya6hcYslGKOiUWZPSIJ2rizWsvX0eVH/B5j3JTPdOrXe/F/F28XI1m
4oGHqpgDi4sSNhpV/oWA01lPSiSiGx/AGBXrSFFATlacxFYmrm2BmV3daFScbSax
tmA+R8bKkWTvdfEok2ThMZZxeSN+TcEZ8/bcsn86zh3Xpy/DOHYrAzaibJvFxJyU
f+w4k5xqT0vhRGeIxoqt7UMmLTM0PoxrW/rKzl77Mkbfto1/NpDPvhFTATh+6EDD
onF3HZythHQh+snbg9CXvxh4Kgc+Dv2KFaGkiTnMOgVPyiecXKidEbTILRiT9HpE
zdN5scnF55zLt7nMp0V1Do2W3s4psFAipl4jAHquz5rNcbjcQQ7BlZpUjs0U+lA2
QwoK/hiLvyMGbLd05u8ZWU1Ew+gwXsK1oJWn2gDUZPrLYfQ62r938/yko8eYDFLD
FTlVrYbDCd41yw6jK4GgkT9umLd0vXx1qJPioSOBD7rJkr06KWWW55nUlWyGCez4
xUJCF/v7oZ8fjS04SgJ0Jx0YmQmYVfUsdNHd//LhswDGa+sYd0sO4iEeGVLOLEJZ
WTmQH74N5thNn5WTx14oMCJ84R6MJIVaWOkIO7DSf+HaZksD2bHXK6XaresODmOq
J06UIyk3XaemGNZv0AcjyYAOip+z8yUeqe2KbSZNuZ3hZWwv1OcRqudtB1g9KGCs
zBQI479N9WaXvc+/O4FhQKjsYH1BTG5QeR2uuJ8upOmktqsLPjm4Avwp1EtfH4Fo
QtJj8fO39oAzBJXhBXR8cZ9KVCFsJBv8atkqrPfU6RuZTwAXjzy+TuUloIX9G6Ul
xWTflgxiOmM+Fl5uh0o4VBthIskopGbgDU9j16wZMwNiXEmkr2bmoxAJtHtPElck
Bmb/JyHZP47PLRkJrbKOEWVBhxTl9BvwN0T3oK5oaFDwG74S2RutyLGRsPnTB5P7
0iqgBmHVhnBR60JeUIBpIsaTt33zEMAALBSBYZllnO/R35WnLqPX2Mb/GkxHgDhu
3El81tHpJ4dXbSdmYC3rBbqA/oVHb+MC4FNvE4s+DM2IIIDo2vWegOBQIR7TCpZ2
6Y0rW9gEz67R/Ns2zrVznRsZUw65kI1fEAVT/euB2fCQNcWeCZJUosPdNNOfWN2D
ITB6fr2R8Lk/mkqMehn3ZRRMsVZCblWuHm20HSb+dbMDsRBRWDN2FktZb1TADfbS
8DSYZhH2ikHme5/6/GFPk1dJGuLJ2T5temnmb+179TBJuyPr9zzm2iT2BpV49cdy
BoPDV6qBdFTru4v2Ys6t5Gj1WUWiC+cFW/AaBTW4E/KAkLxK4E9QV+/qTRVApRCp
2Th4os5hHSfYso8tBJsygu/OuvnSQEZcVIQdp8ypTNSulQ8/VjYRY3OwIWwiSWRl
x2eEty6mN2iSXw/DzfXYFsG8GWTLHwPT2mGhbfKf6wSt/HwC69UruFq33QV7kIDo
GExr8QHVMPeXG3WlIqLLg6X2AwboRs/VRMH4PviHteokR4us8I8DNT3UGqQiAeld
i/e8iWFsPDvqQyccb5KWoU3ePkvt+GcR34uNn+wk+fPA6o+PK5e9kyINLU+o9s8d
ch7jRS3QZ1+KxVkkl3kbKfQ57ZLpSWkQprK1B2bl9qDOq9RgUBsNZGExgqogXMBV
pBWhESjEiKkAtSQly0M1qGG9jM3XW2BjnoThYoV5uzl4gUa6P9drrMoA4sEd7kLH
DDFxhj/PtWDIxzYXDkt3l5nbx7uf4Ewwo411idFO+sZk/bwf/xsx1Wslc2PUOWJQ
7ZMcA0dr0Ip1NhgAGMSk85OAt5jBPNa1M5EnVmHOUgvs1g594OJQCP5WkNys+ZhD
UoDMcQqZzViNRQSno+zK5stYV3KBO4ftMUtVoXUtMhNS9lrs3bgikWZoypltzmjC
zqiDHGIqxd/13fL5INd66KacQVQ/ivCL/xb5oI99QO7gLO3TCjiqA51Px9lyZtsu
Ga5kIUa/z+nnegtwSKEtk6oloWDxWOrfc1ktS2/2Z9VluZvlgW5vWifTcrJ4omvK
6ajHgX5F3z6FzdukK4wLlDI8OdXcBub5Snrg3lgKmcO3d8gZYxjwclHbziuHT8XD
RhLKBJi1EdpBAz1jy7BZH2GofyV8H2QvsXaDXLeOXhoMuY4iz5+zjI5TpgHdCSoQ
qvddQGHclPZfEjK/U8kRfx8QjmMLyGX9/7x5w+Fv0ksCWkIr9AnQP9aaNxt06reV
Iz1+WjNaM1ZvU8rnVB7MHORA0zgwWWNRvOXBcOxErYCtCql/5uk0GthwaB/ziRQe
rjmoOX6ujQaAdQc+ehiWzePcE+/veWe8P4qy4zbps/MDFsb9KceTX4TjpICNJNDf
mDz8j1q+/+C9udA4LVatrbNI1bt1yRBoL4v3+NPPduIK2cP8foFQ8CLOunb2n45v
YJNgXUwlTS9cliKD8FHjbVq6OoEgq12bl0cKhH8EErYEiBKYp7gQ9y9YfVOCN+v1
35umQ2owREg4W2oigEnQnkO96bo9Q5PFe+pxYNZPC38+fB82BLeH1f8JfnbY7z/o
KWQ04LeqMuY8LPE6ki4ZnOqa8pnrEs2J0L0xiDOfxuKTYQVRohBPokY0cOLtNmLq
wvj03juS6qC7WTYaZU2hNQhFNKO5xZFWoHq/gJ7jCj6/H3ltscDnvVc0yGzZQdKE
AwOXAaLzyz+72cGCK4BCPM+BIDH7GTdenPcv8fh2UeDLD+zivHLEZSPgyi5zjeDh
hyvwPXsTiSmFVDjLlEPYw1993QbixneB1QeyJbtZou58DTCq9fQQYUMegZKJ4bYT
JOEZLqEuQdTTwygLFKe6t6VC6rHM16Q97v7jAvJ9BXhTuYPUXpBTB9KELwOwSGMK
pd6o3rzCqHlbnQHnFJqTC91S3vTHiDisaMXbYMdtEryIlGV/x2y7BS4q+0ZzepNS
vjhgpthd7tz07kD8EzSlCysxqpNVf2YOEB1Z78HSl/28a2H9/SOlUxm0e5hcWxHQ
GwMgpxsC0jde9Sa2RLGkyB9ZUckRzOypEzSh0Iy1R4Isw+ppkq2EpcrJyF1DivNz
UmSygHGmL56yHOnU14EKQRW4PgFOvHx6T+hY/Kyi1jH7XEpIMHf3Cbah2ykkiavw
+cNs9tWjetpyB9tCdGjIM5A73iodJbegf8rEFjqU/h9Jg306S2mPuAzE74j9v+zX
xWw5eKKITcpHRVfD+0pnMsFu+I/bJS7w/CS5DbN3Kylhk16zfCvgSN7sO/TjJNNQ
cv3PbGKYfK1+CAgj6MWg0Ouw+oya4OP0sPKmvDzwci/4vTkspLi02bUKzB4PwKwZ
rCgzbjhYWbgHS8Log+E+apzj1UpZmujx5cfisutsWt/0PxFL7H7dXPvhPuCz5xDb
RYsd8SWyWNDtJxTSI4CO/oHOJRHzpe21t9pwoN3rJyheiWt5cgpD0/uKluTTpax5
iFEnuW0s17svR7+JgVviitDQieZu03ydnS+qhWby1smQj9b6iCcYD54DnP8QMsK5
A+/oVwWVxwHsbxGy+nyGH2hl7iYq+g7cxmIOeEu8T1XBY6InakrG/dviasRuBrsr
nlqKDMWqEM+/29NbD58Q0z5W0wPV07c20pj+cv5VoYm/elxJXOWxGfj1L8UTdcxp
Wv/dgogCZRVyQ8zjIGj99JQ/6FBGt0UmlR5jc3lejxWOSoIrY1AS0qzOOQ+9nUdF
F0hRbgbyvC6/4j3F+vpztThKNgdZcyL49zUOAtLjcTU4EhbFkWfhMwj45mMahaW2
s/E9AfTiPsBza8tdiDcURKFPE2VGGfzdHBtoF07axRlyBvIotCyjXX6kqZAUbk68
hbP6mhWC/QJT5ljBE2BBy7MMLgydTcy9vPuAxiTmWujP4OeG/R9XRt/dr/iN9FZh
0mb5vr7dWbr87DkPfjb3XCeHmow96dlcX0IVTKxc+z0fAb+uBVVCD152xkRg4ZFu
F2xaoiZzdsN5R99u13p81+xs4NUGSHxl/hWShI3xllF3MzpB3+zF7odaFKjJWcYn
b2Zrf/0LuyYOJE6gXrDhklqjXW9OcsoXN/8k4f7z0heEJvtXiyYqycAkEZK8uE7x
XF7dfin3wadJu5ubtVWQPx89h38XbLY4C+CoEkYJMMOzf8Ewgs5PUCsNb3ZCv2uI
Vx/AsS42WmmBiDbIxd9hRa3/v0trSVRakNDQ/plv4e3HANl6YijaKYyIqrgTaODm
wA8yAVjg/CWRiUqaEcnM2qJ5tVkxUWthp+VQ/qaZpNRDQfJgYsgSp78/gpZcV/XQ
vCirOsFLu/VBwVCi7GZBSUAOavpl1fVUPFJcjt90JifsC4YEpW3a4SVNojqrwM8i
U25Fra7sjHJWEJwTNscLNvwulB29cuklQpkWNoKmvI/9GUGQLud6q0Te/m0RSd8w
GnLPfHozw8yMczhxq0vNMaeqUYx6Mj+F4TcaTPRkiianCDQK+O7ZhfykIVzWPkIH
pTQ0W+VWDzs39eoXKvHiH3d3yTlgu8Tmsm6aJJ9z5Mz0CEFjJTjE6YtNN6EOYyrK
rJKvtoWhn0Q7Hpxs5+Vez04tkKWEV0TB8gmIT9KrUlp0VMAnV9cDv3sKZqEtRp20
UJkLqINM0rj52Fmx1j1ST5HTiS11/RjiHAGfR5pGjo1N4mQ/rzUshxk8ED0tDyd6
SWcSx6reXEx5j1136ZaTDe3+9ade5p+YHKCpaS9hDmNl9TKUgmCKk4R1eKLnzyCh
gK2GAP0h+vqj69WdHvQM566XnHZbMHTH/LEtrB1rVo1Tbh90auqOajkXcb38aHKL
q4qDpiq885UILnU+TFZKdF8C5w+O19MfdLDmQ1WRsw1uVklGG0whLUOwtz/GSctX
Z6dm09CjYWgxi8isdCv9dwh0QknkrVo8lhnOA7YYh0BStJVzEh4UBHGkjkAj/xu8
V+I2WtMRuVQeWyugG7QRtdRZ6Dgg/p9TYe44qOIySc/SMeaqDFs9FWsGjiDGjyqN
eanWkBM3FX9Ih9NLvxzCVoyzSDq3SGUT5lpdRztVo8IyrG2zC57ZnyKUMpktAX0n
LXiHwrOriJK+qKc6YCNxYZuq1EgGAPHUwjupf67vEqGj+1RYzyemqmzKoz61s64r
su1QmUx8LBMfEsu3583KnLkEUXjq7NwPSrocmyheC2S1b0nEuRPQAWHpA6XZE75K
co8Y1dxOJsRVEU1j2nGYu7trPFH2Jjy99Qij64FfI82gEiUolGSJHPk4TvlzId9z
KIUVHyqGcBAfRxSn5W6U91OZMK85pxoNbTXgrP3yQ2dJC73AhcvGFmPOfvQa/XvV
3orEgVsjrJVVbzFSg1Dy8tMtBp0ucjrk+F/aQKO46Vp0s2VvgM6CP3NEAhM7XJQN
FhZlkRMpnedS2hyrpNQkQ5DwK2Bhj6XT5hrMIBEvVFW3rr88a5EBpAjhefZue6zc
z0ZSqQ+V4K57G6W8XVEHXTn22nJlDNn+JLlNpo0Kbp4ssve6BP0HZPcUKecZRPC0
8P7bftac2kmyevR7pa5jUNazcqyJJ4fPlSMMovi2SnTswQoaLr8q7vi4g/V469/2
/YGSpvPlUy52myvSkBzKf2JD4c5Qoum5rbIuDr3wRmHUtvwyCBSTCLHkgM/5tFBu
IG9syKByRjfNbRg5Dl/L6V7mn3YiFd8U0NYqzgX0nc/5awbnITKsCNKciNF8As6f
lAk+uE4mrrNcn9mNvJGvWy3y3/GG2nbNd19xHzaXk39BGv/Cym7ihlrAZigRWeaQ
+esWQSMLLg43JJ318m1TrzzzhlHBGVM0kPlSHDtDp+CBwVJjdx9ftVGX7wcsHMv6
0OO0SDK0cUvYNtGTCCTnbV8ZezcDSiX9v2Oa8f0CUBUvdHTzE3lyfxeU5OHVJdqZ
0fRFbFohZA6MFJSRBw5UvtCLqkmQ8iUVBHoeQyIM9WiYvwOPosPAMwt5ReEPasUi
QmpfzpqzoFRZd8TVK0MmWzhV6KgVMxcLO4ciOu6qpizOyNiXV0+RTrMuQuXsgZw0
AmdyjB6UpE8UCyH4u9VRhhU8TI64Pu1iXhllAxExdhvqIHqLyvgmNHVCt4jn2vHY
boxMi1+OttwWK6UOxgPep/JTL6KPd1xDL4kMcThguyb+PC0H6GgFy7oRTyZPOxVv
9GJV9op5hjULeFi5My5qywIyiry5E31AqVNmyopDp6V0enBI1IDO2Fz5EjSvIkI1
YGW85ijlMbNpLyaiY7pEOhvqYfzEEA23gzFGYiKMy7HY4SWUObtEHkPupoQDz8Rf
8oYaJX18NJgD7ysh+85jTQwymht7Hjr/4VorCwGzcSstxYI5gAwu1Q5W7FpY7qgT
qnl0UsAO8/SSiY57O6uvWx4TjTePW7oAX6UWhR3CNoi97NPl0ijvPDg044m6KZsh
ozcacoYfS1g1xh4cL0iXLLSx9hEHM2uL6AM0nJPjxbNvswJmB8jKECWgwCkQcTbY
9KtFKzIK2G/gTM/PH9+Q7U3wVG+vPlULK0WjLWh7IMcGiwOPDkhCpYCVkNNG2jRt
B9SO8faYu/IJgZiuM8klUYF2c19CZeCBxoq1SIjYKorwgisLALaK1nkwbdl6fuBL
LCB6NTftYjWj+4ii3evOynZ2KJscb17h9a+a/3A+ve6+Adr3FkCjzBkT+6vfAJqa
QXW9jg/XGG8aGqnzjMYtg76ySMtuo8SoC1YnUd4h99Xyjg+8EVwznMRmtWNGyWsW
yJ8KaqQfaRYrqtWYewLjucWV32lCWrClKQ4A+QYewPxrlzmw+VfEX9m6e5C3m5ct
rZ3v5NVuCqXKuBoBc7w45MmmJCQWZeqL5+E7qG3nhjWnkQX3HUSkY/qEACKtwMWc
pJoqZGaSvtXU9C+lAzotaRHz8ZJ/pqjNLisOf+SYKh9CqF1BKpr3JRn1CLdiChtq
CXLeG4DVulT9uW26Nj1UoH+Dr/WJEhDQsvUoXGrhGQnGUZmMssR96DQu4s17EVZ1
f3evvUqRyJZgDVXZbaf7tUzmU72xu0Wd9Avpg+HZT4NVSdT177elZLSYgVRwtGyT
mVL90mjnGiDOdXdi0CEEfeECTSjXOCkYhMmPWEu4GkEyk/Jmu1+VNv/PLxAwxCT5
SFEUKgygOARR7g3En6vNB5XwNcmu2rQ2aM4KpKXUjmMthBiWsm4PFXrDr7XI50mI
xG0Lwr9vidKoU+Wr0My9/riyeCGouFawSvYXTOOP+KC9KUwkXDj5r5d43m4MtqVv
FhCDhF3KcowE0+TrsTTckoBMV3ahidAVmGEUMg/kscSd9VhRkoribvLBcV7mtJVQ
xgz5lHiXpmPmUmR0jcK5VKdk5TKxDm6xa5gzlYnfHwdUNah9/b7ugsvpk+yhNxDX
HPP9QBXURk80wSg9lpA9jnii2USEVNTAw14U1bB/UmvnrYWBFhsLklSR3wz5KoAc
2Afe72nlGcOLYWtN2cswAceh/pVexWIGNwGpcZA8jgqBcesLMb72gmvfqCAAtoA9
uo7TrpUgCl10pdpYOkZdGkAekX2/ZVjpo08o7ss1GLqNy6LGeztQaOCDUWU1UGXR
kvf0noeCVaRgfdn97oL1D1aR0Y5zrorC+OjZF3IaGLGAA1w0Mvyqxz3lti0taG9p
7BnL3RZpeZy0XPiZz9ApqsG8INMqOKyOEz5b81XmDawZk48meuTPCOxvX0rIOQmF
2FCyNopsbb0aKU1vzfw2rAPyiEWVYGIPnkTOmOkeiSt2j96Q0tuUZRzFkIyx3a5u
atZXwb/F9LvBcY5OGNgumKOeY1dvwwV3PASq6VyQmm86BoZI2o1nWoeq6EAK1+6s
S0SIyK2a5A+4FB58uCHFSMS1XDr1qFHlFDVwN4+dHY4x0TimzdK+lJUG25gzwAdt
TYgcUZWSUk09vm5sHO7Miy6CNCi/G4ysVKTbAuvHQ+uwfPZpaobkUpBVlDYdj63R
mzkeuB+yE0hTeMk9JTsCx1mDncnHaBNHHoond2H/5uRKCcD8O0NcfXm6gmPKUzs6
Pfq2J+uEX7IVCVj9A2RW8OBkhs7YFdKh78p21j1CBB3R296nDkScUT2F+ZzA2jhm
8buaKlwJ9vfEIf/uU+lovHst0SOz5GcGfiYHPIefRrxc2/aVa1wvFqkd0pCahtz0
GR635DZhVqYFUyOEpYYmWuFrQQSK83Naj0iuzdJpX4huymR8c+rEcDE7uMDHQ/Xy
s6CW+B5jjrNYr70cAe250ryQiFtzRz4kKAL8uQNrPvWFLuuMc6N8Uy2D+Qld2dnn
+IMaFDV6LHpql/lIL8hv0dDbjjDPQXXsp6zaCG4idYQFfvy83+yy9jWJ3M0xYrlI
972pdeAbBwsiy57BbcmC/5kLDDxqbVCvE+bHU28SKDovWDH/Rp6LkPadY/G8vbI7
6+NMl0EMx3MFyrxwzmRiuGlto9A3FoK+LEi+48B10Bogh8GSo2XnRTvk64iLnqbn
xuUtwwjc0d/fOfo2rsmWGWCQxiYwdoJSd+LFejOw3WfqR1pYkR4rpSQ4PVCYCud3
gGO/vXreLvH7TDsZM1yMqIW7O3eAxpe3XdnJu1ZQL037sq3XcvndcjzqN0RmQdWg
ps/gbUTKvKFJqU4/6GJXtG9/p3BdTla4S2+H9fCGOj+EucGDAoMj+v4fzbZMViXV
v6L4IvbybTaNT+c0MfTEbA1uUEC/1LRFKwRetyiQGJ/IGY96tjtMPPPXbSGGj64T
7wgp6cSbMkI7UJp0r5IOHuuC2b+UXDogePGUHB+D9n61JqgHpe4whse4lQfaoxoj
W5GlanxWz65jK7IyUieet64Yeimx9yv1KlPC8zVc2FtFfyEkwsv1Ynjoyq6ZBV6P
Efx8W/E6El0GIA6lDM8wjRvREj2SdKqde0U7PzgI9bRpdOGRhdtN57hVieggOUUj
2NtJYSRwa+5MpH5ta7Vw/xR2G5P6TeLF+HXuONF0i0jGSavPY1WEsfNxIcy/XhaA
GhoqKOfTUrME8NZA+ZF8sxEMPtblChmv19Dn0uvCPFzTpK83CEcmLVQhz5cM6GTb
RhN/0ppj6+HoIANfbzZ760cacQAiwbb5iNxBLy5C41zPqmne1ywpSFnQdxo4fwmA
IaQoKoLlUTK/eL+QXAyTdlBjFRlyHE7FpbOhytQEFi0cL7tXfpH7aO5QyGguH4e6
fyLW85aytNROHX0h77SMEKZ9a2zYWfdoE31OL6n1m3GDQ9vZV0ZF1xH65NUYiUgD
7gnfxk25aSKxBq1LteV4R5WViLp/2o9fQ769e8fuRaRW+6/jo/Ocuf7hiQjHMiGX
2SlqxlGacBczzBOeY4iaA9H+cpQnpzXxiT7lY1aK55lZGhQT5xOWgGfU7fIr/s8V
OwuUL/2S5pIc5HaNB03jgRnoUQzV/S1BGUaggXKTr7nqQLSam1uWc7QbeIWJPKnK
QoigBNtBt/Q7MG3TBJTBdYJ+FdrMbig2wJ7Xm1u+Yfb6LaRNIRHg++RAp5TxPBFh
XBNNO1BWFTk2o/eECrZKFEXIiVppAQ+2r7OMoWqHVu4QH19Kjc2jFbJMaOvyHEiO
rPxXT6eDE7mH6Zpj3VXqyAyML/k5fLih8sHUNOFUv5ta7laUaTCPsNhw/NK5gxvg
ejsPKPSbIa2GLyi4A87swUkPd355aWad+oLdL/nC4nSmW4IirTT/coSf4+SdQWcS
xbM83AVzYNaOuyjZ10jdTOqlTzrfBmuQCwBoc9dPKGO1cgVE/YNZ2wZKYiL0PEBi
ZVz8fuLIY+cuX8PZzTHL1q67VAVLZDbtVIwqNwrox9dWazt1EQsAZWVFkLmvdSy9
ii9MiJ3gQQwHY98+IjiC+AgldrCswJLq0EmegNXMoqxFvoW/MRtA/9oASXyDhwZY
Q+xg8Xx4UrRwetHDLsH0bd2T5oDFyb4JHSzMSbY9jOtxZbjVuJnzdNiSei8iMk5Z
u+pcavg3tOgKewnCgmpkY80g1jK0Ka8+9N7wBH5Hagg8LaIY3S8p9AIBRsy3ziWh
9Yj67IvgdYtt9aN11nlzIB/LNi35U46YGkkUhyS2ee29+mWT64vBMyKNo8wnGvEd
X96aiozxnd9trF7Ud6KtzqqDNgBdvYy9CJkk/29v7fZ/IddvKGmV+ynkMV8rj+MK
pR0lk1M/vT8ED94hYMvjf2KTPtXNGU1jNjqgrz9yZoB2NP8IxB4WIhtekwxfV9IF
fnIWXGSbyTv6PVd00BkYzZ5E77Kgj1nJlkSLu4SsZEKZAtvXl4iTeNoAvkRkOv00
pil0Gmn8eXEY+8T+aVGOxhcceWI+B37qAK12zKlZjgBcFDGJ7RNylJeAy4edenLh
QpHXT3wUKsugQXSPI7HYPPxyXePb3dnhFnN5d323rFSHUVi3uerlX7iVaj3gp7kd
ZwwXnJLXA+aSeSGP/6h8yxcIeaMNks0n+ZJDQMRSvZI0ov/kpceKyr8pVfzfR03i
sIoBCZwbohuC9hiTolCSGJwKWSZd8sPDZ6xRi5FIpdxAQuUJUq0NXmYOFh1bY0Hu
51wK+IiL4lMd7LrPqE48QypPLwOmHgLx5guI9jOOcHHmJ+tnanhsBPnbhS2QNcba
pq89/+VkaivCYcNN/iPyBWRyZimEznXy9xKtJXOvcZpYwLzB5tu7aqDdxTHnAgyC
YfyRqc3qBkKrI1J/FmZSnmHRhC3XkPiWIEdCocqJ5FFwEPyuELT/ncW3YjIGa78/
LRFJ/Fy2dfMgUdkxMjuddReiUZKAyQ9C+W3+GEw2jufRe5jLe2dNxFRKOtkSXXWf
V5Bk55MA9gmhVbQsvLInNqHIifoL6RJMi/mCiPZSA3rtXreR4y242/pX/bjq0BJB
mMEhH8AMW6Zgpu0jyALNlu98QSKUMnr62TT6ugiB0ujri91Vnk2M+UDyNwV5VOh+
bSsdLckBD2CXxdfwCe2OKdCSM28Fh6KFtpr/iPxIE+atBXG2nqRyLsAIlcSjOHEL
QKRbIGuOuwGnDeGmSeJH+/n1iJ/AHrXVBC65MPBiPRUbS61akSlyYIeGXmuJzvp3
H/cVJnk3Z/EM4aTz5jTPrSF/NT5BPyiNlBc9oLtERsgkixR1/0lHU0kNbMmzQHul
6XkXPktdNIkHR/vmoSkRVj1Oeta99OIG9VlNL5bjs0KVxzTiIqMY2HJgp3FT3gfF
7fw1QBin2KsP73QOKI+spHd31+Er7ZANLgsDBL65HJARIUd67sN5XiFEzF3x7sCg
AsiiribGSiDP2P/zTwOiZEgi0Tu9WkrQinX/fRO43wZa8mhahXWKhGoW9dsuum2D
p/bjQ7ta7Opg6QdXpwHTi0g7O6AeoeGmyP6RRtyoDMcKr2wSePcigdCHnCqdX05c
mCahhWzWp2ClbBgBC5WZKiJ2eTLj2zzLgk5EX5ZAz3aOxAkYSsOo/aSxaITFuEY5
y0DCewTSu6CYIBLUkaPjPfzPcXRH9sI9lmHflYM7Jj4V+EzV3vqxtXh/oJxLlKbT
DCzKjHHvGylCNUynAmaV/j9BvVHDI0lZ9jlP0UgxqEgSOavjOtZWe+NpK6/azxOy
BW4dYzczi36PmcEQdMJhTrkXEQ5v3P/q+lSWYAIFzrDfx/LEBQtSqHItlOd4IKpO
SMZ9VQHd3bwuahtGtQLCWlDFH2dbBJbTjuFx9l8XEn4jyy/hfMVwnn3q6l4sHtaX
7KT5iANyPtre+gL/eJ+BYlFZPkUToODc7XhDhTFaNsg8UDt1+W04e+L5DgG25Cex
VUdLhDDI+FBuXUsLiZ3dNr3VhJzGcHphJ7wGlQrFqdHn9NtXa5AvpH6h18L4SSvz
WHMy6UDy1a7WwGkkhIQzci76yI4SKLlO6VTKwbdkztqLc7DwiYNyRBusbYhcwyS5
Vo1H6P6RlhNfx+FZrRx1h3s2AOMKhC80IGjThjlBAVFukdZNru3Lt3ut6pW4zTeK
ATBdXlHwrG0NCkbqMyI8E7nGhsd6eJYsNejwSBa90J0yNo4E9TEMXNxbspV+vcQv
xaxUlNfkleZjcQ+HEau34b7AfTzwwlKakGvzwS+Oqej3qKHn0J/fwqaLBms5jGlJ
U1JDkxJ+LI8Pl5srXlf/OqhHfLls15a8kyEmcvo/gce39xRxDWrREwh5bebvOsHM
21UMQyN+lONtfbEFDgMY7O0Ct6lPxhtDTYtBroOGPFBp1zQhZBSvocnlxkENeZ9R
doOQ7mdoexoJ2feEh32VTKYQf+3jbZ0b83jEMoWzgVsk6ALLPDpgD3qm2fawOefe
3IpoekXWER9DrrlBunDt87WJTrYY3/m1tyRxJ0/1Feu4NwYkjB3dSqY+pBGCvVy4
/g/qQKjow9aSc3IcmDvcbFXqcWMH5tM/C61lDa9+4XU2DOkfMAqNbSoUhi0uQ48/
hx8xRjlSUPaGEztevriJGDq9y9ePVnShLlYgbmTsGbrnlqUbfyPtwzn2m4ocYYJx
4sln4wJfiwVCo3jbUzv+TCP0UMuGd8qvA+Pkjh/WmP9vE2uUXbxk3eM/iasrs3k1
EbR+ld0ifSQQ5z64RdmBHwpwVFcg/saalvLGGxb8mjOlxCqM/pOrdmET9F4XvqJU
OqP1FBDvnrgO8/YFjL7zebYlnAROLUouGK7o1SQx7s6C27oFkXa3NCEL8i+f+PCe
nqF4yibq0WbgskQftS8RxxatSuFmaK4VPxYQkmE8B5y2b3pFbxe6s59Ld0KVRnx4
MXRGumTd+6YqvX13FwDE91ZCdqM7MnPhHpIzbhL+Fg+CMr+RJNDrEFLk4ysTjzcJ
tr6pZMf/H9ca+SL0EMjOoEL8sVwnNgYYu4fIwIMzgOpfSig14gHww+0U9DWVbLOu
jOn17m+To+LwJz8GBYcW6G6FqhdTCEKL61EixWb1CzJktpTVrH61hpRyoaj6RiZ/
FgAgpNGUO5R9y9TRczSUYu4rgeNbzNPqyLSEPaOdew+lHmkr21ex4PDtqTuYO6mP
kIf+OmnHYvheeifJrBZQTO4YsPon6CszodTQazzcO1x83XWRauDjVa0+D6wKafBu
k+VXHIiEwMH+liQ5ZIk7QXtRsbuTXn2zT6mx/uUbBwG4HDU4T1DfIQpF7LixtN+K
S2H6PKK49txRaNBVswKwKsXlEf1ghilMgHEUgFJHWnsHm9EPsGoHIOyKnmPPJ+jw
BqBCJq/TunuMp11IQrma3nj1XFltmOCkcaoQ1lEsHZD3VUwJCSXfWXxZA4AwgJ6f
A8/uf/coVdPEPJd2bVv+42mhq9Y930PpP1aHF/z6JJhkCiCbCdktJKnyafAsZGKF
0P1ZpivaWuODktwNBHtpjQXzTNXlx84252Ulz2TY1ED28lUD4i629qTrkYoTKcCC
aAZxISp62On4pNMK7n+lbFI7XFjNK0XcSPl4jVGcrXnbX/cf6oAhKJ3jNjqWJqlC
MmlgB7nP7qT7uObuKxF7MVTBZURnFR+mB3X5O0APq2S9F2m9IGWlxyaiAWtHs6GX
zaZMbeqmgSId6bThH1lTfIhcM5z/kr2L9hkZy+2TsMh3mK5rFW8McTcFR8qpqGVT
ivtrb8W4VZAEIGQWYpob07nrfJ9kRt1ZJmFISqqOVWQKQtLnLVyzTnNJWdX8Vdc6
KVRgEtPOybAtkKDpN6h26TTROPd9EFdk4dYBUXoKVCZfBOBL5x40epzkLU9YkZ1O
tGCjHIL3g4wxAdm79uV/J8tpXj5UUnGPxU2uqazkXxPw28+lkLfIsU+WWbAeCArj
hmXqxBYVCB8Z5ZRShMas25o04iYko4i5jm9D6LJ99pN5iBs2lrTxaxETvi6PfQ1z
1zrK4ex252JYhLou/tH7VoPdDmAmpfr7GvCO84Axw3jALItTUnE9YrqOY4hgjQnM
grnIJGbjkpc8DLhr2K+ojiK5+0w1AlW+w6497o3BoFsanRdsUBXcXoeXJu1xNUIi
ud2SIVTjv58XZ9pg7KXKrV2RxMZJOYF02gbG2i4kzh7F/pzPTuCUJ5tdpabLh2DC
r87pVeOlkF6OFRu/loJvKc23HCI6fyozCJqf+PUbz8BBg8QRYW8Smy/rlpDZyxbk
o1GSE4+Au++SWIqXBSk+gK58yDzhpBica872tNeqDQs06vLFYZ1fkF7dEG70vNoC
EKLSONgQ/a9p65qK7SbMEt/sgTSSZvDWpMkXGZwAzvXpUbZ2CLRyguRcgKhp5tZt
LzOYCFciKBHUHdhXiy+Zad+uiRvSm8hqdD4jXKt1vLrb3ReE4MAOCdMfOZwahn6R
6qweH+vHk4fqXBQKNTI9YS66qSSKd4AmT6OmjxIOS/i/ME6ZmGojq/5eNr0C1Yi1
BeMRVsb/1RJSkBq5ftXTluvlkP4dISj/v4opX1S8i3rou6+s4UZqpPK2HXNFG71e
g5gLpt/G+t7qun04D/4H4ZNPBoZ3HqEOypraC0lzlka1g+tz7apMPF9XTPiOfKrs
v2RGoecsgfZSVJjbIagsLMLkSZNPhJgP9TQ6Jw8Gd5xfCebtaqRnZP4T0v5r/Esq
1YnujcTzmflPJCwH7MZzPUuwRAoU2YUztVMTPb1mzb59FnBlbPYZzOu9Ru4goiUo
2OBcvjc3VfjcSs6VUVcJBhZf7BC3hu9Ie//B5CM9w2JUcl8Yn0S8fjCiscxHlW3b
SEFWxXiTdPTSWhvZkH2JYHb9gB/fH5VHDoI1yk5oHG0vseDDZFdvQdzzuFrKfwvS
BknB2hZX6+HC6H7Pb16KwyAU+a2mT23EPH3glMbCg0l/FoZpjCKCCxiW8sfcfuLO
Ywx0TQuFZ3oL+6oik6mujCyIwpR4k4+/+AGFO1U/dkGNxRYH/vHaRyjrrDXABl8w
Qk3XguKbPGbS4T1t6yRahTrxssmIp5AppfGNDWxlNWsHTo3/02qVujYa2kxzMVvM
jhxF2nDbWfEQh3gqkrWfSQR/EbLzVsBPE7UCINWnEhX7U5xmdt63+3M92EGA874i
y0nP2ihPIbkEuZuRRUb8AyRFg6/wSGDd6GgcBzwPYAt6D3/zHYcSaNWK6GUHBrns
iLwpFx8/urpKjINGSHMrlDuKi4NClaPorlIE5PxVIQ3rzF6bFnMGJFWVpQbQQJhf
4FJynnfaCzUnmm8hsFWfnj6FZu7bpObJOxBjK5gUTdz0p9XXeI5NechkBg9AMiDE
Z5gQZomiSsK5/a50gDWBsM3dQGkfyEjDLeAMAD2Bv8pKSKHXrIByf1+YzZVy1xpe
hif6Sjs+6B+y7RuXdjdRIQDmUJ/J9+gPcKdE+G1wwVJQUA7sxpeirsbjJi7SrLJi
MvYplhwzfqETgDx5yGKwIR0plJyveh4J+YPYfiblpVB/0DbHf5h61PzYWJLODMB2
oqCSvFSbxSlsqrAoghvFmlh45A8Ch/JNhztIC+Qb4BR3Dz10ueUPXTAOyIMBzA8c
nhl53/6W+LaQK2UfhO5FzfoRYfPOBEZ0j08CYKB6dpCeM6AIeU+eF6wHVXHfeZDF
rDruhJEQQyuSZ/JVJJDlUsjsFKF+CbhsWtviPKeEFrBghbdkD1qCHwX0qAKKCbTg
8C4D81DKcF1MQ5WNIgOpjDWrfkSx+eWRk4j2Q3HGD8i3cOeov2AR/PuMXtgI8C/I
jx0oJBlduEfZRyZyyKtvG0FIHH9uJS3LQpXx541WV9o4v3AUCvIREBZy5x0tWWOy
XB9wTOKTA1qii2+pNwUW/j/+HRxY1QJKOI6FE3nUzs+I46t2GWkAhAH3q0WGcwoG
8KAXVakMC36a4i/YEA9lVtJ1Q+PWH1819xEeZ20r9NlvIPArWl9pAQciErGokdaU
NDPn6T2S+BhesoarmmnyIp9ELkWoByqZbbwKKUn7BbY32qQoV198QvEiLmbIpIcN
qcytAISaD8L6vHMdNoYOX2d+iW0m6EC4dV5eTZzMitAHy74/JJlReTvTvihnJLcY
kXENZkDmH4MscuNWezku7uSGadkDuELT8Hvo4FYV6/GALjo0G0dCAWbDxBt9Hla4
kjrJTdXgDd4r0DEE+Oi21YOT4nF8x55YktnrDR4/Agt5NopDuswOBqqkaasOH3yP
8B6yeDSqY5Kio2Wgyb9gBjbgwfU6KJ4Y9+ho6lO57sSpqyk3p4I5LbKoiBKdZEAR
75E6yFiIosuoxjAKyPuhaFvqVKs4LHuIw+K3JqLXIwDhUOWcFcV5Ndb6iH4a1bTj
YrcqSisdsVslSlssnMExDyGpsR+JfXrFsYE73tkU8mU7jwWvcg7Q6mt6WSKEgxMx
K2IaD6l1gnY9crGCN02F91inkwfBNvIdc5AwkglNaoU6HjmC3mWLA0cyBu4b3CFj
APPCZwc3JRgD+3bCtPncbQhrvrsh5ZK4EhB06e9la5lUjCsitx2sV2RG3VGcRO/1
inlSRp0QYLioOhvFoT3N+1yluTvVN1T70NL5PDRQgQo7IZtHMK3sNEZAMiixSVeB
ehT+xdbWblnnfKVPvOd3Qf0tFvfrEdCMmsq5NcUqBNBsdkXGKegblyy9HcdqWbyj
s/wpm3vpbKiLTow1O/n7EbXtsMxEeKNixgya6Z5Z5SZLUNYcvG8WWMFEZAXfbCb9
mDaMaW0Tockg50Z2S3o8OR05Dmc5VQGnoWvOG6t0na1xBxV8VPBgqd9KnvANuSFz
oedtFkR8IusaB6QQTg/kV6GAor3yXxLUF2z1TX/Jc8kXAEJJOqE4HELpdMooVZ9g
DpHcHEFzH7h/2g1Uo0nkzYRrwqt9XHRCUmmb3q2eNFX0g+mQ0IjVYCbFGntjoKur
Z31gN7WHManRXn6ROVG6K1YBgM+xNcu/ivoY9hqcAwoOkNtoEhKD/rVMK6MorWff
klVE9YWcsTqFcD/e7SS0RwIpX56Ld39t/dKvrvMhqS1xQD0jNTP8FkaRirUFtNJR
9bgLtPCVrm+3zdACzItU+XE1CP2/I6Jwqa1K1tNu42zhz2zMHE864hxXlYsQj73u
k3mL6cw2ISIRiqsyvuUVX9ys88u+GJIjvO7vwCuk/fQXOW8v+7b94DU5FrYYj4NL
k3L+LGpzPnVwrrH6diBCe7VT0T7lrSXBvWXRDDtLZQEKijL8coqNOjzWRzRqDFRB
nZhlOT3A9HMsl88z4Rd5QPiFTTW/EEWhz0pq7Ju50CG6/QignFJSSGLqnk4xOFXq
AXUcDdzkB+XaQ8tDth3QNviQcwRmVXJ21GcnLRqKmdoe+vldyhaCIsNw/jbmMHNz
R6VxVCMJV1gD8Wpa7ld4ianJ8zCV/3wN2Ea1Ct7WFC8+Ujw1hca1BY+/0U+0uH98
wrO94gFeb6w24Wi7wc2NDfSHWsaTwlnSmlJ5VR6tsmG6nrIE6u15ehNZkzcWy3od
/NsTyCPVnjj7Ra8JD8JsJs3NKXbt1k0+/PClp9VFmzahdp1RNEkr3cL9+TRQHAJX
HhIEudOEaIfWRxEgjHAaPGISO68twOTqhoSI0CK2UJ2uSkV6p7amQGWowgKhP6yy
wWzsr3v7bMiQVDhdLFIv2r7um4dItr9eXJIQj4SZr5zkKv2/kJDtyuFjHrxwe0bH
EnmumDycxULyfpCy9ajgVfjxYkuLVMfmaqAHUyXRtwdQwF6WiBEUaZu0OrtJbR5C
E71zNoPfPhHr9FAJWJfUV8DzTlLonvBWaZGdXWzJCDPoVZ6nkHU3WnaF0m0HWC/A
KA9IsZHETUulvHZ726MYazNqBhvWFhvNQC2iHUmHcRYnbZ10lgBz3Ns9Uz7dC7kp
gfP6iKeXGxihtKAQ3BfMr6WB5UYCx2eUIoHpds/CjB3mBzDosmqg68XFqNGd9jUz
jc0h50clnQfHoTQcP2RcsNWfPoqaTblvOAx60olTXCEzqurU+bcRryl+Xwv5xyyh
23bwSyim0j+2f5OYrVldDEFwGQKXUl2YsFGGXtu9+nR2UrAlKMOgFxk/KjYSg2jV
YAJiKGkl7sJ5wtjq0JntcDy4IVX7ZomOc/tE1729iM3r4TaIuM+2oSEaHVQzChF4
iGysSVgBFSyVhvKVJVPFlwKcUxyAUepRgzchZPzRI9ouAIK3Ooy3nl+T6mA74BuL
prquIYgjq9DYLHGykwxPaEg/u9unCfRBTWBmMPpJM61p0cu8Ol0p3yd/BxI3NdeB
wFncf+GeoDxfHukm4VEpeTRBgLfzLtGbUi/wrZyU37Cx2wIljkZba4B35AqWXPWY
0JnQenmAgD/hUNe7C+yvqDvvDv0FfM9W3vwvt7ehtOQBRYCnUnkKnUCqb2QtdvRV
Kbx2A2CmMM/mokjg/YqejKdGkC+q7f/pEB73zW75R3/XSUvC2RIt09AzZn7gmbIc
SQgSm9+HQZu9i5OIEFWCBtpCUcsa62o2pJwev6vnnAaryzcBjQ+CMIpMBwbnlZmG
Lm80cqEI1H7ios67n7dOpMmYdKbtjB5OV7CP3IGmoUUYjQufWvMLGwFxuTX6SSo6
GbNHLXVVRCXZQPmB6YchtuDkThb471buTgnytbUotd+zIhdfvyEqXsakMYB5cH9K
1nrfyha7ZJB0yTSDZcCOxdfPLa/1VGAWvril7ls9ULj+yVltWNmPsBaHSi7rblk3
j6lm8kG8nC9e1tVeLhpqXIk5L6V2UgKsYLyJEUdskU47L+nuCaI1+RghRWYz6sGR
EXY0cX4igl8okxRIAtcMCx7SU8B6+feicXDc/zOBOPOwehCSV+N+N40JPwXQaVuv
W1qiiUV+m2J/i138dNFxi+/VOC1cSmbu6OZUOhrGrvz5o7BJ2MJHYyOsQY2nsWOK
RmoKrKENoP/U4wZYgPKgyon1O3m/TnI1FLtwwQhNljuzcYqqXXPU6qm4yPVr1ZX5
SHKcOUbil+onWRCfv0UxAj03iNRasXgaJRMYjGxOxD5zcTqKBvuusVrkhy+Fy2HA
WFtIhSRzQ44A69G1tkLFNqys+oyifU3K6VUb8Hwm9V5eTZJLahh0NnMyqDOk4bNw
ln+AP1La8JWtseMB2ACeLvvUHBmFVPyC9usyFsXqIRQPGk2tB6QessFn6Lo3jW06
eUJ6e3eRGi9zfQd18wxqD/3GBRFVURfyeLkTD5PTuA319PzbKPD8zIruQSGN9NDf
d2i/4hbfHVPgDexA/ZlvZgKWdOVtxyHnBOmFim5EkEvdjk8aVmog7AdVoEiCYMAW
VRnwZLS3+u7lgghIFvExx0CAvs/ZYHyZmSjpADZHunQo6vHLpdKZoP3xLoBaWtHN
e98xPYTx6w3PbKsRqrNrwhA9UIZovSSLAxkTwRab/9JAuVxAJv3PJHFQTAJOSFuH
pKFeuZ9q2MRtpoEcpS0DfFlY30IpJQmz6seBAHq1pOdtroJtOemGPN7isE+7RL/H
xKd6pGzu3tDOVBu7ik4BruSCthOtLGit7mgZqdm1gZDNsYt06bSaBSWERUX/x1h5
Bfk4InI45ovT8KkWQJJmstJgqRdv49HgtWDRDl8kMK9mRF/7aBTe/DDKQQAsYXKE
1e1cEi3SdJ3qMIzoH0TIIR++83gX+/KPXSfTyJeGDNknr5Ues8dlZ6F3Cror6ibl
8P+uae3gus+70GCEuiYedkyWXlz+U37jKiPo+5/Qs1WHELtgtOQKGlJWZGGdpj1v
cjLgsRXf5Fd5wc6k2vuLQdIcoclo0KEXcftCfO7RkVJhDOYNMDCPO5KWcY7+hzqO
B6nwQ7Na7TomE5zd1x01s9ZUkN4ZdE0SlBiyDibVto2JEjKlGfG6zfnQgl0k4+OM
TLly7ZXySHOayKAuIspoBDdzJwzHZKWJfcvvFLVHO6zV0h5ID8n31HJX+FACTAAW
oO6XPbbKuk9oiJ7WWS4Mbs/LJkObxLqg/NS53ecDDqrMCCiT6wpR5S+MnPiIQaDz
zNgSwOIJHq6ApAi/8sv+Yk550TpoXqwhlAJ7BIQBuVRNdANCIgXV4WoHs0/84gcQ
8Mb+UU/mMZCwtPX5OMpS9qxEmdTgnO+ER5QPxIcepK9nHfPu09tmAYDNmMzdxfY6
cST/wxkCcMdzHLUsqPQNYaDKQapJryPmsUTLnwgOTpJrF43x09Lspus3owwmzSnc
nRl1bDJfX8Aoptu+DH+N0OHUHOcQ3dXBnS8c22uAjjcPJGLN+O1Mhfg9oBNz1Oxc
bMJ0W0v587hSMX/2Vs9ohq6iBBxUd14KuDrbwvZlITGDFLj4NuFtBYoORKxUF2BT
IiYtanpZWtLwPwiQBxeY4yFPNqWYpLoLedozhSrlVYz4rfMKSvogsSDPrpk2EQD2
0rBlVUszXMGRmr7tuAOZNS5RhNTjv7PWY3zrPPtPKZzZxkvDAUrnjm38vHvNZkZQ
gZwyrRRNhjJj7P2L5bTJlntxMi7yaFJGi6Rzn1cPq4NRKc1/5rkHgW55lzfrCCcV
mRaXRxoEUlRE4t+VvKLPjTjWVM1M8RBHT4tBtin+Tr2E/Y8VsquV/hutGIFUC0Ue
foe+WTrnbBj1gxmY5SydS6e+7w5yysmtKyZH6XFO4Bt19mOyR1kYMYF2PNW0FjRB
jAiSMAlqabNBPsWfx2F77QgIlTuC0fT24pHfDI3vy/AeTX4KkRm/AALrCEjL4WVp
VzgIbDTRlmh0j0gDpDyOve87w6Q+H5aqEOUPh05dS98GuhJbYi/taTm5Q+KhGjlL
kZhz7AyNu3WCPvzrMWNYoNav0Br7UV+BtlXjLE5+QG09qLtxLHvR2yP4Jtu+9ado
/YBkT5KB99kP6jv8I5TGFkQpMuSvL5b/dmsyTklyE/tJbvkkWG85WK1fhRDM8lUt
F4qusVIhc8L5DQFNYmeBsG8jhgo86Z2cVWp8SfiWnAb0Y8w8eeC6kVzvzz6pJ8xO
mEhpbneRlb2w9T3ySGSbKPKoElWd3UbqlDCkvgxJlLdmFo1uGQbHiwDxHG7vfVo6
uAfEw5rGAhxVxmvUyx7F1ZglHT9eQ19udlXzgKU3AHZWXh/wq/p/9XsNy/dAO+wi
r6yUpuTFbySHmyT2TSNylbm8ikLNAPb1gm7wkkVaAdXwVMZT47bRQQvJY/jqaS0p
4BPPU/QAeUk8AbX33x6pMs6mQejzWfIYdgOU1vaq8OkMy59T2NomgKLfBNW+HGF0
FdyME6oLypaAaKoLatKOiI3A+V3OOOOuXHnbIC5t1vK5fPJ8I6rJEy3FlWBcgN+l
gJ7u6TdT9kXmn1BBz2eyNsT4frKGx/kP86mignamiMpF4YQeMZcTUTlC+EHFmcPc
R+X4syjkCAMqbyKTsBI+Gm+PwuqUssATWZ0lFKPtLxyJwijd6OXKyCUbhcahkbb4
OYeS0lI6Jy9bZTnDwNB7hN05dQ66+JUJlijB/3HTG/0fL+2kdLTvE06t1IhY4YEA
qINaiF0uxoGuL31GIKR/EZm/1WtDIqnTkhFP43GTWAJNYjt3OTzs6KA1IzWzsPYN
gX1h9B5U+rhlHByBmnjB6uI61Qi6AJQlxA2ZHBjHazxJvBGWYLdwFeAJKAojOnIr
+hpDmC+aLjR5Q7CAzxzaG4h34d8f2qF8hEbdeQgmUY4T9fM/ELGJudto01gnXz2J
idmH9qMKjqQr4iPvVdEzx9gLve4NqppP/bfsQNYSwgDVPQs3X4pRZCzd7OPkPVFq
rvJyFs04xZpd3OuxwoXEStU7sNE5piVq51XnOC/lzJvWVQ/pNlRUEtHEtQC5fZNM
0ahE6PA5aJ8eXByuyBitJk2BqG/R6VVMl79NOz9FV3Kfg+cwMLLYP2RnVPCVHMrZ
AyCxhjAbVpxQnn4vJf0eMkd0RZEZ+p0BQHVADwJMKqwzaQLLlu4yILbWz9aFeSMb
3Kzla9Flx49XDtaWvdKK4VidvQ7iupSYYx6GoIWUkUNrAsjzhyO9y0ARu38g6kAn
mtr97BB1z8fiBdA2WmM1nXAMj2Ww1z8fkv4GHo9ko40Q+ZRL6eh6GrzqgYDuSp+Y
Fw6hQQB7xKyKaGEaSS/DI711aVDJMpzQjTmkXDbxhz3nn0XD2HKp5a1lNxoB6e06
C8U51le2hw37TaOljDU7Pzj489ATXm9texMybavMGdyatPlODkD4OZ/Xvk4cFgwx
eTCl4A7bXgD5otVjgJiw73h4gZr1zYzskk4EYdWb/BQ6ljj+kiQu0tpFch5Dn+3j
KO3pdYkEsafj6aFECng6MAeC09pMrtXmlFoQxcuiIyZbRgCtbMErLuc4LGuy1B7z
+4gRXYqqrlZCz8u6ZLr0zrhNNBuESHKJoIlEspG8jvLJFfIOVLw73/bHRcJXOWSv
3MYsdczBrV5pfE6GDDZG0rs5kuC7QQtKuv67ePyG7v4GAPJhGkwtUI35/C8tzCo8
Kykg11PBC/GvJYhZnIAyi13C6JOHjk3N3iAUgKtvFLNhTAy3ByOhug2ZKzyIJxVG
rmnTsPThFlcLgyUAvf28zLY3B5fG5WAn4jRhb6XSIkRz1gpOf7OErFWVvZUFhv2Y
p5Zonx3jxGTvHDPlrVslvJwdre8CZ6uPuH1JSqNPPKh9+FaxCuAosiUtuV5PYgfM
bE4F5hNMfm9klYb6Scglqtah78/rfKtPmH3aPaQ6D1fK473hYwTjZRvYhV1bKD6h
ZW+vPjlR6+uRKvGRMk00+QNA/heu050bYkqoTu8pii1+aWV7jOEhw66htfV5rlYO
97cqjMi2Rnr25mjEr3hIZHdTqDwMlJLPgYpjhLhzBVMWag0Cfo6wVOO0sK7OrW1Q
yFJC1U0badUtO7BGZl5gsEBTUFCxBYlA3Mz5he+W8DyCLLfufunmjMn3U0osRkCV
t9wzCWMUQW0QjmW6f0LSgv5MQQzdjU8OtJeo/LLWtIO1yXqWQM0pzJseHvaSy4cP
40C+xOqVK59OsI+SASj4nXmKF+FSjy1cGAEgS+07o09SQYLHhbLAkSWhgd8jdqox
J/XW0XB0CtPQMPE5n11klfQ74LmKFGjPyxBsvs95OXrTXgA98EoGdi+sYuEASlmo
VuVGR+DQVah8xPQoHGL+ipTn8TK9+XSXL4Gs8Y9c31hLLADRkicjBFz6R6E7oCdK
8h4rdkXe4BR+9Qq6kI8JDZQ2D7tC8vzYTEcncOf2+OeJ3/Cd9AyuWobDGeUGo/vP
6bBRFsisbMtaBBHPakilM1RoWj2TWifYCvTEE/f6v4c3XTwDOE8eckojWR1x/ctG
lXTRyqfBoEM9am2xX54hDsTsfIirw2b43R7zislo4I+TstHOXmSpqkHrzfHw3EOn
aBjE8eyT7KCKBQuGjo7sZGzSqizDTtrEsRq4XbpqsXTWEZ9f98DJSt/csSKaB8di
Z/3iJE+1hafpMccUbyd42yreZxApzm+QoPRUpmHjK31pdjY0yHYqIT9TWS28AvfX
uXUgTcgpAOk19mYAt59f27e6faq+LUFo3Mlp69q+dHFMHpkAQ5DnN4nFru10fFyj
SFSTE2vI47obP8Cp9VZVoeSlD9KhXU/NLYTB5T5sNtzXf8koRxCr0WRAq/nFs5Uh
SQSr096o50bSR7agn/q+Oyr6zLGUKnFwW8W52DXSTB6InAxhKyCIh/7AUHdBRWIi
nY3XYHdy18COToW/zPabk8G3l/f+UIeCRNwM/uMJjBjmWBYpGsBS6kKUTo9lej8v
95HptZxeLIRBPuel5wR7H47f2/WWn7IFs1uHIdbShy2Uep6JNz4QArtFvKWjFQh0
WbYEsCwaac9/ralV/7R/T5dAsJW8bkGCszTR0S54KAC7bUd1ozVHua5AbWd7DoZp
CKHIueGej48xQ/GKeeHgiXO+dX/Ri2FUrrez2745tyj7QekvGE90ZYzjUH/V6GEb
UCVycnYi97Kbot/j6ZtG5YnsvNMFbg4/cRtjBaGjEgc3yeSkEernEskF+YP7V9Vb
W1ersjzJn6itcnPrMrQfhXZ/rqse6LU1zIujrud+t7cCJu1hWkB3RX5BJgdn6SXx
azoKAip1THrPggYZzBP9TjaixYPkf5vLinqJWxy6t0FePTvRcEwkw5f/lCVXwnOP
f7VWMyXI0Yy8EVSv9vjpXakKcGzGmouiE3ETMF3+yZB9takKTbWXT1Euh/TXu3YJ
KAP/+9sMDZ9njcRufCxCQzHqrzT0am3CGaifEkpVPLDrosKJw9tR7o+fFxkwptji
/2FDXxUGP6fnpNVwid/kH1zo0K5lkmBfyqM1ddVXuW8/M9N71DXY0cLob9+P0mGK
lU1IXYiz2zphbtnjbfhYaNTb36QuoWu7taama1NZW3V2ApytCzFlDP7InO/OZy2g
+GCex8ro8AIK6599HkMwFvboPOmRxcMAAj0T7HC/b62CLbObjJuy1nUFPHuJF7kH
Sizyilz7vLn+TAqZ/uFf5ApXU5epLMctDZKhxixt7zvsUawsac2W9rjcV9+SM99o
SK/jsiW7Fh+PpE7JZ1U4igr6038C+RxLPvTwYNmmQC4bzPrLpHrYcuTWPZ6P31vD
jbp6dQFthkzTfh6WVWB/8z1vemJnQez1xULpvBFdvMFqq5f+myCIKn+iG9667zy+
7xatgTY+0xHnpZGdgNTL0niNcK0agp1HrmPD9gAZhw/pXRXNU2FzRoH6Mq5QTelm
Ptl4SoTTW7uVcpsv9DTdzsndLKFHobEGuwVHrsw1wplfPflZH/S/PmmFhgDR8JcQ
BWn0Ztefr3gn2PlqGsKeqv9/YNJOu73iAbYsjEfFr7sFImVztG0G7cAY7hA8M7cV
G8pTRsiKYpMwUkyx3xOi90JtfxNf+mIDq/8tb3dSrwBiO3l56TjVutTkuHR3uTfF
+K0yMjm+32YlXhAGmCq6knMcwQXfYoofdxgU6AuZYH6mR//qL7tLzrrTfh3bg1ST
1b4GIVBIBD/mBBXROqeClRKmsXdsupx0HRuZuqzjwNVqbRBvhZuPxu3dgpcGRR49
EWYIO4z4N/U0vubwnuVFmm3rbcIs1S8k1WPZUXbGmcqj3WlGPv1biWKfScFizgx5
YhgyCXo3PdkftOwX0ZQrDg0HmK4nrGzpYHQGPvUV3+y0gj/QrztSk+fidxm1CcHf
m6G2LaNpJ+7OqWlu+H90AXitLexshfh6qpEWQbRYTBXNdgDXkjBMlG4jpM0huha5
u7zitpxIUYUB4JH/oScXoOQnF6MG5YVhpV1WSuhnsrsri+CrBOGm5WRE85KWPRRn
n0A+pb06DRWJAMFha46Nwnc/EUIDlcwPK14I2Rgm0f/ts+z9lL6J5IY2cPRU7+ks
I820oSnA8xvH8DL86tXxc2Qkpz/LvApWw5cNfRnMR5LE1KZlv1XnZmQ6KNDBDo9+
QvSaoEnhtcE53moH3PQyyMGl76llEp5z85EmHReQmDVfg7rxd70GUDWs9+qGKEgM
l5x3wlVrldj6g43aWDY4w+l1F+d3adkZID/8zZT6KscyGN+0/1kJ9vOt+TFuVfqX
FnUicGsDLYXaa7/JIK6Wk10HsSkJEDqo/bLGmbI6AJJfEItmwLaU50rnxKHVaa2u
ZcaRdaXsdL2Al7X6oXYwrOM2p2/h6zjQv0Fu1nM8hw+upiFEfmNpSfl9+3TxbhOw
iH5ADZH+lfUJWForzlxIqusODlDMf3D36urFqw+vYyz9mMlphJB5sp8lfVjGvHGc
XhD6ACdct38jITwpHHqHdpeIpK5Z96tXa7NcCIhaFZI3OrCAWL8zStOHendc4PoJ
WEYrBv0s7EFw9ejAlEee0Rp/c+7kAYvWHoGUqpCc+zaZzVJSm/Wkiei8ZmDtAgJm
P10vn7CWNft/dp7frUQRozkgK6GTrHc5BLmkmgJO9Xqp37mJII/nHyLWurqk+hon
N/D1JfA+oSLOJ7Z/Tp+iqrOLPaCT4mfybNWC4Z14o0WbCA0lHsrM3VyUmg6O5gjE
N9Use+BupmvhmanGMZ4gcHR/GOaPvuVJKzSE49Wp+o2deT2drI/1Le4YcF2cQpRe
efsK5DObUGC+oHLjqBjHuSwwSdQ86Ll/2ma33e/Rgqn1S2rEQyNYESqPOldAL8FO
+x8+UN727axMpTKWb5U2liZZ1NXc6WGL7Vhgz+kHZRK4VbCQ2CEjb5vNTScQNtZH
gflG2LTokp+inq7ZtScTjTL8VkXUzg6IRkb3InPbIPO5BUZJedVys4Tbyv2fZdjU
k8050sDjwNbrCr00HN54GJzGMcS/E7OBeb+EcbhrPhjMQWbid6osePH7EnaUNw5+
kX2Gr6ETdvMe12DJ7gGNpu+h2YO1ckPZYldbxdGk7CZUb7hfGB57zV9mdV2erWU7
FMLImz6HWNH5C2aAeF1FCh8RYa3SzaCLIa+Eqkq+mG8jT8qM3wBRPZAGCo8iDmTB
hw1e+Pb9WF8LXFzqjqEbAyGWTz6TV7cUUtuvWDZAHG3dPw+X4LO/yy0m1z+8giSS
eq5d2poYQksPi0cPpSkjO8oqZkgdPUGeLFxk3UDYKL/s9+UFeR5/6WFvfrT09STU
nXJVWqE74iAkKhP1YFqfeANQ2u/z6SJTixNhFatx0FW5Wfrdtq7P4b2PMuPKkUEK
C4g6lqvQAa9O3CCKEYPsJumzgr3Mkrasp+MIPoxugh0VH7W0WfODuzssFMT26c45
sfq2Man+WUvcHNddUnjn8dr1kbIjw23NhyFYS5OKn1kjBmg4IFCouifLJys1IyEs
A0R2dqTwiQ0+/RaJdh2ITEAXo2swVLivCT8nRzenhqKT+Dj3ptDaQntWLRbdHpC+
UGJQdj2uysgkunc9g7Csyv4ZXnjt1evBz98/YivtN8YOOegjhK1/2e8CnP+weMjV
Gg+naIvH9EoDnNwzwYubDYmzGKJY9Fvor7A1SlLh8/jPUhBxHrS04QFaWkAdxqC/
HNCyz4fOLguEG4Hk3xmqGj5nRh3PCscvy8uOJupgrD+ahHH0HkrI8L4Ggk4YRm2z
tJ6rH5Cgo4KmIbdFH67gKq2yea4j00k9p/B5jKsR0I3TX4BTXt8I6DWb8GkTT2cy
xA1xIYAKAodaeJp1SxpUslLJlLXlaSguVdFOpsGcA0BHp1/u9wHOVWepEAbXwVcq
Rh3YL2c33dTrYwxYMU0tv6J2nRy08K3FGIHrE2JBYX33oW+CKdNpOqkwqzkUI0do
U9AvPzkVb4vnaaLtjzjPQfil3n1+KyVOA4aeSZGauhTCRjF/BoM8zFUV8c1K0aFQ
3sM975G+aiiT11woRvl9fuoeJ1e+ZkzFIeGI5+CpPp2fsGb9l19xCkrj977hf2r0
PiwBytO5irmWU67bf1fN0J6yVCMUcQEruX9KQJr5xz8osBSs+X37UtHIcJntbvII
QGMKdKqmDm8OKP02m2ldCNnAd4kfKjKJhFSUFaEDbql2vw3wRnBKk9pnuLWGbvQr
leBWFsPdTmIUbeA33x5gChhznmSnyyXXVyupkACqzCK1q6KCv12AdcZ2P9SLlTFy
/g8G/j/IRXnif6dCigiM0ndHkUnZ2Xdf0TrFHrPD0kQ3M9FliV0YGmzGDjTVeJDb
vv5fuUERbPl8FPqLL5rPJmaCLNM+mNMR09f3AR+XvP+YVZHNv62Vu6+kq7BwGNZt
cKvXYRsbiDxAexZpJFL4lnXn/UNqBXF0FcI6JLBtTSlSX6ghpDFQMHI0urllAe8F
oXR9018Cz5HmXPBZyLVt43wLDzQmDaKJdr289hQonAb5B8O1jBvQVvZfc+YlkNei
/w5jvxQ8QhbZHPtCWXj271irWpwxRddSAVCiZuggeu1lxZzoHdNy73JQ/d/aPK3e
1XjKyFu3blqWgwn58Q5Afd9dfxEaKbe9UP5P0VV35GHuTBnfPoXpet2McmNG85nv
1i8L4Ds5Z1Gvd2mIzKPKvZzZXTvb2N9gFR09tA7MnXhuShsJBKi+mDPjRFdIe7pU
LzdgJrpnbkDlIKX8kw0Unw7Rme9SzZ00mCLcc3+xBy2xEUtMd6hDFAoEWDzVv4jg
MSdphLU11hilf0mOsaZDauf+ZgVtDxJ2uy7ksnGUCIJa9Ay3Te1sIF/HV6tOYUmX
7QxAMq/b711Ggo2kTFVONY/7CD8FQkUDfGeUrShy2WaItfMOObinhHq9iMIl2zm+
Pl9l0pCcvxbuEImO1JcqHTvg70XBAAI0DSwpChoIkDUM7lqoQgyakaRFjxs+Bme6
pYVIPZSf90Vis/taYGrkMxWdSKPskU7w/33+9ogYbCPwxhlSrX/CPIz8JVoYj3Gf
bpn3C2HqJ5ru+f4Vk0Jii/0vrEd/2V5m53rwZyBsvrynQ2b2NiXkWEXO962JZ0za
l7q1/epPg3FU+RwWE9OY4Baw9soV0uE+84MiS0aw1+ZByY1zUu2qn5KlrmYu6iov
g2/8YtQxBV7JimKF8Qii7fg5fD3eODCMI93qy5RIT6KizkNMNfMUmc+n1FZCqiya
9VufBqfBGq2Qh8t3iat50KdO15F2vXk1YuuvnH4cUMEP8sRUj6oJs3hYEw2PnbNp
wyEI46ouLKEYf4bAfGFj+jKEJWkaO6nqNHjSM8eMwnGcMUxMz5ZizbqDq20SylLY
9PBK63B0Bs6IhVaG0yB7HWRcKO2QkiD5/K671h8yPAByCq8LAycrjxY5VfYbRC6j
WgXs5B06FvahmuNtmgCJT2v9qYPAePMzhga1ufpRQY60dpXdnFr1F2+sNcLgGWe3
SdxYfEPR07woqgnfW/WQoGZgMtpbR18GGI9oy46uRNj7FD9BFS1zv0MT44WS1D1u
PKQ5pOrZErJWg0OGe4Equy3zUX+atuKHlphsJih0V0oUbHZq0NSlxg5fnF59F4zz
j1EcKiGbMmQF5UoFdcaFyHJbdIcQbJl4fwin6Vg9kGW28RLalHbsorhM5oNkb61Q
59MHcOQN0TqoWIRHLPY4nfWT3btkCtG65TIuSjQf+4nzYEYgOnGzNqyLwDiRecro
/XvD7YdfaaI7gP2NFZXcTp1uPW3GHXbV1KVecmjDngIHxOR3rjjUOtakrjuYC/6r
aAYqzw/uXbptCHjzEEMHHE2cNxYJsCtF5j/AlpixX5bi3GcrhJW/PR45Acs+Db2I
QZHKeyeqWQk35MGOdpEz7v2EdGZ6MeaovW1lIr0ep2miSZF2h3Oi4Weir0t2/eG+
SxKiY6BwBl1qK5g4WJM0jesGWu8nziiHln1Bv17FzaXmV6IOQgCIPGJArA/lxV/M
vcTBoluhf14ouJFxbuFp42EckNClb5WiU4HARt5ejdVUZVAGh/yE26mR3UzzXwL3
kEzp33seLICEfVOSdaHZEPmKNKXr5UjUNTGP5yQWhAGgWa3YyCrU6dX9EoiBLHou
QxCzce7nolFNr7uT4WqOXRoxK9EoCrLbcnvatwNcry6w2ztRSi8ZJDlTXWydWRP4
ty+IDlXNz43bsg/Ocs9VN6gBmwI6KOJKxX8E6PAYhe5UiYLPRziS7H1tnEKJQYH8
001v+mEbm/aM/O1FkwGzE9PIOku8Fk5OCyECPEpfVFxdQSt6FHXH9MEt3uv2FCbt
JhoWNmJxxbp6dR1XxLmJpGnhKcdFYvJs5Rk3iMpZWsOI4nwrr5Is3zO8LwkcV5nW
aFfmnkH+6rqmVHSd6cw2C/7d1rHCTTXbWWXelvS+JNfpODM3WMpGFkn8KxbG8IaX
XzISgz/8/hm5O7b39c3XyQnu5PMfIyeOihkpKFIyDiFexDQ/cAhC92ewkDPW+cFI
7W+vkoaDdz5txNM7sRcZVqVGAFaMPBYaEfIKr4NPkdHoZTatHGK/z2Cj6nnb8KLR
8g+/WlrEBZ3bCTXe+Mu9qy2hQkGRAZ9+yzgGizt7z3peC5Hu+SN5vVp9wGD/UI+b
lJ6TxtQT+LyNRfd/TbVEfjl02uUTA9ebCfnbMj2F6ZpOonrajXs9/onlEho7mbBt
bpz/PkAcAaDJQNWJMNVVMVZhQlYu0G8MEAbCMcDv1GLB047wirHW7OmvPi+GIW/F
dYzibFR2DzQWgu+Azq1J2v3mXTjLKokkxOFJsUqD0cGDc1NTfI1mxoOD6YbvACtH
i8eTsfUPB+mh9JPKqn1IYeJWllui9/XM1/2IhMEgWuEgaiph1uwPFl5oxQajKHDK
odFkJHxw5ABm53kbtdpG0yC4EF2pCPKZM7BHsOSTOPKKc8SuJcIi5AF4Kq/ggKU5
rW6UmUavMCUERXR4E7Qnpl3swTE7qAGO1V5q98oW9a+giKX6AgujOIeEZdzzXC9L
SXq4sAD4Gb4VwWjr3hM/ksEnLANvqBYctVhPou3NsdSAVJd2iVpWi51tQpVrGGOz
339Y6XplRG0VF7c2PKsedWvGaYYf+sB+lo2LEdDfx2yKnsoUlPvjga+vAU6eV/6R
dvsWBrpU7moMLINYBKtsZoghCHw/okZHtV5hkCvgifULxRYoJ2TumDgAiQrlYs40
BYLzag1dShuUtiIH14zmpgRJqXHPr2FkaSF4Y1pP9lBMGO6x8kd1LVWJrNQ93kCs
fRvjSb/brZSu2YWFVz2TIPOumw3E309E42LUGZq9ILJgFv+qd8qs9FO1KFvJ/kqY
kX9+4iuGrH91tvWnHnMidApr4DFjRYG6VbpB8LA6t2xbWhPckbDn8/va9IuwwCaF
Gj+b7aou/+oZd5i8u08LR95x9T8qlE0utlc0paPtepvqfTgeSIZANURJCxKmRLrc
x5CLvuuQUjIj/ulh6l95h8nKsLOaQVLYjJ7ZTdSmB1qEl/rIroBp1C9m1zAmR2O3
WqRSwPf6h3MmlvqZarBgV5j7Z4wa6ljgT+WvcIfSM/MXEvJs9IyIvC65wPzhLo+K
twpdxlPom22IvPUa4MvDcZdo+pv5//jQgNE+RBF737tSVdqb6fMN0fuVVWrHWGOo
4cG5bGskoH7lzLtUAy6weShngapM4C08JKREJ8aFyfhCGw50cKeM8FXwPlvhXX96
2n9s282TaB1asfWwKxfO6jgxYM4CvZjYjZU5XSyeOTK3VCyOzr29zTVJHKTvdMz6
r4AV4ZHl5PcXegeCjMYJln5zefZvZdRZul/EQZWOdbST2F3aN2Xrxokh7ALuE/Di
Ohx/Ee9ajJL75PiGZ1GrqeSyJjSDl8C7Qt86xb+3FTY0irMxF7Ojj9e/6liw2Lqx
Jz9sVIOfJuvCUDSbiDU1G28diLe3L4Zx92mo0NVP5+IOTirSDE8IcxgkNHvZpPy3
/O0H+Uyn1Iqu+pWoKg2yfCj6ghriSQahcUV2yXuz7g9Lfnl8LgApYOQWMvifNOVM
PrioYAS08+6F+eAB2FtR/NbCltKUqOTsbEcxZdFe3fQuvYSMBLtrBiIxWq8E5Zoc
slgtZR8bM3virIjWuneUKnyeTWxEMt+AuvrEN/dtZTwSquQrFrdBAoztOVpgFVzd
nwDwDzl9i+MMlfVf1sIQc91/u1Mnw4yimRE67WokTdW9J+0xxxZUUCh/ODhXRiZv
gfvhkm5XRi1+yufyRfdoiDPfKzRevsVDMoGQ3BCIViDWh99Dv0kxe7YgsP/fH00a
fG5ox95mqvXagi7b6JSMF+K+rN/c966qgWLHzf1QMnD1juzcE1BEQ6Peh0/f0mf0
w1+Lc6YTQE3f2kxAtWD5+Uc7hGZW5doltwpHaE0pVjT8bBMO5axl8zZg+NdAenhY
WExOmlMsx9nkr+KuNwoEwPEMC87ikX+yoavJd0DNUSKosl6FI6w00RjUfnicOcJ4
oeATEqBbF29ycF/0B/GPV+b2Zj57YHVF149bSu1GlwNJcULQeD8JHFVwocEvfNiu
yTiMj5QFTOlA4KNO7ydO/q/LCsnyxfDTOaYTEKr/D7vxy5nyteQQ5Pt0ChcD8NyO
aZt4mRDl/7oKTCjtQB/Ox+ubgv+cpY/tXmBo3NFNRs5Eb4zpilyTH+G+EfN/MSJJ
hJ4FbGbBycH7JSii+BLTeSnkFZRh9yMBieG24jF6AMofNSk7m4wMbhCBMo0bLWmN
GFaPYlIBk3B1wY3/LpAVK45B3oaq4I2EUuHAKhm+3YvXJFdRY7PjPXc8ScFKCWw+
eMAorwXO7tLnvOEhs5cmli17bP+u6te8OY8FepRchJqSZCacDhNgFZlykm+zQtje
w6JyMPKgbcST6snrjd/0z9tvfLS06HK+0AHuM8Ud5r9N6SF3tlpPfHlT/z2/QqKo
MMWiLPOQKdWYUUC5WPeF1FTRUf/TQRn7/OYlWUo2bFhUrTGGJLxrAqdhfFsTWP19
mI5Ke6gC1aXcg7IwDmDWBqF4hp7ewXjlejc6Vl7pqePR5D771LszIG0tuJ5O5Wv4
GMCnXkd7M2CPDYjmikEQPGgSb5msbzeXUTU1LkUCJliDTDMyVa+k178z9MQt4sgk
JWmR357bb9jZj4+7IXxOB0qI8j1Kl2+EQ6pgzMnwD+HNPFeCiIwbSRNFk1Jw/pxp
eH2SSZdeG7g14joeMDK5n9NHuSAMYhqP2OtNXnHOaH+EJ9VSMz3EVim6KyYb/TuG
+lLrGbzhDIsLRxpv0DfGFGIh18kDOAZLV5R5Bb92+JYaS3j/hmcEgDNvHR2A5zCH
DzgITQiqjY7st5Ws0ab96C1lKau1PSfEwqcm0qRpTkDNrcujQHxDGpVif4YHSbC8
HdyJF2CrXUWjlep4tpfaJXMwnOHmfT+1R4WkDkVZO/HBal/WCbGIsyAwhvNXlYMe
+gwVusLMumS/kTEO6YMOCrFH+X/QfleApXXWL79cYKLryfHPD7C51Wm4BjYBeZwD
EKk+owNXpN6rtry4N4enCLoBvj+EyT6NoXugcz/isSFCXb57b2jNlNxGW/BDhUFw
/bE3o1IiFsseF/Op8wUai/6sznsixbIYV+F7pyh1uz+eTiQJ9YREF+P1uas2jDiV
tHgocycNI0V8Z50u8OIzCi5RXgPnT30695E7QdCan9Avqav8E0HDC+2zJ1UHUdNq
vfVWHSzUrDry9GrksGobF4oYkjkqO6fJJueveveBi9G0g0iXTvg4HgQwnNjr6oIo
TAqcby2jN/jE2nA1hCA8GJBLXFMT5oR4NAPd6yAoslBRiIYj14bLYgGGGzLZW0HC
PRX6cZ6iTeoTlDiY1kEL3FDc3AzR6N2wGwmxAPukCVWpjLcKpJuvvEBwLDRcLSOc
HD0JFO/7m2PGtlFgyXTm2joMcqCCTPJZx58kiLEv5v4d15UAPqpQrVsY0sxGc1jO
uIlp9W3mu0XwzYa/UOcNrk2WloqlgUqEYZ9krNwPbwuIjvUINWGGaGgS0i8A/UjL
PacrOuTOvoCLTzCwbmj30PWGJBkE3zQ6gG/hB+q/Zn32BHT5N2Qbncg4iU529ddM
hSyeiGFgTYdwVUShdDSZIiUIZXH3yYRjaXylKa6yGODbI35QAmOVjWnwGORtMWD1
Td+TwO5RWCkQtLNl5jAkd+pCpJlSc9kkqXuuMo1ISKeDkDLVNx4cVrmEelrsb00s
Eu5fbe1W7UMAEb4gaDGI03i8hDBprhx4EP7xeKUqCZykqDAOvTFv2mOP3iFKoKm4
qVoBn1JTVoJYVNECB/SoonjjCpLO0vFeXVSAlpzoCBqweO3yxNaBJLQAHwlf609p
mirOv96364o24Iw7vaq+dTDy3LA9jusoqFR4mHyjJX3oc5cARhKIM0J+r93cLML0
arVjeDvgXP/Gq7z2CXHFCOozWqjgSuITsWanIDCe5NkLy5OX+uhgHWgsJXsCIjCc
MUz7T+W3KcrXhE/yYBCzopZ4GZvSMCURdx5m16BNSYJ1D9Nse5zpC/xpxnysKvEg
yu897jMmDe1xViAQPqmziqN1BML2lF4VyU5D2eHuMzM4SdTElspXAEOirBh0KnMX
TEEAGa1uiIRRWh7zqIbyxNlyPIOwYURlhovIm6MkaWn/x2a7qLgc1QSaAyPjZmZY
CFyq3epOmAfDUwQOkfvSuk47N5bBwTkEAQoXe6lrfNKkIGEyT9FJYLtTSfey/r9t
EnmUbvZ9V0hc5LsJ2QDWMIEX0W0jNuyOJrcoT4sqq8bBBel/phWx2qONG0qZvqdX
vDKpwegOvB4NbIV0I2IjWkebPy18jJovhZQ3Ge34JnGtKl+9NCv8aex0AAUO7cxY
uEF1dFoCu6qmtvZC8b51cJRqaZDiH4hOwb22XSpYHJ35LVeyWr2ACa65Dgki16os
d9wSNYbg15EmFzASzIe55QMyHjv5YQM8546F2viHY4tzBQc5jkMYqe3zEJPa5Bp8
RCkR7TfMZ0JME7BrW4JUAqMm8f3jpJg2e2KnRB0vdn3njzz8bk43I/vrue2Quave
0iUDeKKHb+h/CI0T/WzzM2wCMFIDFhZSSBeZxP8koqm3uryZOTkXhmBq3KyrgTQJ
CHWw1JnB2EYKuLO22WfhdLJEbsYfo9p+5vYEigXojhHw4/69cJpEG/L6p4PvZjok
KeOhUCjdZWqXr/jI7e64x3YLlB+rJ++M61Hii3pvyt9SSt/zcm+sgeM/dZbRLXSd
rF1i8bX0ni1lDUudtGXo+4kjrVHHxx7GQ89Ie+JStBwT+2/+X+kf2uIvAEjpemZ2
tV2LNVG8MyL/IfLqApHRdW5es3teMosbgLiGKJ472hcBOIslpFOFttfKWBy05mUR
9o1MWWbyAwzpwjaXHc2WoAHv2qHmvm+OtNqvr1HvkqqCVaMenw522Hp867KHIl6A
1NJGTYlCAlHupUsw1bD0I0sEw4PGSVTgALaAJceqtYwQ4h1iJ+2FIpzaG1eAatA5
RM0vghVxmZ28SjixwmZ4OcsV0GRn0JOZ6wDR4OlY5ZGPVUQc+jOHmf0eLFZSKDOU
f983ul1aVS3rG5597N+T6I4ebFNTZeViZNHpoy14MWmJGntaTPLtnZBAv8b1OCNm
9XHxhbHZ6Aa7Jrn1ccbuwCqeDUPK20TiI1h2sasNDDwwHizR6ezFfaXcyvhLnCse
7iDVnrikzfsvWETJILYv1GwPsdf9l/1SQU0lxc1+66ny9DtCuRpI+/7Q4AWX122G
SnIbhL6pwokAUwu+VNHIq6Fa9c21u4DGZ11fB5v5ZEQ95D7MO1JEJcU9+MPh2lwJ
d5mZxGrkQVu8vIfRfNnIaJSxDfcJS8TufElMOXs6DAAvQlb4etIOFO0BE5a5eZmu
J9mWRj7wx24ByH7IDa74Wbes7bj5ky6hTICCjqrYWSWQvxYceW1s8zIuRd2H1n28
SXwJAAJCbu6TNDp4eSteiksFg6iXw02Ky9Nq3nIld74aRxDQvEkg2hJddhQvTBfs
29cOd1ccEqJveSuAHxVsKcjUdrgAZRvAQ+m8mHIX+o6EkH1m8raKMltMz0Xdptwh
xH0vmhLn1U1uUIm3cuVe93liFKhR2FqXX18ZYLa6Z8sOI6C4QmCX560W0oTrGlmS
ekpLQnHUCxCd3dhvGo5kMDpHpo/S28mB16bR4mFzpBzCoGauwxoSFdQY0KCZxtgP
SKiwDEF55yZDdE41v4sL5BFgmtI9fmlJzTftqOgDm55X7iVitZX/NgkjuuewtUhf
ecr2kEIkM1j2IMvriOVkL4bfszIpYoGb/xsLg5ddj2lgbdV5IRIHuqAZn8wESaTY
ktUR0RwFT0S/2rlCYsQTsgTb+4xz2pu4gA9y9XuZb4AIiGgQepwUXZnkG701WWgl
+nu+QaaK+Pj4o1n5lk1PcFkpirG6LlQ9zpAxHv0dT/2QFKEJM8pcvC4U868yKTy2
XQyF3H3hrwD+fz5HWb0R12dlkkJ/ILbzfZPEEzk+3P1k0jIB2z2aZbJyLDa9PdLw
v9RThPEdS1n98VIPF9Gk2yVrep7ZkfOUEV2SKsXt8nIraUyEt9lrjTFmhByrbQir
P+EBgxnyb6ohDIOFwywIJRvczG3gbDONTETQqY0LotbwfdW/09nasX1mv1GlqEBw
I7h020OrGzWh49YPFePPGRRww/cKnBYFZp6s+k5X2AlzAXPfN+U4QdXCC6GC7APX
oYAEo4EDyRstKm52ghQ555CRxVO5T5ZzPqsqkdZhrhsYQJZFbL4BxO4uce+IcnsM
jN50yi8uh1EI6WWZzYw8YjtC97ia50k9QcHuhQl94AXOoNtNlXeXlnJWPdHTc3qM
dziNypUACoohQWDFn5ZhSX14V6wuygOWG5Dj1vzzj6Wxd5cUkWFwkxoilY4IeQK/
BXv/Zdnvx94qZYS9AGXdER7S9YC/eLautPl9sdFZlDJ0/wPOS/pFaiUHufeJQk3b
1ZwJtjPuChKwzS3hVLgZ6Ng0V5mbejl2oxUxTZJWH5jcwuzYP2ECmkf4VwvN5PHL
Xhv61B3B7NOqHlGIf18RGTj8Mv4Hn0oSXofDfWAp+Hy7gmEpioCiRzhU56Uz1smE
4BevfrLcxmV3ML94ht2K8PTogCtlDs5WcaYlmclTb/S5w+bbgdeO2Xj1/q2qoRSq
pSsDI+pOY3eNEtLGcqC7lQB/wnIw8K69Bpfyzdi4m4UOFoOJTWZSdntEzAJJDrDU
aHzYpffsBbOegB7fM3o8AL4LPaPP0u9m2SHwTlo+2bdzvJCQra4DdZy2FlaMAs55
CGVbIHxk/8UrS8PMxl3zheZzgGunxL6I3ykDD7f/qQopDKGGKIkP9NUoKNJG4CWu
aiMhVSbjEFa/LiBAthHdy2ZUrVei9vhRjaSsTEn+O631S2Hwqhop7bBTtjZ3A7/n
mhhQGZ4M9u6XsvV3MC++WbqaLrlAQW2Qxf9sR4HOEjwQ1oiBTvwywuMudIDzBc05
/YR6zF+jpqG9LZJMu5IG3YJIzScUfKVWtM8Dn6gh4Ae3XciCfVAf2/J7cbE/GsL5
na18Y86tzRoUHKxifshOlQhSvG7NDAvZ/IRUwQrLVLp/xoFOnukeHX8WEOFi1qGz
gg3pxrefWAPhfONi4DiF4fPgTVtQGnm4RJwNjcCIF0FlbJycjStn7bqPDGgFt9ri
VEKZVKBkhhsmJVkbtmMb50NZHlRGObKIQOqB+Y48exeil/M8b7dXlNV42HC6m2T7
LFuD/ixfpVOFo5ME0XrH/Uz/4r/FvzQ76kaE6rDejjm2dHaP8txFoyePOWA/o6BA
1zPId3aoGkxWMUW4/zqJS0X1EYqJHhyw6zcXJjawhUS6X252eLfAKG4ZlJhoHq5e
YFmLjBIbP+0dYVNxdjaEYo3SrvHnvT4rvZVM0jdTtZmiar9G48EuexNobbbW86ov
CuiKRN5Rz2Gb6SY7l2AyATFvHMEydsLg5vFl55rAxUzCp0QMm8deAQ5ChtRF9gth
Zw28m3oTKKoLYl/7fWSz8Oxp/Xo8wKOBVxN+gy2ZG1pnlNam/4w5w6ObKXyDoxUO
+DjLXHWcM3is4PUyOSxL5dqWv3RCTt3APpQHVjpkZ2ZbpTtXsUXbNma4gHf/SsRW
epft8r67temmTFrMu0Rfoao2KBOL349/blVOVPV1lRg60/Ml0WkLYSVfGoEpx7j5
JTRvSI1qF8jTmcYhaBBUaVjn4sYBMczrRycyygiQOEhrSELBpiZNFOh0aNxxM3pa
P4D9uZgNWhKX6uHIu22RP2CRlM5s8D+SYjkn6AyI5LxVkzeeWzP02twU39ZeBJn1
Bx7JzCL/6n/2W7Q+i4bIlK4s7zLHsPFbdo8GYH+6NyaX2VwBTDtaa1MYR9CoT4UG
cafcqBKtlHxFTppHMfOjIQ5uXrkzbx+L2VtmxweBC1+nPuNv5HbiGkm1AwBuuWyk
8QdZ7qB/V9k4mFyZvC9lMrklzS92PZ6Amr4Q2e326rGHMtoJ5SRdtoScPq0/wI9R
JLIeqLZ9y/Zf98mVsyKpRwZp08e8GnpHOFP3DNOVc9/QNuwn+vxoalZ165JufSih
tUtGoxii9yljlz+OULxLMNflXcBGPoCofnO7HXWwb224422GtNgHWlPS2JgioGye
MQk1PwdVj1ezZaTI2eLIOkidAV3VkvHQ8QfRm+Ydmo0GIEbt6ZfFnUWxyhojkVfa
S+DugpFUMEShQ1a5VYB5mXz6Y8V2SY7pA/dASvGIimg7uk/MKpqZPJjtKQrBXFKa
WtU1Jl7ZaCcunN7M9NSnp8PPV/3k8UfTzP4dx9Irh/v8CSK6Jdyg+S+qOL47mNGl
SKvUJhlNXUK8hd6dnba8bQHE73nqUbfqeJ1F3UkuMbGtLjUq68mVvtGsTEkSC0Ci
cjqbqQjf16RdtyE6arLmXWwZBRqfCbnrJtiahANmZILSIaRWp4VUZY4NSrawzkHt
LUB8ps//bXMey/r06VWQF2vw+jBTDepdhBUiQLw3776cLm7U3Tj6eThgeks9BAAg
GbKJT8Pss+/h/7wZ4WmQiYpVeHo11Nz9hMQCz31bhLCT7BoeDIWZ2HuKcGh3+tIF
h6l71KfbTKBTXaS2nzfpq2BuXnxwcRRIkCs/A1PDRcjvA/jAi+7gbS0tnTKBMTbg
nhNEM/jCGa6DXVW33cmEGfdXp+gXzsrh5eE/ty4AisyxYKLCC9uzGAiU2hI//pUu
damghDOCfqXI5/6oXYkXh946SaOYikoNpbQFd88bMFqJkTSRBNuoKAQkXMM+CDnz
VGKyr8NGlE4NHszEyNyYmQd+K+sy7rCqSwoj7zGQdpUrFE4MLHfLGU0Hl43fbQ1+
72qBEbW66h2X98QPCpep45vze3gfr4PrniR/JJqIHA2yBIdB7dlg8yOZdK5+8Lyw
MvpLSHJKCjKkqfTyYq8eHX4Ud0Fh7cBbHa04apGzU1FDgv3GsvcZIWsHvZmOoCXf
lH6+7oAjjMI9y/vaxeww7u6zRXuBoHXPxGznvxZoSW9mab1HT9lL8zWwJYiB29KT
zghsgNlwzlJYWFqlNsek4XAFk1fPlZIxEHjb7d6DMtf7B/7s059qZNolsPKA+Yvf
X81o82mA0mqyEDfrS8lex5gxAL85xArdDKBNqPqEgEEvWxkvH2LYh6AUxPibNK/4
WFsy/CHebyepFX3yFQzMhlLN8tefUXs+DkwN3C4u2d+NZUompsApzIfscItCRgQX
Rkp1z5u5MiUtQdV3HqdNI3B5NDw4TVjYNExy9XVTAESrQr9P/C4QsQXLX0cM6nYt
qnj1jCaYw/yem6EE5XdJjt+Q4KW+XB1W6c7dmBDhcGi+/YR+mXtyBeJdRoA2W7QE
CvR5/kTwkpDHBjN0SNaTtDmyCr+02xOeeyARjimkknJ2hFOZT5lY5MoexUm+qDwE
MbyuQw0Zni9WNEL2Ibe82MjZftJ5n60D4UatrcgUFmgKkXZFeuN5qnP0BNQcy7YI
fsX+WELPQSl23ih6yzvxjKZh+oyH4uWZd3v5GHM5wyaI9apevEFxBJm3jEZqgwh4
/AL7gxgXg4GqmKdgBoMxMBG//biT5u2bma3+g/15qMr7e+LiZTWo0mz+wFmxWy6+
P8I63IkXB73cwhDxJmCxE9UeHU6Y3H6MERcnjkF+7G04l8anquSbSdxIsdjl9pbQ
M4kCwI2jNO9vHiHVI0hrGDrU+x/yMjKH3QVqPS5B7Y4kUzECi1ZNMS2d25ZK79q3
htEzKz8DrJHGnozWZaK9QQTLe+gxgkY7hdtMq+nf9Yghe/oWUyXbB3tPHmiP6+sU
DJyBer2VbpQY1F2TNI/uSbQst1VdXB82ENH9kr2TSw9UOi8hOH/GOL1rEaa3SXQm
vjCgx3gQCHlUdGMecUGv17NmsiGwCGp9gBK3wEM1f9xuAoIMMx15G7omEq9QBpEJ
RGIJ/p101YKMIMge/eaMz1U+7dvCwjW2IReS8BnfX6ahHUbhf/slWtup5wrlUAQC
GgNQfUjRCN+6fTupA46H9aNm2r1VgY73Glmay8P8vsVJGNxrWSnmeGcEyWWldZgs
Ht+PDitSzjW78R69EAJINjAjBs/uDsKZid7Sv23XtAahKpjs0peZUcToBwyNhDKO
55/artx/GPoGOdv2YyHGKgdeZ49k0bIgbl5MnzD4dfs/Iw9JYmXiKiyqZKiHqim1
wXXTtR7odzeXqx8Ginef9g5NWEDN1UmBH90XbC/Qa+E2sle9uU6TU3o3I5y+lg8E
iTg4kj2DMVs3QCiUZobOonVx75VyLyx9Yv2D6CI9YDCcs1mq3jCIkFSh3yyJ4gz7
qFvSh05sQzEhFWJCvA9oE3APj09lPtCZdD+DMWBAZ+hpFydFw/hvRDa4It2sY24N
u1qz1aVBtZS+55kKihQVuGHW2fH3G64WDGKLvMzSnlyRVXbxg7OFGpbW7EFoiukW
tuRuAG53cmN9i0uy6fWBUYujOgtHRCDP+vo783UH1rCGEDawz9u8FTkkeMnhUBKE
KsxgeGHiUia54/z9fBpWMzck8WXOSY+Y/4N/ba7zzq7MdCfn4JRNhbYrCPbr2Y+V
kZLpCxceNtALXHGCbYtPtWNhOWJi7wRrCGafE67YZGwGoKmOaZ54jmsMIYPrdy02
RPAAv6Fj1cSxJyQhDDrOc3tdrxvDRhwdctNSc4mChVCwLHCptkyqunihaXz/BayS
b45gDY580b1Sl30r2/0f3mUfEttHjqfZAQ6He6nj4kTnxqkIlURHG0fDyuQvb4iZ
0ABGP6PD40sLdChIqiEfXr0UFrSCmK7cd5+Po5Nd0L0C7MCXYN1AksWFNUxqR21M
Pvsydyb1iXrzNSOP1rbig/gu7Bshea43HlvttRW4KKRrCVIovOedL/PA8J2kpseD
BpTM1TcIFgPGV3AR0FJkpoyiDIUspfORev6olPOL2ZDlSvxbZdErjkQ0mjRpv/cT
mDIGCOdjxj67Y1H6GYHy3D0h6ulgb749ruA4XY+FKY/ppCwsMwUEq5Ilx78kJlh+
+imFZwDDEkXcPl6c2SMc+j5BzPeCBnQZYcjiYvQRX5CQZCTcYsNAbYKekTWRPy2i
i4i+eBk/kJtA336epSSta8YPsjMQmCuqbqZXdsDGc5ZrV4ZC0AWYGwt0WTZqS/tN
NPGWqM9k8jOFrWzU0/ogkE+lZBMwS1bTR2zknyzOExpR16LFy/4kTWvnSyXVRJCK
SQALgUTN7/G16g8WBB04LKDu85d/drpCKQiQjUE7QNpuXVR27K4dm7FfJn1QciIM
Shp+b+8TZunkfGuTIFrCvtvwlL9AVijZc2xiw3o7RnUlifAsxJRkIzCn4j1UeTwy
daPfZaHK+8Dra+dsCMID4GWZoMoIy2c96DU1vdcWWpo9L3TfvGiHhJJVofzb84JQ
I4HSMFF6MA746kH/PqygDlmU4bagad4Gj58frNJFXowBG3ZXaKSkzKwGClrccsju
ozTcddvVlfKTH1OryhaX6QNezOteyx/6HnnutEw4+cGGU1gpat9+rPGpk2SolZgS
6mirrtrdVNCFJ9/yvNvSQhiSY+jp2X9ds5Oo2Mb1VaazKWNq9aLeEk/PhYrXPYSX
D2I8aR7qSyEM0qKAvkJqlMfCJj+v1koLy0cYwvCsTPkJgPDX0adv5knmvUkFwCRV
PlstxBCrKaRCGcWt0kxF4hb1G3M4C3fH5BQ8Uk4UpcOznY4qIHJCXVul7jFmlco5
98GHM/9tsW8kz2yMSg8Wqz8x0vGTVDCuMyRp7/2YwOSOoz2yYqqzk5yjn9UajV1n
DEGU41dLaMWCfwtx+KXzDD91bkT6ADYKZaPFkCFbfMg6oK57HZxXLTC/ks/WbZeT
Ey8V7BZAv+sHOdpay6IotuXDQvGokYjMGuFvd2uLbOf2HCDFb42I1mhV9wRvQNn6
AdVkvbw0uYZE447UVIJElAQlHV3UFHYjnxsvgJljpWLoKkcU4r1GvwnCu8ibAi4T
b59SkTvWUao7hGN+wfBpo9vP+oE1AMKkpWiVDIjwQ+ZOhUbGjCWw1KIXK66OEajs
/C2GBegsAGZ2WKkCaUrzYPlyRJsonCbUrlmNBk8B+bAzZwmt/NQISLpC/64sWfpW
CrzSXcHHm9J6PISifaYsXiJ4HZZk9UxNFrEfysMaOCxg/avmbXwG0Uk1mBeR8ZV3
sRxCZNtdYccpJt6tULeYgA/tapfRbHZ/G0jbcWN4RYWQZR6vifTXWHFimfHkCuFc
a+tRParCP7LnCDVS/BoC55dm+kJ4QGOO7wJkykmfY001BVzm2OgNoSxJVjXuwPwr
EjQaCV0TBLkxJx97SD+UyiC34hGDgE3AABk8ATVq6EP3CHGHG+bgqhj/4yTIYVvj
xNlNLtt541QZKloJN74NA+OoyuGadEmocj/W5wT30HOl5Ro8xBhTKtct2hEwHaiu
FYzI9h2gOJWtmtb40tQ7/iSYm2FqYDVabTaNesh2dRwNziVrOae58fyfxOMdQLvV
v2yjs2PjHx9AsE4zMCuI0/W8R5DqYTxN9/ddUkROJhmUIuWZxplZev9t+F4jPdkd
tZ6n2u+OCx57O2T/UJXVAcZ29gAW+PbpGDD4hsDIguNNvUvir7ZJ1+lh5fDkxktv
zGDrC+3qaQcVe37GvlGKWnkHrXIQqY6vS0Pp7bZnKgLvyeUjikZU69p6ulda3W65
UsCPBahMZkmSePkPZBk3LH1fIroglxD+Hzspx9Pp6KvKJ2ZMn/IpP2+cMI7cP3Sa
Qdn6W69+8kGCAdZIvcYGlCDxYaN9x+B696pQ30p1c47dbEOU58R+kHjZ9cnWFNhi
Ri12LLbfrLqLVtX3q9oLZZRn8/zIpoW74/8nSkhBXxQp1O8EDx06dTD0lWfmPc04
BPVyom3UsJIXYdSkWVDvPsFc8hSkT/8j2BxzcB+zlNITMmXfXVVcsBD8niC7Xu22
JgS4oJoMiMQinH11j6HaaJYlCAbl7xVnukkts04f6vuKHEYqV6XNisqURwS9ZGbl
UtHYJQ7q94NnOCsO3G2EYdtprYKHvZ1yHeGBc1FAM6ZG+ifi4KTlHRpEyx+UdIIP
fx8Uka5iDzonmeaZMFcCUIpyGgwzN2uqxpoEixIDFJ+urkORK6OlGfz9QU9v6/bd
G4Bg6mi7k3CfLWoh+T2Hqnl1z0TooTJhNqZAYXwJsKSYFJt5aFbzVVSGPOvLtNw4
Z7bAiX4p1SvM5vZnJz/RflE5qQRHVA4XEu7CmBHRjnnc3jkX4aOqdkO5hIybYsrZ
aMceZnKRk/40Uc6PxCDYwRzkpke87YpXzr3el4oc3Nf5l3SqjkzhBIZfR9KIHAHe
KvOwKjBR0fPU0KllsO0Lt5hmMgJYBsK/s2qENudoBWyrBTiHZvH0f+DLt+YBT9o0
MUHJ1oY9TCG1jwdAANTP09lvM+injONJhJfVu24kC0JFs17+G8rXoZ5aPag/Af5N
lRAvbFrXnAOVBlh7rpCxxM05OG5lwthdy5xcY72YRggPq5WseuXmka5osVt/zpB+
32Jm4kHJDvntQ6Hxo3OQt0QUJ+w7ZvVbRscckAxwF5zavSf+UIaJ7TZu4pld78p7
smzRg3Es0BQt3s+U1sKAke49PeBKOYIWv2jt+TBs8FJKTcTx/BBcF/0beuPa6YvV
AlJb51MVsbbZx8XZ0gFJnrI9Ln+p+6o3bgonhafVllTOwK9ea46m7OzaCI9/M2sk
lgf5WPKYlXyYVg+k0dO+aaDImXHtxL0hXsHzBBdfYy3ACkstoTwEvkJz5OKgcaQe
/yVZ8utB6QIMNmZR1ATeNAfkJpsS6NnYHEqDXGw1HgVklWMc7ZkDlMmYI39re0tQ
JUzQDHC0kzZvpJYT/rVyUvaaeEm7K/jQC8nZBOnjImvfvwztzTNAirddrgnA7PZg
gNubBmU3SwQsHwyXFrNl+HE0bnCorHHn27965jAU+u81AxK9y/j8aJNmEupmygxh
ftrx7uFTuCRTIzfpnWDbBCH12znehrXazdvVwdoUZsDGGbdxNQSp+g80MRmfsVvC
HJgDw0vblu5rJ/5BdNfcQYCFOChQ4nFBcgdEsncUiLsgQNWY4MswQHrXEfndFWpw
a4sDZWBIRxKR3MV7Qpb1CeG8T7Pk6dRDgvmQBzWtW+m1Z2eXqxrA6RvYo+fXjowk
znebKtQA8afAgDOuDCTeiYfnpibD4YNd/PlJqwDFt6dc2zDQKJu8tE7FwLpoO7nM
T80KLDvcQ/fFjp1h4g9m+SqPB2cW26rZZSlpvh/yGPU4BXMDJZbNhtJpEsNI/v1l
6CLRA5sHPXxeCf5PAPLrXSi5+ySYAlwCXQtf9HJT40cQ8EKXkLLUk9im2Za0ovwv
uWd+Sk1s4gdzcEB5PfidGHUkDMMuF0L8+R1aX41D8zqY2yqnPUBWj8OdikBiJzVS
DAT/z9ZXvPeW8SK+EMHG8eN2njxlCl5wLXZmRD5KyDdyga0Kyyraq1jGvm+zDuaY
9Rk5aTOnUTzWpGcL0EXZ5Pqwv3NPyfDFc9IWnVAIsOM3dgaWwEc7nckWfBj1r4A1
Ls/eQHylPDnnFt06f4SVOQMbUuB8/mMik3P3rwuv827rzrdIpYVj0bOEfzDH+Fz+
YJp2huWAmClvsOm9xPd3Y4L2zttH95h5LpvM3LvRupQ65daCy3IvKjk85h0k1l7V
DU0fJmRDYCrAjPw3M2fAPs4aJFUdZZN2wwNGixQCYRkRbfOjdht0NL5REwM0/meD
ETTCcSy+sp9S+EHYRuNZtMOGSNopJJRnDvdPnx5RmGiGNuKopGH/aV9+f6oZgI1b
4RaZe4IR1pbgdCSQo7zXXB5dXehxfguqd9plP40IidxtpQ0Yx9Gk7OFPxE1wXcqK
w2lVJmwTio3eSSczkexQQb5M/CUyQN36kZYdKbOJVFWDC98OeevandwB6RUxuZ+X
6JBme/yj5YbZ5J7rGZcdAiiSeydmjRSg6rslNuSmIICtV+2bJspFD9Q9psAWZR69
3aJz93ab0c6zPKjC8m+mro3Duy9P49waLWLRssWdODwSj9dfHJ8ikJf3S1MDO03m
G/SQWKgWglh4Vw8orGqgOZAxFGBqIJflglzEgn9p4Vo/E69i7O7rWDs3MHe1fxpl
lHvlJbbPwVuP2zou6C1yLouzHJnh/DwesA/jT1BmFLGkv7FrroLc9/ZjMeJjMkO9
tXt72nbmnID8kMvvutly6DhADOKFcC8veD4fEI7kUB+I3gIBNGdN8eAhucHLFudG
VRiwi+ZPjeyTKpmRf1QmJb8jc4nwRHpsJzP4P65cEWU7QvOxou/FSiON5DVsFde5
yf8gQmLixD812Y+Zay5+zdgLYtTqwoj2GKO6MfQmGpUOi87+3Hwl79FsPTDTL5cb
STYLAvx1d3auybUgqjAsBhvM+074geqXlMSoQVldMHeGjH+K31M4NLxogTnqA8SH
/0vw/e1auvTMNX6kTOSGsJWOBRucLaogRpkcs0oRUt9iQYprSiMd+LtXyon1OYjY
B/IcZTWKDFC1u6I6mOViWYcQb2h517yqnAdMf4PyGB1y6NkVkeBtuTzAlg06zZS4
RYcWzfcry6DOJKjQ7GrPqyEWU5qFqPNsaCeCl/m3Vw2w2N+6bGkjy2XIbuBDj3+1
MvTVGD4B2U8Uz9wct+NdTByfiCt2z3/pRWyX8hbcMXM2aOBuR68LkVdDiqmXToIa
3JfK3/7ZnrZh2Y2Brrur5UPnM5nEoRmLfzuptMTB2dIF4BxAigIE5CVrM91vPqSv
eP2JYS2DVHJqiPJ/Ou+r8zak5XD4++n8BzyeLaVRdp69PahNPVt1NRx+X2R9BfoZ
3UEL2ltY+qpByteJpUpZhpZoMf4hfDxzWnPGNnsI2kwyv7ljMtL+lWjyDZxbUieQ
Sj9pjyIC1nW0Pqw39ZsResvtwXTNPWMt8KaGQ8hXKT7ZNjav++n40qLlr65hw1uO
j98amuNsl5SlbZEDV4zp2MmWtFxo+fMbUdVX2PNVA8Xz+OntKSv5Xfrn/2njYxHk
iwsPafD1L1FdR+qP9mq/amfk1BDz9qxVAhHeQgqCXvC1UHxHqfkjGHT+ou81ahAp
zCxLfRKATgGoXjtX4tubqBOhuigj5OJotihpm+1Hzm5x8ZpJaAQrOVTsNv2fUWKj
+xo7/1chup8TngqQRuts+JdEXMnj73q1duLDB4YILwHocsGu1yp2Zu2CiqNZ3wxx
kuiqDX0KHD30oIeOGy2zf23f43+s+gZ+VOZD4QA4bTIjProX3ZLQ7lycvr07DZZc
TbNoYT3XIL/PO7GW3jn4kTmM8jZbksYI4IaX7olnRODl/i4RDGh9pSYloNUi+q5R
kJoRWED74lGnhAYuFxp6hReM/8mqjRSVwNWJSAa1DDQLiMh8uPYwyDyKmVufhRqT
lyun4NjC8UJQ/K1EFPTNKbA83IGqwvcDqDCcuX/bE09frrYBzMM8BcWNfTRWDxxG
5RfgK7/nbGBusclQPJZ31slHa8C5zQZIXwCjex952SqadtBIXmLrooMgg2rIDRsU
FyHGiKi5hHrtZqIHQPxfkrZ8jmgA5Ww2ueIO2+a4pRYz+UtfH3rFn6ykt83A50Km
CyR2ru/b5+o1gHtvklil/fbmKExJSyb5gljPvebPtAg+Idr5HC4bEj8b2tEgZj9l
9r2Kvf1wIMZZLkw8ZxTCreo58+XM4LwzcyGaRAqIXpZWHvOGyv6jVl2C3odikHlh
v46czok9iy6Zdv+WEVl5e9sfOz1G9HdG/CafpFRU6U/2wfDZzJ/BGFwgMX3Sgy/J
uNrdeUW9OBLoBEvxfz8apfNjiK88grYOuqkWxaI+AXtTFzgLei/pJV5XsZW3sA8n
Ge3k1+7DwWw/pzsJ6CXcLdXHFRNnDoEu4/GzyJz8cVJJ/jmXydWu4az9tbXP/f13
D6H+3dxogu1N/MVCD2i65jlN3rCh+WDf+WOyjOi5Kh3lS1VCmRBKjLqDn12XXRYk
fk1VB3b7Es69Ky9NTHfxuFaaY9ds7im6AIsd80QqAeH8kCjJKp2iD87gwprRO0Z8
TEL6/hIHNlp3vTTb7MLyZvVdzyP8hlbZOmhtB+4iDzHxjxFq5jhfaJTgiDTIez7g
GPJtYk4OZj+eNgqySVwb8Fq9K0Sp1v0I7nnYuKjQIpQsRbyZENmGyNVBOxgT0K0N
8X1I3svtil2pFeft1QZyJPi9mcwrZthAeYmOyMhoiHsgW1K9plKjzLwflnyoDItq
jwXEl85RpThx3jrGdhQb3U5FOJd8oGvJpkyf74PWID10ZdCRvVG8l7kFVqtOKzwx
C4CUvbTb7qQyqe6VVGuJbRF6lKopV2z4aTDyUuA5Hd1lrV0NCL6dtmkDeA1t3D4c
6ZoKTWhrqJpnPWiCtzvKgv/s0Z7kpNEMGZiSLL2VxxZ9M/NY0nArKwnx/1VLtpuA
Pq/b3f5BEE2vg4Ty9VKg342UfBXUQ4BAi5kLilHc4Wlq76UtyFueW7Ki28ywtM+X
lBbOC/+lsaKqGYILrWMoon43sx4b/J7H87ir+r7FZutDZC48hq+hGmdh5P3NMIWm
6XdGnFQmeg3Jnl2RkvM9ax3u1nvIcZc0mE7vQacEVE9pxpzLxdeq+fApbOVKPspi
XSRayNbxOHbx1hw7I94Mi62oqK+rURtzRDQk4nOcG63XqGplg3tu78xzqW3Jrezi
1sy6YK5vKD31Yo6yKUDN1IB1Esi96tRJlItuoaLDOFBdmdGUfL2uwbrIRqL96miy
BSHkeYyNf4m95YjqKeAQBHXUJg+vugHNIhl0PgI5sU6dHOxBsh5bIz68vcSw/4xK
Cx9UgoSIjyunGT3p/kbU0kmnzEU37VnHxZs48u1VcafEs7z2bdYzrzY0y/QZMVyz
zh9+vhAx9bvWmCUIS15VupV+k3wE3NzI+IAw8N4o1kk8Ere3orpVEAs5glF4UEX3
9IDlH0/ou6TZ1hiDsxLwjkEam6/Or/RODMYdj1agTKIcZP8FQzkIAw1CSxY5357R
4JGoxBfD/N9h9sa8hhLZaEQFHeZqyHOG4B+FuyMR7jb9SIXyX7F6LIz1jUYA7PNZ
wIKRi7wbOFOd6HCfFCDLV6NXmJ83lwXf2tyXAPTRQq5n1F7o4kanpaT5cHF3Bxo+
02OmooWwTGoLxVkOGBJ/6IOHWCN6OWohFujmuXZD82Ex3Wz1GtCbLAgXTgdOXl07
ERVvaXGxvpCG4V3HLfOQunsYjrkSMZi6++bFIR4gz+7YFQH93ILZChZroyIz80/M
daRH+xfcIrDMa4HSsUM6sXPoOxYiRgKkuItk/cHvpeEzEVf+Dw3s3de6G0tg7sKS
7sVGBO8PtbGoJ9rQxndcusFEXKmpV+ur16oZOw1Ee+wqI3mDB/A43MYWlXQVsnJ6
eEn5zzeTaQLeA8MH84j0jsVG/KE465ckyjYi3z/AwwH7/S6b3UEYAMQKo2R7Uc0V
5Vp6IQ+u4mVrkywHxfA/VV7pwa3tMervEz899WP4k9btJiNzncwfztXhRL+gmdFP
EIeYto8fDdIfX4xqq9YvKM9QIyo3oAlG9LaowWU7ROc81RYUIfG97u+oK1Ip0u9i
0bthQrV+JTdbQPQXFmHv1OvzOUqzdokRpKhQNPVswxlJrXoIB3tbrQfvmrYeAG+U
Haarzfxk/0YawwQdRjnv7ocTg0lKMNwu5s3wm+bBYyxuvYylXpt2z2JScTDhIqtd
zc2JHDweSNij9i302XSZGh7u72XmJZzJHjnnr933iIx9stKFFUBIGZeEAcKxj9us
BXisMinIhU10M6laG585GVsRklP5WrYm5NWk0KGaHefyBmoibTt+LtGDXbJbycou
roF/imTCemAUsvJrHZ2yZURxuypSIMw/QkV8SXn+SSIM1iHahAmt8TdCgVp+Wc+k
By6JW5zVbX0oWXpMRWAWWuEbg3/B/Mw3FJ94aQiMlmmK7FtVErjNM9BUpB73xJW1
x9eKtz3F2X+xBx1iZyHAxcV7v/i+z/nwz0GlLecI4x8w+ibUIjlBefDHNP/vC5dq
W8uSeP3NW5oM94BAeC7RdGUiyc6EULEaXn8t2JwQcvXvb1MGjlu0Yfyk0vqOfBwE
Dxf610kgpfxj6fipBusfJ4vaoHfgatQEoobBhJ1LZX/OE6ahFnSwvOequxqqHF0m
Q6Pkwg1OKuE2ndGLRpm0rjeDIhrvZXFTC5lbRf8hER6nGkYXYVUZ7uRJCVav/c7E
a35xr8NbmzMU+1Jan/UOw2224ezRQuDRFnZNvvGmu27ZcbeTlhvWaBeiRiqBCsfR
fEq1pAImfV+LpAtfR7dYqo4qZU/zNcpmehHSC7wpjMgrStiJDU6pOy2NlPxqiD8s
oodQ2PVxcJxHEcxHEYv8toc6g3+Ua9zk/EVfiRjEzysKBTyyKArUDu/czu93YpN2
Bw2jy03FAd7M2k0JOjC2mqyXsPYGrnbfuzUpo7wPB7QtY47+WS3tWCm9C/DZS5iP
1+spTldMDPT8ZpRCIF5XNnkz2aUDdGlzldc+SJbe7serj3z3pfk3SFQQ+6BA9UJY
7FCArFj+VyJMhDj/VsT29JGVZ3xXwppPdTbdoiJ5QzD5Rd5xlQG/gURlP49phPII
FbqPKXJd3DUx359pSoE7WzY+VrUVkpq5w+u5mRnBuH0vg0m/4/d9/m1p9Xvz41jj
HZTG3T6YzOLMLiQtDpXoJklKegtX/7rBjpItkQF71I2BhMcH7s944QYtL8SHZgmv
EUT+dyOSguG4APU6th/fXFj5Po695KPs0n3mu6EvnT2+ZE9zmUTPPJ/bN5zccIF8
atQ432ZMSLr48zpWNmtnmLjERdmya/Kk77kLAiGG5UzyqS5TpRPolxU7KaCtP2RH
zxUdA26uxZXiTIqFgpJCiKRlwN0H40VvpZpdM9ccxbiZwdcsSIbenM/ojKd8ZaeH
ooekH//CHVjPzGGTa4d3JJQu7fKb/yZk35rSE8FQ7OOjFrLBniejaiJzOGhu2H4q
bsHFabaANBJH3EiUgLlNhqgJcmNub34xloMbLgO26yS/NUhYgzWQfKI2SMYYEVCh
yIIcUYMVr8wkAlxBCGHbCfExNKh5xIzM99ZVBohOztogRSeg25dzD47tzOmero5i
7pYp/lPzOecViZ+xf35TOkOtKzJhOwjxG1Mi+CeMAehJKfa9SLRz4WPlIgEZVtpO
kjS4tovULTY2OkOrF1IYMmbe01S6CbytXo11ZlHYr5ZYbSXQn4NewwwgzlRsHMEA
PuIgTYqIbTZTPXia67/y1PWHTNQAzUZ2aZnGodejFBnzh4NjU+/aUffPNVI6FNTJ
YogosDpVGIpv9AwTYT9zrraCS3abg3Fi/IrGKZr+bRAnUKAO7mDBt2agoKrhqZ4S
ttkPyNYUaxIX4eLMUSZOY4cxi2eGEdX9osczFoKsbuplOPR6r5aCvSmjn1z5d2QU
sRKpKOszvItMJ9+tVtDMC89qxshs1BwR5am1fwfFpjOE5PpENYA+g18F2k2rQgb9
rY6R3pshnEmc+C1jqZSIVNENBbQO2Hem5hMqAY1/fgxg5/XsNL1BtJdNvMJM3NJ/
GX47Rqr6cykBla4uT/8HAfhImR6R2wkWb8dDNnaaVzpBiX6S0cpeBFG9ghDOgZeX
nyhhcdEd2g5RyeBmV3VcqSfXaLdnDMC3UjiAd0whWNieVdzAJtsYfk40nnuD7FdB
Eu6y1tu9UD0JzLVAAC2TDaxBCvXQeYIl55CzBgHthZF6Djc3xN9vF+pfAWoPDkfy
jGs6J5X2gh97XhR/pKnqTEN95jYcdTMosABzHfgQQLdxYu02mF1UzHtEEQmWOMcr
z7sb/rN1NwUJ6TeiH042+VzluyVBwQGGTtFdbk+0+p+HbmIvFThHs5YUAyDL1WHD
P52Km/nOO7fwgh716M0xkHREJIInolyMpWszr1OzK2rXsdrwrHFrz0cn+8rMc7qk
UVI4pHyKLgfSewzPo8r8t12Bd0keN0fsHsNwiRC1lD0RNz2ROUGMtXyqSiPKVpIV
+Gbw/wDIdAzP/0jVY2AhCv0gAma+HrANsK/t8zPliTXh0yp1soeAhJKiktkBbCD0
jm0nLmPWJSNpByjnJz02VJT3U1O5Pot7t5LOGacoLQcO0vH479EI482QfLmDmuHI
ioPAfT3YUnXtnY2Tp6Bcla9ud4MHj0kKO/8QIirZjKnXjv3M97P6cldk1dl3A3tZ
1YUxWhBTEC5S5qG8ikqnyxaotSkVp9TY5t09jB5MYFD4bG47RHeGgqZieDXxSOV5
v19McCv6YUCSSMFNlYQe/TCwvsUyv1le0HqNEEq+hveM1rQ423HiLetamQ7nJtfq
mojEL0l+baYAM8D33iY2Kg8SuRCU7xgjP4rr4Zh71Bl8m7OJcv2mKxd9sSBgfdaK
XwEA11NUvtDytniaw805IxfHxdgjJ/W7qZk87Odyn/VOVv4jWTVeXv0uQr9VsUge
aXc0oDdB4AcCMzy05sWKstFB/ohlgHC04Sxouup71EL6D8Lqw/Cwf7VSMHb/6YM2
JDc7C6DpdTtIvACD21IXp5HON/XqYFSG20xtCWJErlQsdfvDWGxRcVYnCxX/rVZs
uAU5Efeb0aV4DNsuhRwAAkKeWnPot2t5HP0kUyqbXOt4j34HiPg1ao0/3kWD2kfx
xiK3KlbEBteer1cj8C1TIlaWQTjU5xBQ+IjjGQxcj7LuP/2YvwDls2KpmYyw5zR9
wKSNI64rVYLch4+9Ot1jCea7ngtWph1a9ZpFKMnn5i0SpZD9kYtv2BYmojCAueIc
dwFq2bEmapKztzs6iToAtQAeaZnCB3M6t+a+CJkTrgVHGPkTCm6mZaHBm7HnsCZQ
dxo9HPxg+T8jK1tbImdewFXMd3S1nIi/PkKOv+jeZaqeiiX8e9bw+cJxupLkllK4
+rTLmbiYFDszavcgCvPG4xX8ECifLRUd/n35OfE0SNBXbM+dxV3lZrdOdtDGBeVU
L8hITDLFT+NKczE4tVYIbixCplREcCZdPY2GFoepoDiNGk2+lLvq/QQLnfVFwbqX
QoehwxCY3ppZVQHCKvxbrFirrpBlK8+365cdhJN1WCUdumCPzzBxW84p2W8EwWkl
JxlsFH8+xAnCTR6U29vC0tLfkStN1IdAeAx9F243EszZ+ZCQvUhl2Stk8i0jIdFZ
N8KZX7B7zR17I88YONKQ6c5xCWT8zWunPSCiaS90IyEvE+yKXHGtGVWj4SYHkzN8
o/IfA/UKzb+cfpCCDHhn04ebRyVqP6lq/ul7vBZ0u32cClUXiCTQllPVi2Y6JaUm
eKyhACgU6EHawL0YHlLM1YnvVopxxauxY6cafO32IDNY+uV7JomLc84axKmLAoHf
AMM7iNN/mypPYo2kC4sTrAoZNg5XpB0dU96x+T0ExbVxywKKsTgBSRS/oV+SIf1c
zW4WspNLrk38SDmaUsegIX9l+h0MXeyy2gSKI4sh9CQn4ijfZYWA1tDEB2cnFf6/
tJAIEDmL/oa/KCMoe1ulAHK/yCWMWmFp1+QRIQfyCffJaWkEdj44D6sbRYfzjSx9
aHEFimdLX0jfdjXul1FBq0gvU7ueDTu/yw2w3YY/mBu3ysDeegcOho1dQN62eA/z
0rfthpQMTEGct5ecqf+aHfTSo12H5+pMiqv8G5OjGj9Kv95UtZIv6+Ow51Mul8Ex
UIOEzQdOnbnaFrSKf+wOtvODciiYRLNQtJ1DkqEfBeNud/YISYAA/aK5nEPaX+zU
hhcRRThXxM/BQbyp7BzD75otYM6HzwrFEdpZUzcZKGG+Jr1Hiapln6HIJnJZlTcy
w4XK9lMthG6i/Xbk3r/FbtY9BASeIXh5IQLpZmEPsDk9f9I3wBqhTYQk0a54++jM
Mj/QeksyubhR1Ja754kZdptsRURRWjdSdefIFnPNF3IXtlUK3+JBaNbnIFhTN7xg
gzbXcqqNvHiM2Oi2fx/RpsygZVOPenNdN78rxkn5gZEAwtCFvC2kqXOVGo5XQVNe
Q0lko/9hmRU99qG6JIuRQDpOKGxMDtfkHe9qI2rOom6oLozir9KFzODPC/YsQw15
0LSXM6DgXtEMLDNyyzoDMY8HWv3ig1Wj7pgDHj5RRRyrWWENTjKKao2yYir1xCgd
WGAnpgz95MZ/oQipswY88q1YGfNzeI9fDgy9JfrdA1Z/a6BVbHHnjr0cIMoa7eMc
+4via2dYOkdhS7levAI48WeM5jnXSM9j1ha5p/TEOqdh93cXxzrvgYubuATfoOa0
yNUPOK0Fi/BxFMVWqoemEG6p8nhS3VhtwrEnYSPO+ZLJ920KK93ArujInJXWL0hA
82n2p2so5KYd44Z+aYFKqIoaRytpLWeHb9Lm4YZJYg5yseUvA0lQb2fVeRL4Qxek
2THeUYYsqvQBLiaulRHugVqSWbt2yCSsp7XhXhr1IHiTUxzliaHAXfcvMYN0OMFa
sI7oiGZ/wiR9fiWpjvRpJYzthscyY/olYu6tEqTgMfFZZxqWUeKYi9Qg/slrNszz
k4QFVV+BmZVmVThAZm5ZqUlW/hEfXl9OxdN6rj4BRcE86ZJXtkAlnLxBrZA3WxBE
jucGF+tIhjP/ztzuym1BmaFMzyvPLNe+VnTglz0uFaYEnFtkEHKa31FV5ajMhDLJ
OmSyqXd9KDsR38NKN8vKo6UyabzDcN4EmfOoXNctneUqedLxSzXIiJeds04AOEQB
Nw3YVocEzNYxK6ZodUDPsinA3h91KagJIynbXVVPEKX/jNzEBH+nCC977glw/3U9
VckVA/tJjFNaYz2HiSX1Lw7RzRpgrh3zbPzaP7w6oSsq8z8QLORiSZBIsavm4Glj
rT4r3asY5XiHK4THiU08H8yXw2s5Z6cx0ZNvBIh8SPLWaF9QjeP+9BgK8y64PANp
h/fi4ghNrv9LhA9aAbzRRx7t6mhO2gbl8CsCWNd1f2lN0Rv90cQzJIsyeoCvM/Jc
FlvVM5Mdt4HaDCSMehrKUn8F1/dN0whUw7yIja7Lgi1rCueOjzzrNSh1mJJvDpwl
GFrYS3EJ19J3hgFr2l5PEOM9P7hqpHHrCErng9ds31r/k+xEOiaIjaLVjNq14XO3
k85ZFnOBfFILuolV0c/FxlcfKNW0Yqg3YHcohNDLb6T+LNctIoL+xdjSlhE9rTyj
WqBq7LfRcO+O1bsnvUhvqguJshNIm73p1FSbecDkMmHLp5KaAYzC2huE20YvFJEv
KVpdXz0Ykd0Tp6mv15hLfg7s+yQmpwqt5mGE4l77dabXcYEP7J+qfUOgDw4P97Tf
WGqrL1KCrtZf6KwL2fRS3/7Bdqkh09gn8CYdWOW2qRwQhEmqcyr7mDLWxQrFzQJr
19DS4cL0kOHKuBlXKnvCxMvRgirIk7LPWSD8eFtVFwLcJyJTG7Ebh/hLvCZvoHNh
Enw7WuCA5mtjX3GrQUvey5s9uWv3ujTaoSF+YZ6Ht3o0S6Gs8BL3ZIqvsUyV8Fgi
UAKdp68Cj6xmj0a8oZYvaA0d9cefj8z9Yjxe1HZsV1jOyJHJ5HAzomOxx/XokyBW
uKHmDKkVeCcyOArQG/inWWwzVfJgBXx8QKFcgdylyq7vogP0t68yT0Yiwrrpb6Bs
FTY7DFmFp4gRRPicpSQkT2L2KcHtEFs63WAWa1T0KnjiVTmmo0njCdfgSDtffM0l
DCmUU1RaUW73zE8Osg2xPftj+Y2xK1/Y+n3h437qo7ilr2vrdVeWJMivYiwuoUmk
MCQqARgcnFTMjJVTN8o7+5Ey0Q0tdc4lXr3nFI1aGHZfC0VxZE7QikL4Yu01UtNY
CX0YS2EC14YqbcNAZ7uw2OoTc3nNz8ZFIB6aArY6ZqPpij1MG+H2Y0esAsUWgjfH
LBwKn4NvD4CeqUV1z3Sz/QaupfavirJU4pDsrEsqfsAgPTZK4uxarEzKLPDpljTz
zQdZ4BvdBsc0gh4A7rQZGIcFtLsof543BzTJXKnBzR3AVPVDN7jJY/Bk4ebfNPk+
3c0/SNdzm+bS7hQ40xh6ioTMgIfBYBouBLRO9LJgwF22HxB1BPdtHEF4XYMYMVD4
CKBiOT/YUb6u/RkQh88wLi7NmMphXB3WweliavxXHzjHvhoY6hmhij6H6TVean/z
CGWjvZwLWBRLjYMVReLAJV7WYEQWlfYBHnmaypk/qCRWg1qzsb2FgZ7oGT8yIbQx
yjj/F7ppHMXnCsD/F9EBa3dcNUZWLJSJ+FccrUcu61lTv1w2KYYwLIwXU+RgborY
CgxrUOr0IWGhL/D7nxSVFLjZXx2r5ymcr0DBPb+k5Rfd598BwYj7Vfo0mWXEWLqA
TSDnPMUbA4yU0e5Yoz7Bjii/IL6Jp63LPKguHt+BJOGcn73z934atXXHezCbFjG1
vHii9yZwJrwxhyNOyepfOrfIyNSvaEl5ah2tmEM8FTfyHs8E5EpvBwZArnlg89ut
r8fyDUwwO0lUp35v1Fhqjl3iMuPa3u23uhCotGQbWMsyp0HOwuhqogS2NHA3VlBO
yj/mAWD+iQ4Ln5jez01U7HfsSGRxvjXOK25MmMVPsHIYij/c6S5KijNsk9IK4+PU
ddH//ocIMhB/+ziEpBQTVHCyy8uYehteSvghEiIeYsFW3f3GGW2UubU4ePgaEAq5
5o/sJaK3lZRoQ5c4Zm6oChUGY4M15uxiJ7hHH/+vnGHXbtWzI6m9Bh6aTXlGXfY2
SZhlp01jVPvhXc47X/0EibG1MNBgrEL0peNpEjP5962LwaeX704E4/B4cvPH4pOV
Gy3OseariSp0vfgudNGGx/V+D/HIfuQXaRU4XagL5PvWn+9dOry+AvBTgNvyL7XP
Qjh90bOpgkKIIdM19xef0O9e/1UlgdRessDaRWTI/ynH3vC+OOgV/SfgFeo8wQav
wPoO4Ms3AmtS+NYdCGpvMxZ1lgwMBOxjf2VVXPsdtD2aovkqu21cRsODV7Upg8ML
o1wL2qJ5habql8lNJyDbivB5IbBkpr2kInBdFUIaomdod3GzQ2xP7i9qsqYCnAuQ
wU55gdJewjOXed9b9HnmnLaBsfeNOle6hhGKzL9EriiTSyyMGYVsYtC4/tEPmNV2
S1xbfgvRCSscKXcorcIbu7oemqVuljap8DNrV+C+RNEoal+bLjspmZ7dK6hZ69K8
pv6c1e6B2wd502iSwV+NsSUntvuSsFTR+O5ZEZFB+fGXOeMlugh2Le2my/pn3D+n
fNL1RZPIRD+2CoP3l7TphbyJkeexDHCfbwFeggKTR0lUel4ZhVbcd4Sj/Duf9fUq
IV2K9Il2mjIMCn2orqTfj7kMoojpsXrw3HUU2KZ5bYyye8+8HgkNUNDGaEiJe90t
54YnTVk5YH4mTCAXLtouMbmbDGw8C0ATEp6U//iPYYZ3BtfrMVUQvX6LCL3zzqfg
QXIrVRM+nPiw5WsHBRgEyvQqXwPY1JwrcAspd/XXGx/G1svGkP1b0clDtf5zevHn
rcK8e4J4nOzKaj6oQyv722bPuusMXp3YjXmnJKrIlAGlBlE5YhoLAEKDHR9TyMlH
lqhoZiWLMojGX12uvPbsl628PxnD5IvB1DDsbK09ZLcRW/flcF5jfTVO6GsRrVDB
26Hnh6vF2YsvvYlktq9JRrxeuXr3ufcm32nXvtMUjFO9uZzOQsQ0CeV9hy/qz0gn
jYvr1xpUtT20kzdC+GUnpmxGOshc1ycki4J1VgoJguz3JTHtjkwemnwADDQz1VXq
FyBQVdOfAQf0+zajsZuXrEN8YsH3GZEEkma+VF12zCJ6+fbsPTEw/ihMkV/0raKl
g3Ba33hd/dyNmPXLi1xLGN1emQCSSu+YGA3SaeUe/BwTqePpLiuXqyFk0easzVcX
4sE0TzB8BeZCWHiW5PQD6joReZHTBapm5aa4FE89yKzS9mLqBiNbXfpSuyZzn1bY
0HDabB5+KLctJFtgLs1YuEG/q8y2VawUHH6xx/5/fsQh2+OsLtcJVeOx9dNHQGbG
s2N+x5TXx69TYwOEKMQ7WAKt7vzebZ/JWzA1E+YkvHdv4o1yMWLk2TJ0g771UiBm
M3ZvDG5vkaQx7/SdQkQtv1dUs16ttAYXeDuvKW4V5OGbDnAzYXKiGtlMyuviOhH7
Ixt8FVBbBTZPUMJyQb/uYUsRYQibkDbMJ4DrLWNH4D6zt+sIhwHrFIpfaJ1EXION
2VvWNAn4liMRjSlTB002FjztimNjRMFNRNYidp5Chu4t2TjrxUEyeSqDJBbnSOpc
aj/ZrAY92/D1q8nOUcdY+frSfQLwXFaj2rJb0ktF7sPYic/cXVMJMOtPFjdo+R10
SlxKON8VwqeDK1Fed+ZOu0TkH9MoZ45UpvwVG7zxnnZ+CAvS60tYSLr3TUXNTPZ9
RR7dHiwRKqE+4SS3IBJBudulI3cwGCbGZwIRqUE/aRaKAFCgcjbkn8v/92Nbvp8b
td5RKYvd9+JF9gKB3S6cjpwepovFG5BPhrJOTf9sU+f8TqpuwgwsBElfQ2UFSvmm
HWLhz7Ol9DG7eOi04KGAPhnN69YJ4BOIm5FoqV5aHjV52Elaem89KL7p51YnkcfR
aKGCdUp4mzJGRY6qGLUEfSt0J83G0Vr5u6pVdTe7m6Yxjp58Hwrq2eHgQ2U/RBT6
/NSn2pO8X/8D+3/iqmF1MEq8EVkJ7vBS9wA0WVuOlENquLGRGSNGnwmD/21vYsjb
gdKAuAG1yAg7qqKGj73J4EmcTb4OCwALPKeU6OkhgXWDPDXBGvGszCG7V2eCeG1C
eBzBYvr0fDitgiDG+mc2l1xUZnG1gHDWmBYIoKw5jmOcr1pt88WdC1ka5E5GSaj6
KI+0MECkQmKfQ73pclIWgVbb4rH41MPKPjvdXP1SxvBxMqD0+FIOoG95YAFGlSnR
rMJBrFeQl4yLDZSxOM3QaCbOyR4mfUEYFTLA093liw2m2Cam288b4atpTOPUn/dJ
Hl3lnvyUW8GtYCjsR9CI5USXCcY50GRtph7Y0aDXfY4Vi4pRNILjoAtXMzG+jPN0
mut1gTSR8BMRqBaq8Y2UHkOqMrOSWlrPPFU+KKfIXXcjsMO6j/b5xiuswRRYmhPl
pXyNb9OaCcBuDRK5otDOjluJEoIz6hqJWtLA6D0oKesh1OsnbQJyX/o9RdcO9AZd
I79HvVoJse2zDCkrhQT11FpyAUHZZyQues86n8JFH2cK+f5OfYcoxqLt2mQ0/tIm
3SEn5FdpHOzWLAvKQZTx8hnzKU0PCVQcSVh0N9O1s8/cFdEwZMb1chh+7y84t3Gs
0xMUi/2wCvrq5JjsmRqVz7Kq+X/tFfa6Bjh/trHjqqH+zytpLxsnOO99i4QEO3Ax
0alzHpE+bOOUbSA/4+3zo5rjPEAbvzDOlGkCwSMAcjcl0qU5f9EWuby3vCskrR3F
PxMsiVXYJREwe1Rx/mRvnj7NRT2RHpps8vRXMQrgG4aUtZu8/4mjQCggmczhQ3Hr
svfw/LsftIKzYqsbHlSpCnKpNAuX3YeMiKZTjQ6TDDpC5eQNySpzgAfNvHx/2QoJ
Dp4K5oaWh3e+HrKNC8dor/i3aXsCEoWDwobHNzxFBshglG4F6oXiqK0zqYUO2hDz
nortGqvN/rjWhlpMoPghDtrr3BN7I3EdyXMSb/W0AHV1GESYsy+xGChLSbUGtt/k
B+GTYr+L8nuGR4mgyaTWI3VRh5CHYNlNPuL3a2wACw92Clh1rWtRC58fk+ks83j5
VrAFjrV2hfX30KqIW1SW9E0CV9UbH3IV2bWz5QDIaytC7PJnsXAZ7llrew0tdXnt
iaKd0dS5YzZC92VcENZ84QqCl3k9+0Q/O5p1yU8VYoKTfbcJShuKAeizLYvjjbIe
tUW6TsdU1Spz2tPzCSHhWXU5JQ/3S2NlWpewp6fuo7lpNMq3v11tTRQ6VNYboxKN
HIjodZcDG6iBdnr3BzMq0H+82N45PcfC3PepnLQpU1gpmKfIJ9UkMgGmW/pFCuX6
Kx/wB6mIwJj8aLxZjQOEh0PbVkwhHsMmE6h0B6bpPejNaICnBL7lkywujRL0APxI
fdzIiXEhEpu4kD66k2ewYGwKE2bhr/Oa85A7HyuVCgBptAL45RejilxKh/LNhJGn
WRb5qyvrSZNksYVV118D0hSg9KY4ZSsgwdHwcW/hXl4DZNHOtm9Vcr1OplPnjeJs
/3z5i9ayzmkl0SSXbwOI59GBuMMkgoej9j+ktacavjxgK2qzjFoIV9WmgLmMjzVv
GUMAD8whfY5u6XkxBLCrUndPpwpOJXgvgPwKHCzA/nXZScPVL6obaQshes4dAtRm
v/JbQ+WtuQCulgTfVptvD8sg4icph4eUsxpebGzLE03+ybAaX6iqdNv9RerAojvI
IW22G/Zve6hM7JFALQGtllKBRnufjbHK1wVwpC0ig4tGiko48QXKeYG5DgQrOH+9
xt3KADSOc0t8PXSV+e4UnHAqZPGeosQBg/XGPPXIypwmYlCr5DbUXUpHI+5lnymB
ZEqg8Vah7jBEJCsdmU9Z5+1U3ZX2c90e3Ec1sQ7W+xgVJDdpADvUkFmghXwX3prT
BwrVgwEeDRdJePFNySEq6rvQuoqw/P8482EiNdxssnx61U1xYpHLQx1drxTCOW4F
rfiq+BJutvMvaR2KIIB1p9Zk/na/HhHp/b3d1myhE6STI5vb2A0PUtHDctO5kiXf
t48pGi4XEblnJpvyX0fe0c+t5eMXv4CBfQERYEZ5Y1jSPSqwMIvoPnWoRUvWDd8S
mwvVIkt/aqAnNgD93eW92ce54B6WHxqUd9Xz8CygZNFdzf0emeQJ8719k0LDaRFe
WUKSWhaAsNtQgV0vXL0s8KPcFdvO3uo74DmAWUlZ0SpJkM+BBSbXNCm0rVyZ9+uS
mdzkpa9QwsXl//HQUKZ8oPFDaYpsYt6h6W2VN35jJrwpCMeigDjC/zLI6y/kf/gG
py1zS2hS9FNCmX1gdaXUFPlOZHDQF/qpTOAzrFLmpreEq/GrKxpyKPnfg/gnMusb
ch1ln7qq53iJB99Z1ginBYHj9sS/+txvcPmAJyilrLWTDDEpYAOfMG9IJ8W17qb2
u0ab4W0p7k3DZ7hu5T9uR1OZT+6lnj+hlPjmcWmAiKQh1vEzvcT6SEPfeOik8B9A
GSE/L4+WUCWilNLMZunufq5rpwpDi67AtWwmnA35wwBViSyrQIhdguop01P7BtmL
+LzIwknNXW2Ue7uDway/LIZyhYrlHYsR+pY/61AhDIDN7aJexFH88alCnHVRAPPy
EgsU+LVp+fKHzA4E34iFE6P1T2DZvusOHM+wQUwELju0gpS3FRR5G5HIet1Em0DS
aBpCCywg0X8SCR0cMxTDvL798sRFDcG+52Wyl/PEqIqu1fZQLAqeTnf4s5Uby0GD
RU9uchikInNQMY4AJK5fP/LBiRPZ80woXMggo6tl8LuV2TlD1cJSw41mw15UrjI8
oI3g2gy3f9iE9I3banev2WYg82TE8Iotfyzeg6xaAs5vO+dUOvu1vaW6KS+bc8E+
bbaSqOQDu/DvoHTjElhuqfAd9I+zrDNegQYU1N2m6usV5A7wRtMrQPBEsV/drZdp
Zlc7gjoumRI5hYGMKbezqQOQGneOJ4cg7jAgTZJZ4WSc3MpKVqOvaMxioZETQpUR
n33IRynA1rPbwRe005HNXcio1pOgenrJtnn2VPcR2mHTJYfHk/uiRwK/83npUN3U
ahu4N6e8kTSzCgA852QfyS04qzQjfGqyIbRQBmofCjLSsoG24qmw4MWtofFkpt3y
vx9ySlta5w0COrGwp2eSREKUYxUjGC60N3h7LnaG9/hy92mCjX85sg8qDTE1I2sG
cO5SGLB7ErkA8IxvZ3FZPLQB64UtVI9IwSJjRnA1KDNzI0HnczYIBDl5wGoX+z+3
DiKAd0qlnVZcV0MnQPQhx4lEVjhVq3t2WwwqLQbPbxhIBfV0+a3iJqtZ3pjPFtOH
i5K4puTXhnLi7YI6RcOKZEHgRNF/L+rbYNwC6EG7/UenIeJQzKJ0FIICIFT38Ukj
Lht+AS2rg3dCTStjlsDYbATdsH6NB6n6ckYOz9MvYirn8b9qU9Oi6Pd63i+32Vjf
wxQZpVqO3VUDbZkchUpcuo4bmOSp2oOSaMZI0TA/uuLpRxjFLILX5isd7vmB7Un/
zRXqZ7L9Ptha8EhJ6NFznq0erZ+bcAmrqoKufkbXIbi9xfObmtjgmoFC1BmNyYJ/
/KlVx2xfIjzfnWdlnFRbE0w1Df/65OBizHG0Lrcw0y2pLqyubaBeAlv49NemTolW
7lXgHot8RJ/bcd3+F/XN3MEqULUIIN7vjWhHauyoV3UVMfsViNoUj2t9/k50uPyg
fgCxU8pe4H8HQ+jbwJZ9ZHNojbETCI1yWngNE0pqw3wmxErwJicnXUjP4e6FXEy5
WFrtOTPFDLQ5PMS5FmwD69UM4hM0piVQ888ClUb1RQTX8uGfStZ2122q5TXHNxb8
SxBbVs942qcj8X6BSIM2ujC8dUrd8uXkUf/vTLCQ7cZNpJ/LE4blJ4hFyBFgPu4c
+NmSBlCLVMP5Ut0NhMDlmVJ3oHMpCSD+Le0elC5LFBN1Ywwo/yLv5+LQBErO1mq2
9pUHmNMGsLTPGvzBW0hN1byZRJIlwa3dluZGp9LLXTkwoPhQLQpSrLQjp04+BWAi
VXg96tBD9ukYWMl9hN5Bw8strQWQe4vp1jem3foSziclPi80KAk5BTimxcZQQKUk
+/k9kgIHZJrVVj92BG2omYtSt1kvCc+DtcuQ/MmsplRr4EFhSXzWL1XHhsDGAlj+
MDAEtFshEP1JfVoW25L8r9H3q/CBaRuunXF9H/aIdqsA6nIWoPASpKCC8bSYoGe7
V1ZVZv9XrnuKUZxr2YqPvpE7jFA1adPA9GjurLtPaTEvA+e2NNXpwqeHgiO1bq2Z
0Te2X0cnVp2e0lyNO2lhlm8Nj1A4PlBLTkyR6dn1j0DW3w9P4YcTsLGnnG+iCAId
Z8rmTHsKCrS+X2VujshIID1ZktPPR9wDBdnx3arnp7VKBhz0yfMCsvAyPoQ3T3YA
fR5941yvt7CSXCGXAkhcxANQkpxNSq5SQqguTRy+MUp66RbHRFXzfwsfK4R2PruX
kOetRPjn8sDoLHD9o//KHXC5X1MIIrhCqKtKSJt+YeTkNj/REiVU+bwJUr/n/DME
8EzPVJHGMvY+vLCusqX39qNlEZQw18M1KGWgCPVK5Z5ooZoD9zN555myH2nsPflz
hJQcCn76zkjF/Tqx/2pcPehR1m3vYGrS0fZpsjs3pNiqLECOqyawVybx4nkAso6z
2cBkPPmvDG62Xg+Lca6UpLAL76t1IUwuCeOcKDd7gCZXtoPL8bjp7xJCEsN4NhUo
t1BMZkdkAGEsCswHd4lxa/rAcqA+GLN4mXgmBhncMDkF7IbNigZkzPMg3ZxO4uPB
2usVTMErIDTU/BVWzdiTTfxO30StVuYXRoGnL71LuJybrkVgjfBmUq7hMlWah2yh
VSUkSvD81HSqk7udQojIPGSeK1J6OZ8Fi/rXErH+ibHkrDMXLw+D2sfOK49U5hPg
wGeFVuTlXdB4gV1b41gxZCBQM5f6/sY5Vseggh4oUD+43M9YW9pA7YYawslxQNqP
yhtCzZ0TqrgFYfZ9upvXk9HBkKqI/UAIEx77lj8yyWWk5L/a9pAhAzsWx9IqSe0k
TCf/NhvsKXNXurqmHf0dtZ2pAKNaxaa8Tw/EHdvZWIiLWvnQD5P/6UQrMzPblQFP
dGym0jFvjAKycLsvHi4x3xWyVUxQgFD3xnHjeE39LkvPhV/sOqDk6X0ovsoaMX1E
ZHM65nWVA7GGnbsvyXyjSf4WhQdPlM6kBDSVByuiObmK3bogtihufmuZWILDlRIw
V5l03mkM53kPSSy/iflBlUryWdRnw68+/nU1uFnduHZJFG1fVW/KBclaF7FnpBpQ
tGydCfno+fewSA/TylIOGh4k7vK20Oh5p81/EpKM2sCD6ssgXlvICP9DTJ5KTjdE
9wzmn/sGa3VmWrZZfXZsAZ3HU9aVFkGgdom766gLRr7oPnKQesUwFfFQ+sDIQ4sO
jjHOv0LMxKqPktWp088+aKiXbDARx8ljPCud6m3t12tZBznh5PqqcIHZwBCaosXu
wTnO795gv8na4Rb4f9Vzi+dZ5+LFUeT4ZVF+J3ygpGoUg0EHMIEdHygRX6P00wkY
F0ovqDGP57KKIf2kQz62Nv1DVqKIQJF0Tc/w11AyhDWW3Fotp+JtIvnL9KuQPJ1M
uWLUNYpUDiucEaOMHa521gYIqOPZmbJEnjppiJt/b22KtTKJNwbDylrmIuDdI2kE
bQYKT/7pELlvYvULzeYdEAv9KWnEMxtJJanV/UuNkhJzCFK89vQITrSvJhyx45Ay
zWUUGf5sfvlZvrDC79+hzF6kjpRM+j14W1XsvsW4F8Vc2SV0qWn9aYPaDYdjstFF
U6IPxueREYOHaShbnEd6Sq3vNvztX8emeXnqKWkERnowzUiVRzWG9KqtKZMrj4Y7
gDMDs2ZVYBxPJSBdrty+E+Tt2vSM2uBYsFs0l5cuXElGvFSOMdV6SxsAtSx20in0
cCOsahrvaEcQZO1P/BoP6IOpQ7OwHBJ8rl6dEW9OC+nC67Xzm8sNBUY+u/hlxAgi
LPOWWsK+dMgqK2s+aIMIrHGmUpLc+Uu60xBER7cdKa8b5039UDH+xIahEiPiAfou
dWZg1zvi9+gDHb1RKKyF2WClsdSwU8pk7Lgap4vwjDX7uCknfoJjguUHsR04sw/G
d/ETgj3G6n0OZsbmJN5CtFLWcCTs5obPknRF4PA1F/Wb+KAvkLBT3DSxS07G0FVH
vQMpcB9RTrIiT+XgdiRh/L1SnX0BKc2oziNqgHWX9XyVpkzObIFHOYKWqNtZfaqQ
E9Z7E00dUaiFGirN8/U7AjWmSfH8tMmLKF3U3qNFo3R9e6vhofYB1StjFsklCHhn
OabdcfcHZ/KArCb4NsUAjx2fvOAvLCS2Fkc5hJoaJaSTfCeaxikEm70MUC8ftIlz
ENtiF1A1r8CNhTbtkJAwGZnwNvib3obGUztTj5Uf7HrcDy5G2tvfG6gxh+nGlGHc
wCvFq6f4+mPhQNE4M30VaLERBWOR+MIWnFK2sji+9xix0iZtklEY5/9/6zzLlmI/
B14hfqYzvabJm8dnpcSWnJAjCkjYwSJS062cd0g0w46kzZCLzttuem9MHyAiqCDz
HTrsi/NjzfL6gR/uHyPvd6HBC4Fidzw/ytO1Ez1UhughIYWYQx0Bf4TOYOfAYHub
IdcOhiVUJ6/+rxNx52dpraw8kKknTbqWKVDneAdKXp8UcGMt7DxhhnsyNR9UBonZ
ku238UkLY4IEfFaf7CfXV+ooG8yvUPrS8DfjpqaUDS/dtn0OFZbSsL/Qg7e2wrNW
PakGgkz6DP2/TJjQNHxgFJMvmz8N8K/Wdl+BGJJkkFVxQdyyhcBN2PhmK5S6Z57K
EtJYFTDd/Gi2bjAgvAPMFZMQJdlPW+UFkFYMvNRJPbo8rkGv0oUVhbD3/F6rWQ2q
gsWkklOCWIiBegdUPn/RkkFlZR+6NCH+YXYftGpRDKjKFmlAei3jR2rr104513wj
JttaLSTMdkFVMP5FphzHy0HWvhkKgTmMcfWMZcRlMIJnYVDo9Q8fC2ZioxHAnh6O
IqLOwnVRRwt2VFnllcstBaYxmULhkoV5NU47/dcc8n8boZgZ66wJXpp7NHqZxNyH
BLHqxklwm9itPaIq1YVrKpExNVXOBCh9oVl+lz5Sg/LVJFwNFEbBbyDLQ8pF7pKs
LFDkuZXDhaC4pUdWkNzrYNBqAkLy4R6SyPGWXav2pcbk4lcLtqQaDHoV2Gn4qQzb
NapDMK2A33DlQRcci+Guf5giDgHevzrQNPd0SS+L5xvIORhutfuLGf7tyI4uyGF1
xPQlydIrghqg9YQY3LBnCwqkkmKQyU3vNOEEQorvVzHRcAm2r4MkXFQl+bkygLUa
JHfv86bf0g5RwOZdtRQjAJfZ/31L7pTCcRTnOpE9U1RT3A8xW0kUOChbzxn8yxt4
DqUFkq9v0jHmriaP6qxYrP66sLIhUIfzNFxgKFbKQE1xbW6OUAkgYUxtWRc8e0YY
oFRtxGPfW6S4oy2rkNvP+dEqBmrofxkRyF3EfMrd9rgriKCjeg+cwHCAhjdlTwVj
0qG0ifm/vrLkoUp1U3RDcWVDwv9QPYbG68u8w5XZYhFaRUg+s/wV4kizwwnMe0YV
/PUPwgoZMiZ9WpWd5niaJR2Jw9KdiCOzf0xFPwfDOkH7uJaD5IuhkM862XOXAYtu
JyRsIGq+iYV3dBeE8AMl7oTK4M+Dz0n3sLhOALs1Qq2Zg1IXhlnFqUMWthkd7XKq
MTeAmm05qzmMCRrMsMmQNiwZKL90+EkUUVns2wXP88J0ZDL5pfNbt873x9EYnOB7
+VL12MPuao0GSh0XKXsRxZZFk+6taZA96Q27ivAEdWEWFdNzlw3aKru06umQF/rW
zrSpA2orBHYiKbo2IQKBu933t/r6qe7j65KRtRakP71i1fPZJFXAAngKo16aiyMU
zaVeuECYcxqhE6a90Zy684PrOOx6YFbndUK8Na/a1f3YJqUaRfCfa8h43o1U/Olx
sODOFu84VAFHLNSy9TJLf7oSlLungiJA9NbkJEK/Brbtxa7TeTKZkXiHdUSP/UUV
CX4a8+Wu842ZRy3aYo04QCpLZ2xpxeDeHFw44ZFS/U5Inkki7ItIsAVKK26L6iis
72wwtk6/nxWyP/spNP27lGHTcvSR4e71USIN4Kro54JgosJuuWYvm+nym9Jg/lVP
6dR4y5Mx0cVw99yY/stJinRXOce/nb3+pOn1MsBygXxMsAGtM/vvZPOVB3y+CGa6
UWTnetzZpCiJoMDxkzQEzFBDcF2ZKBTwitiJ3rSCdjzvZiKnM34HihUdK8lV7APU
xOGnHSk7/52w8hi5I69KRxdCVX8+aXjkhyvd0Gln7xZn6Y111P3z/2CgrTJZnU79
qEnTquRBBBxVabYyvNy5iwzqBmLAFH1MELYds4u50XX9Trnc+dGo76Y4VsGwdjwI
Co1U1MfeEuZOGGYYL2+m3sabVpDcgWkEqIYf2ca1xhDi9InXsqwv1B1H8PlbnZd3
Y7feSfre3LWvJxCTPtqotwfY3euiNHJn4rVDLLZi5sYLrVQfY7qda9CgocbstjE9
1rN55f7Xool5WLKWYZpTiLipMboq+JfdzQH6kfSXX72Nu/gq7+nn6AzPX2lr4bEd
IW9wxnL0w5gcZFWumzJthquDE91zWQTSI/PjXkfeQcSRMqUxaaf+W4V1q7DTi/7K
4zp4aGwUaD9ncSLkNTb6HiYr2aFrQ2NaOrdiuspSLXDqwulFPdgEATvjGDhp7D/e
utpjG/1JQCO/N+9Udc3gUr2gnnJN/T2UNQ/YKiYqBzf49k14h5/QrVL/6BLITNSe
wFZSioERJ0ogK/1nTX6IltY8P89oMHpmIUzi+tM0IW1BWM86KjXG/8XeCDfDy1Dj
mBolcyDx8tIPrwzpFXqqVYbBV+Y1A7uMBIuDaaicdz0rznLDVz7yOg9Kc1Ky8v0t
AmBs6/qFOlXbOGNrCNmzqsIX/jPZyzcfRxa3gicIoagf+M24GHAsow3bEaGaAtsg
A+sPSbFMR0/1wGY7ctNbTprRzPzoB5n1Ka2ZVZ1pbkgX7MzeelmFBduuObDzMOuf
5Da1Uua88m5BSuGU2hMoru64MgTXtPPPsXCtpD7+emrbOkpUqFc+ew0ApfFgqtNb
gMIoUPlJFRd5t1YyI+BKl9YIhhaFysZK+srjHp4HHPkMNczVBqE2t99IqGWoX5P9
C8bvC7Tlhcav1zHT0jyEZXOXQYs4gbw9AA3uoytvM3qX5lkugmllgjlJw37xjicr
KrUZPDVwZXwhlSjWNZHM3Zanx9pkk7xHccrGVFb0cpr8mu9bcJCcnO71X+ayaJn/
wVmMrwxmZxtm4bJCdM/wRJrpvM5p+0qSgCNZo04WyFUfCaJslHCfEmedTcqs7LtM
K7rn6iwhe0JE0SLfbsI1VRxXYUpZfnpKfXDTuu0alddOj+tk/9rZQ6jKDd6khYJl
Rxscx14yElNkpU8XodVeSjDKZQzdbSBIlhd83FI/Qi2NqozgUkGFiPhJFSmfbrng
Way+YXKccZBjtFhQsRGuLYine6mo8Jh37OpWvBRliymw8rl+IlAkPd+kLtAmIeMH
pdBgS/oPYYpw62YbmzD1QtZzLi/2cIi6kFS/e3Jp3huH526M3FmPxG7//CZNtRnt
oVqN9lzC3SDg15BUxRTnJobi+K8IhxKPLpnf/KKwj6Z+LZ/SCasEcixgNG2bSQq6
nozVuL7GlajwpMZPujOCJz6rFN0VnGI4BesL1bZSC25cgt1C0jzv1wubjBWTJwZt
kC8F73LgVb7CETBxx0Mikc0rxCMj9RsIq/K+SniZdLkATvpElPkTDstrGLmrC1B/
LooZkhWHNEt+dCslvuIMY0GEsZBC0Z0togj9INKwltKCB6BGM2TaoFMrxMgoK+nZ
KYu5sGlMrDJ9qr4dGcmyg81Ascb7tnhMXV/rHJXH1nTf/lmYppc71hz46RWak2WG
pDTJFJO5TeNGcx/4ktZHLbczBZOJF+gnWN6kzp/zhoVIXN61Ihe8MVqjuZ6VRxnQ
f7h+1l3FvsfwOOGTmp1ety+Q4LamTnSBENbCRkPlNLS7+pUQRuZD7gsuyW5Jfo9+
4upnESfHsp7MunB8FvzMc0XasoMclEEVNuB8XPjz28dMxFoRQPeJo0svSNeIViuh
bY1gBUVFlccdrLLAONc6/TsarPXcmA29Fb9sk/6AUOz/g7fG/8btTGo2VRTXsEi6
brfwRIuuoky8pkqsYAkLMiZenIYxT6HLedJJbtFir+IFR1knEELu0fh5R6PVE/tH
sLF23R4yd9xLha2a7QPLkuRHYwNuS8ipI4k+cpeRMQpmp1UrapIq0XHOfkigus/y
K6Rp+2Ga7cd9E3kg3HTxNxV/HXbzTss9yEswQ5Tvs5TeXdM5CiHjTMuZnqMdSi1X
+9ByYtOUsw+RYOwnsY4Cjv733mg6yYIvgErgNl3c+bFnAExDpw4qrP+G0DGP9Q7h
P0XXL1rBy2iMRJ1FMMjKzIKo2CdqNxlLEeFbimxvrGiGEGrnPqPuxxk6QgyDgoNi
jmrtMHJPmQfSe2/M/JXiJEGkPIbdTfjPIQA48+ZvgJ1H4NPWK9ULrw/6wfAgFweU
cj++ymk8dOpbubalo+R/iF1gqFmf7Ga/haKkHiJkvWcN1ZjrDCG0BoMyF80i2jGV
F3BhrxCp3U17FAQ+7aU7GHNwgs/a9KGGf95aKjvi1Xo7G5uQyjuaQWYOg4gBZ3Lg
2Yd3aOSXza6mBb20fkROxg02Z0E5qH3ukqXg1wratFq+/u7/B3x4lp3q5QLaJh1R
0ecB48N+RO2rHS6qAO+EYPo2/dPxSoxJPxYb5ri6POPsL/4ox3doerdI2eBZjimw
7s0stq+p+hRNzEW0qKL0cIzlWSdbG+knzkgGeoBeAgbIPaxVU9RJRo+lwERm/4jL
Zm4H8McE+Bx/Oj6vZdgjfYR7g0qm/iyRLSKSgrk+s0PfuiMf7uXGcH6wYL47Ime9
yWqkLoe4T8mmS0N49ovxe1Rsll4WlINeVlufcpZEx6UGfya/FkpoY6m/5aZCmkXI
kgucl2yL3Pe04WjXWrP8dQgzLZ8QfwZc7rlRXtARxh6PgZ256aLt3dGzSGiJx24M
MjKimg03EuUyQzTExY5h3bN7qxdb3Ekedl65j2wiO4YlvnFWVHHA/r1hOIAMAhL1
Otp7tFDjvG+6NI45hCcW9X0Nh34ZHw+NQUJAr/ug15dZS2WRGQrxyAHLGuJ04zyU
+cVXXworwgLXfiZuBcF4qGtcwxl2xfob47LUxcqWzpQo3qB0PTfN6C5ku8SuOjwt
EE08Wv6qKiG+Le1ocehdJ6aytEksBWM7K2ppJRNLJ+bm3IKvv8hFuc+75Kf7wPIy
+BGVLQ5fIOhw1uUYw6gM04RmjCAA17jUejvZO3U2tBxiQnRIi5CMvAADJjdRhlgr
35mIAqdxRsCBPjwIjodGT67WkGupuIzdz1h4VkPz4SI+LiR+MT79ZMGM9YalsBbF
JAfVOd/bLZQRBIm+Y+IpHDEpwfatqqTBMLkmjK0Ub7nRp+kJy7SXQsIA26dyhHm3
iudM6F7+x4YkDsZL8zmsyujznVL7K2Vanukq3sCvTvyP+/8Wsym+RFfYHf/WlKrk
mJRRkjtZpweZmi7WdDClXo2RuxynNXirnDf7U9dSgMul250WwSHRcTdKh1Omc8cK
PZQT8ch9BVX0uCZ0p3o7TWfNjKrCTWzzDjwLAPQvol2qaVQUzMA+n7AtNIQsNcA9
3Mkakzjns0uVW5H8VO3qzMRnTzKpdcTemZZ/4IKcxejBwv8x69JMeLUKp+pLavqm
hhfvP59tpT/J9OaKrouOqYiKF5aIJaRShp/A0enI7jSPhwu4TVf/3REd7L4x9Snf
obiWzzCzeFNS0luXjTz+hJIpUdvVykJByXrzu2hc6EjEvv2rzV3mU9mk44EVhWa2
PQUTqsRI5AZd1YC+wtTibrb0kzNJtAd2UkC/aBg8k7c2zio9Ex9z0YAqeo65Wl5F
YE95N0ig1yxhA0jCr9Rtwvo6Ljd3QnSNkzR302Re5OvkUvecartDGWVMNiAqEGem
76t4jKQfPvpuikHuGAIG5IeS+Zp7PQgcHLLcfBn5Dw+WwKqvytxpJt5xkAdT3xT9
pPMm9L4dPT3Zx7P6dDQc0Uvcf+cTGypp17MSsjV5pB8AYzRhRJCoV7BCXgYZ5qss
vPmD5mSWpiadM21ernDhxWfs36s9UOFsJBEN9Frw4j6C1hI4+DTh/7FcwQQNFuAO
bf1SMfRGaqlHZu4+xkfngwskxVEshysjEaaV+SPuiix3UEs2b99banYHkx84NHRe
MUP36vC7nlpbXk4mzp98DctBAtBojaf9t9QKLoPKRdspS6JUebwIBmxzlX/zIzUo
aPbQyF/OHhe/WZIlBfQ3A7igEcvTvCpjz342e/DdNvnKw9rpWjArqS8boVP5zm3P
zG2Da7DsyPglSgX+7jnfLX55hO+gs56Be8pcyo5UqboAwZodfR26Iw1RaAL5qr78
muT9KqJ/SrgBf4BfVST46UnBIFZpPkyY/MGPSxEp8ToAZAM6jYaGHcD0GyM/Tn2i
vM+XVRMtzkJxeEyfppeBo/iCZ6vucDcq+85+A3ton0Z49F/Nc7DIKmKSiV2DgajB
7BClNjfxvfSgYYDL6EtLeX5SF0Ey2t/b/Bs/ySG75s5Sv+SX/K9xk2g9OQrtQ0To
dn3kblThchJCJyQ/H5B31fBBqjWN+hemfuX1E5k/X3QbctJc+QRe2Fd6BBfSF41F
SjmseMI2srQAZr4+YC5baXqOj/eQVdFUjB1M1l+NuJmulGWByaziSqvWNNIz2Efm
hT1aXuG1Arlou1s8fhFux09kZFIMa5g7Jaj7UEAZbAY9qV9EDcHClsZwMfbAMmK7
1eDEYki8BysAkWtOs3E+u8QF04sRFFJlVYBxtb3e4oTzHFKNCz/M9aIjRN5XeLMT
SAaMIEQgaP50eFUDhxYEtoS/ojW497Iv8jIZhwK+LhHgkeBVtLUxMRp4GI5rSLfq
783XQwTTFeehPaDe0sz3a57rK9C/wvpDoGzxJRoPE2jXH78TlQfWvlZO4hdymivD
ndmSzLNRpTq4WeE6xncieA1GemfwwC6hVml3y/c7GKT9iw507bCzU+VBnnUag01S
hmKpNJd2n39OtpEB3SLob4jMXeoukgOcGf0RbyMnhlZ/YQaZ2GkxaYQQZHFztn01
OUGJL90xYtz2CkaMMVDQz4mkJePwRXDzJxy5b+LItv/QgVzw4eko8S/9Tj2QvWR7
F+iTKomq03ThnDU9YddRwIsCnbVIZorXkxqEg9D+DAm5e7y/tn+EiaXCLKRJmWNw
xEe+JK5MQOhv/NF34KLbQCeBsmCNjMZ8KHK7PUOTr953N2u9mKYWZXnw/3KW2+6/
BdySl9AAq6+l10XvOpyN1ZKTmTcgdHf4jmS1gTVZMudL4T3m6Xn68sXj+JX9ZNbH
K+1DxcjXO6QYf6bAZjiOYi+U9tflMblLRzGbh5JavexwllfLLFcU2ZHjV2lxSBJF
4dvo0LntLeiJ2ZQ8C4zMAdzP1u77+dThgMsdQPHt4QNoQUMeL/KF2UXQ7khwXjur
IzFdrIWYC5ciJSXTjqq+z+k79Ntok98dAcCoUnYc9MRcl+9OZwLUfn3liBi81D3n
6IqYQ11J3iPP9I/7X66Fs0hhDXoc5PI4lTixaBTZXpMifNc6iVT+RM2uENkAjpzO
MLs9mBrUSH9378V+i/JREPAN0rWiTkxPk0UU2JsxE+1lSm7VsEJwapaTJcyRISBa
op0w0/7o37ZqhC3L4LwoK3vosSUAKm0gxAZnERTFJbV59h3mNwggbHTFjaC4s/bD
cbmv5KZDaT0G194JWxiIN8QdLdnFbX6JVNNm8WSA7MksAcKquskzGnRocgkJxXX9
um3NJCuLZ68GE4B0jHQP0+SkDUJkf1R1WPfkh/vjv/Glns0x65RwL7S0JKGRNfTq
7rm8pllIviq+FqPtS59b51KbqeFcBwbl3vHzCv5kT+W0AbUA03Sk8LTEDZ6NoMyS
is8bTXqMu8t5Jtbs0GmNqfZoiK0C/joFE+5WWZQEL5rrC5Z+p42PRArBbwU5BIUB
Z14yxP4YWffhGtSgHisUmqfIUjfA8SXLAl0hKDZUQi8wXOU9o5UumANxuGnBynNp
tJfCWAwKpMXj7uP7ckalr4cN9qtrQd07+7j/Uv/U+iaCFEXD0ZOx+FqZSdEC/2rJ
3r08FbxokhzRAUZR7fntHeqTR7VLp4CBvm1xVGTQ/zonoJIXRFzcbtqfHx7HX7R/
dwyg2+hlZOlhgwGmgFjfBWsnFzT9eHU61X+l41eXhDLevEsJppN2gxelqFjwfq8w
f7/5HARGbjrgtNtkbtZ24osBLJMUmHaX1dg1OqidjwY9nVGVgJfXHAp2L1rOJqti
D4ENdE9/nQyP0+ASl2gM2UqE9v1YQxRM6OwIfdMd4J9qLCRj2R5y5O+N7gWItuOW
j7VZBE9qgEcR0SjkjO6J8ChVHD3WXM7KlnP9SlyAixyZ6IHUE08fFqotySrh/i2O
72E8SL7gdziQKKp8mg7wKlHRHQzWIkzdBh4dcNskAzGqMnBGqNBcKll7dUOHAIHO
DM227UrbTS+emR1MauFgMgzD0fttB4doswHW/q3RynUUGOsYMh3XDFF54fY4DVlU
lZb2nhoADnHPZd/7jbc8G6rcMIapyPiGEpndd2ii5sr4Katu3qK+JxC8cPscd44R
Cut0VgVLoMl3aUHcwTE/CrR2gxgecjzz3rTD6nxteXJfuyEi48gSbqe+NYDW61M6
xf32Gx+swvPQ6QflpMPOPs0euT6en+nv/1x/9QWwAhKfGr5qBQiSuYmPqy2DLlfi
56LBPWf6RccEKUk8VAHlmlrHnZ+hYJTV3bgt9+C9p2nUFxuOUZmfzeWFT2fZD/6k
3tcmUzAgdzgI+/GJ8OA96/VAgffyIjBK8570rW1IkvZZAqaBUSm3vWQphu4vbHMR
Vqo0QT+q7dnQFdEra6AbjeCXkQhf2o+UHv1VmDzMo2luAlVSh89eg+wW8F8X5RUS
ZjmgcW1UhJJoyRVgDlBozvPKMmT/FJGfN75Jzq2OdihUaq7wI0jarx7yTspd2Vfy
LU7Vjz68jgEPNALXMKLqSlrB1XGCQn8Qfg5pabdwSXpNtJ0Hlj9F/l2hBOtYMvvO
pdCeekqyWeswu/yXTuJY9AAv3wIWqutDJvzDic88ZtEks4eDZzxmtPmPf4K94FZn
AlHZT4e+4AeWkurA31DBM+JaiQ5WDZLJjVonJbdHtmN0GklCTxm1YBFpZ2ZoZzvV
MBBP70qvw96FSv5rgEe4KG5Lri+J4ddu7wWS2vtO9rtJKOCdywo8h6mBNs7o4jc9
f6xluBXfD8XMI9fEDL9SU9RZTdO9f2+5xrXjhBrW+jmXYztss82qZx4gD1uG9wKo
kuwPzfrTKsADtA+QYTvYw4N16QP0FaH9Plf56kfOo+mT0P3yeb5hjXRI2ejgh5LN
xGVYgyXIlMTQ538/vEg5+suFAdiHzZMzOZLII9E+krqxGulCyDngUL5rST3xwfEe
iIFTjTo8vTMw8MtBWAJuVaM8gX7I9KjRjvfPJQeXPzTdgd7pa+3f2ITHKkJSXUI8
zSLalHR6DpAOWbTCtIk8jTVDWtyrxKQEAouRFiptGIv/5eYkKTWc9pPIP1yiaXyj
uzhyJNv7qv7RajYPDq71UV2QJSQQIBhzsa94zFHINoOyRZK+e4wf89ckqoNkoan3
0HNvlVw14PV+/WeDGClok8fyTwEQG3zzqIavdi6QJWZtuEf+dBQh4BiKyDigqb5p
mIfQYkj499ASv8d7ZaxEXKkrsAvZihBD6BDaCItKKnxWzvWPeJxYuyhYOJW7Wyox
JV14C5vokdXD3qcqOU1T4J/ympoe5pOWl7KiKqf+2Lq10zRtuHR/PT4/PrIcg1NE
Z9bVlkC3u+4BKH6ncX+vxsR+fU27hrElVVHqTzA3wDwg7Q1bv5sFu3QtKvqsoIpW
7TAklhNimou9UDtkOjWVAMLbbn80vb7fegzhTouCr7NSXAzVaMi9mDrGi4SUs/u8
mwqHi5EKfYnocYw8SXHNrbTRBmNIURe1PE5S5c09E7Gj1H4s97R+m2oE6QeabFt9
J2egiPh+D9YTZ3bz+43Gi7oyAg/hqGJlEs1j0SZjgJ8NVEh0V2JhI0Dc6CDXGYfM
JAmpk5oXVgNZTO0/lzbPTXkl8fgaUxlHqK90zz+gDgkt1r9q1iF5loV6EkwsF7rF
eXasCPgmkIHAGcuP7ipxUarOZJOAIEYCLvdiXKFtTsqxLCCesCRjCS+YMrsLDVna
JUWuePbssjSn6aGHw119tJONnIzUHjwJbQ2sJqrv3Yyx/tlsW8OnaMvzPtYQRYj/
Q6DyHGwURV+Q9NoZ9FkOcRuWl6RH/0jeqaj+lbqBISuS9s+3gZdi1ETDtL5zT2HY
RN96yj7PzUrKtINBfviYIP1SXSpYa4MGNTF1za/NfPnKU81OGZKYn40Kll5c8+0p
jA8cpiB0bLNmN1qvRkURhn+JSWbk3zX3PssxaYbtxGuDpJyXVugz5OXWJDxEuCyM
LEfEdOjYuG81oSBITPbRR+HCxPixSVKZ29NhXnJ25U9Dqp9oXLixWd0HBHk49yNl
YfocpK/SugN1JxrKYDjZ+Jn6/kKVW8b/o7y6GXQoBwyJlPTB1oqj0gWQczi2eHww
6XgHEhkfm6h44cwo9T+8VdnK/GFUYLEm8nv7YKJ6sqMKP9bZSwUKSGs27PH67UPe
UrmUKB39xVcoPjuM9LYgYRGWmGvX6ibXLR34z/KtxwljJHGp57jisyCs2vGarjhH
wAooH7PZpRWfg4EaSLgcM6TLeQSIxSv+ToEEogpX7OvtBQl3IQ/K2/a235qhjxSZ
mN7FFjzcodSNp0wgm05iK5sZ9mh7xyEtDqTBovMcJa3FAuPePHiwdyaEujBOJ6Rd
K4gMPLVbmR99vnxSEnlvmdYUXVfyCzDwrT4rW7wIrq6jk2HpVFiSz0NU41aB3ytX
P1DMFkQhcfz4oZAO6LWypL6Uz1ChRMVBdpleQmWXXqvRzFFIhS80oSaNIyL8Vqg9
qEzoo+VakjJ/e4iqVMFZ2drpBOmB6/ZweMszVMXMfQte6VuFE0iNQ/vkTo7TKT1/
9wnuq32M27tSMhfjjT6RSK8ueuqo9iSPBTmbaRXiM8njJGWiyiWVnCR+/jihROrB
rWxuSu+T3Fe3PpjEFWFYCeENr38E+xUQtyLXLvnMARCjIDFZXHG5eMvt6Z3ctvTD
kFycpM++w5krgd+oVq4u33g91eHrVFGd2STIL39cf1eJegQUF0eGIrHdLV035mPW
1MORCMPq2wyVx7bJAhFEhwbDs1GIBq1M+SJQQtNhq61HV6PBA3HtydrUGwZSWCsG
5J8AY5JdU9Xhj56RQMLi2miWCvwKyp2A8xt9nzR6SNoVpQ0RqKphav/DMfVxXtoH
60JJ54OZlKKZjreytUVoq6i4x/sqJv3pNhzNapwv7wsVztrbpOKZHhuBMDX+GsdK
F59e8OSXNkHtJNJU7Zd0/YjBfd6xfDvmECNxGMr/1nFlPtIrZZ+eyOk8WrOSZVlX
h1oEbK2shGSHR/lV+EtoP1RQq4JMRPZqeaFE3o0f3dxRoFhrLtq31hT3JKOTemX3
awNQQj9OuH7iW/j9hGoGbWA+p5+6cvm03YTY7iSF57w0DVndA1MvMOiP5V2dqvHW
Z3tJH1amDWi0GvtIccJZJQ2glc3lLEmntx0uUpI5LiL0O0kkdTPtq1CLYyG1Q0K3
z6Zqd/Ilt1UJgz278Mn+x1KxVSABYZ/o9kqErv6WaM+QnOkDAVwDw9Rp7GdQCr7S
S1kOe53OC9ia+FuJuWIeQiES7rOlRc/8xGxfG2MB3pJCXWLg2ePk3UwIMF7aztjh
kaPElAS///hk16C4ygZeYU9A5TJyw3eY9bL5scIOh7lyhIW1LaO6eeJq66LVmwqu
4aJkX9S/cVpqi8rGApdTiMkzXS2XcGq5KzcWFdPdNxyVsPtjaPIxfmeKnVgrCkMY
i6brO61ypDC3NvUaEotZ2x/f6gG01kQsQpuRA51SEnbejb+GdwR1R0NCkjSwXtXs
HDC1Yl8RNAxIRMSk4CCZrw4YB5LKuIhmhY3sGmDXPRR3o7PoOr/jZduJUZYKvHBq
BJ8w2wPZ5CMPJ6kURW2wGSX/vY2DU7K0qmOjpZ1pzwzJeCii705q8yswv9mVKfvg
wylOfivcGizDAGLvhx10yYksQvQmhA5OYNBChgbL4+cZeHERKk5DGWrLbXE+YZ+I
ehpeoiAZk2ik2MGwWgAwT4EnMHS7ORw6Vu9A3TcZRsWAyAfCILf+mAy8Ti7HmuZe
6gqnN/wXIytPCazRZHoxPINXzhM/+Vwn/gM/VM5An1TK1ckC02l3u26186+DIZbI
DAiK5TcXBNElJDOj+gn1kn9S3sGoGLWRgV8NN7ax4t17yqd4HRJbkTH104ZdB9o+
xEuQ8TuFmr+Z9dBAF66kqns73TYzoL3pcwtoKf45TIDDEAPvf+vUjNIU3YYNV70r
6+UuZ/doBWotePsOzjRIkSoVRfrkuBZYaYMgI32zbRfzE6xqHO6NTaRDuyD+e6xz
FD+KJKrXEVES3ZLRXkV78tEXmFMOJ/kYnm3LjJmclBKtpvfnWYIVy76LhJczm2MY
qd9AVaqnJFM9AgOXeq+Qb5REmmFdqFpca/J/qYUzLvA5UzKAzvF+T1uc4mteuCQc
UYZYmQZ0arE62Wl/+7zOwITeU9pmHjzGHrqbQNNqBNAuWIo2hnLIlFrd6VqxzUW9
jqTCEES2cbw6P2UvgvXUEr8EovvmpI6q2KEG5Dzeh9wQreMA1xbCGp6FxFnHNLFt
WEl4AvbKCFaASM0bz6vc7fEGG9naGc9mYcvC1D/3JakKpwl4CC2xsamRSTvKMtQC
Z3nhvputr9TB3xKdBT6gBBnUIuGBV7eEcQ4oQS6v27hOP/8yeu9D9AI2sv08JhAP
FE9kKympSxpH6rS0+nRJTA09RuYCaJpy7SxnORMqLb+1ctNo5WNZc5gqJErxxWFa
C0C1BdduLVb96NiQHgxftDgnNsp4M1JzHpBB0dH0Duh0n5m/06sjDfx0BRJ5aJ6n
Yz4RLF1XiDkDUE9HWGukmCPp0zt8GyTzI633CagPu+1bG0q+MWU7ZDvVuXglQbc3
6logHuXmDBO9nWU+8XM2aWFjT8UnL4SNxesAtCdR9EfkVP0lolerceTzSxbnJH+o
C5lsw3R7cwiJlBaDQLMcgYl7pKAtkhdajFWx/hsoreFm1v2AHDOVdxH3QPBl6thr
K1ww/lJKaYs3vzNbHPf/3T59+Qd5wJcrUhYKEMrp/9RZtwaWp+1orUWBAU4DCZex
m0iRt76liRjHerKahE9uM6kftWfaXX3Y8DeHBNGUOQPlsGNMbG4PKQ6W3vAsuKLv
t4984WCIfmHuU6RP9tSzvnLcEDOxD2br3JeRiEPo07ay/xsjT5wb7Q4TRf5+/l29
MGlkd13tOUy68m5E9NwClLzDLDeZUDSRMExdr2kbVa1CkA+OBoPigB48OKoIEaBs
QxfrAnCSIJnVtrG0EBBTzFH0gFoYHUgJ3v/cgB6WuormMUts97s6Vtj4EkMVWJKc
i5CiLN4I3TExRaPUjS23FWVOuTTcaptUsed2K3qW7bvNbLK4bEmKR1Emcz16Fsg7
c4CLHnRsApUYFiv749orQP56etdbBe9D6odJfP7/e90EUuGRiL8YxacY52I/jqMw
gYyR+gMvke1DpHpWV2HwQJqnc2d+WEgzX6F+6uQlXcoYAAobnQCqMYCd9bGTTohR
pnAHAJz06POcsD8VJPWbEPVJciotMNe87mYiZ/HjTZam5yHXDVBhxELzLw9nM9he
yIS/yglnmU5INgeVTKwFtUhXBlN/WN8gN0/RkGiZyzsqnMcoAT88Rj+ADbOFvhEc
FQuzieY8wy49D8CbLjhDkAgg2FyeaA9xU92Mrt9V7jy3CC61iJ7Fa9iyCDkW4YLA
47ram+eTtXk1Mzd2ssvREkY3VKmsNOsEjUvg8vlBvuooyDv6kOTP0oQzuhhZsd10
um3jMzvAfQA+j3+UYamhdRJVvvAModsmP/Ilr9Mg7NaZKV7+MWFj28IxI3kFQ2rH
zKzHhpgUPP3simUq3r/RHNAM+J63lvoyjlDoocN74GY6fTYXKkCIIzhMnUfGxkLj
WLhCZ20FlZVqWWgr7cKAjamRTr8Nm2jMKyF/qTziGHatsXj8RXvUzUnH+WlUV3/2
CaMORuHFVEkcSmRZ/i1Dfz9qejL+grNy2H1EEnt2peSJgP0x4pjLtqeR1KrG3BL+
/aG+RVu1mtuKpXoxmkZsiKwLWIRwim5wmQMh6hwzcoXOaE5xxBhNWRlM1ClpldlA
88mR2bpJp7jVAMu8n4qoTkwfFsc9M97j/IpTi+NX0NIv2u2NVD++DXI8akg+uoKG
el+uiI7cmfzZf3Y38TepnAED5iSQbcB4Isi488ZuC9je252CVHuGfsnZfLpY5EoJ
QbiTwkxY373u9iy/iLbrcW42r9gztGc4weYxFO2mhMqPdQbnpvDmvVZBr+C9d5JC
dpChR8kR9Yq+d0WRbLtHL+ljVqwvOH89r4avOS2poMN9EO6RkFn5lHX7zCsdnKDZ
Ve2CUqUB8/8uCKDhA6YkHjcqHdd3/fMWid1ZXAVJhFiRrf+paZof9KNSTqdzbF2s
fhGhsQ4zMDNRFgDLL1YfGB16l7kaiw2fJRTEKRfBI8eJ3LudWQGOwzYaaiAZHh1G
AaeOqi88zvHybsZiaYVv1trO+SQ6g8fs8eDOb5HcaYWEVYzyWL7MxzFhKHDcc8Sn
mYxmt+jM0sgE7lu3SyePTGehVnl6XV7YgbJb+9IYpZYg+GsXchTJplGTfHQ4dl6I
Rh2HOn5AD4ibd+d+KKEuNdO2x1YmMhaXtdkFAF08qJ2IUsmXFVDeyEvyrPZSQf3I
4iyuLxK8PbD+DqspPgSIIklPruU6eWywiMNJc6rzk247gdDjrYJIKBEBwgGFyv8N
IijQo4i2EMuRUk1hJ0eOXkJxWMe/jKJj4ykxkVUYEC5ngIeDR+NVqEYXB8ZLsEwG
DQ5+0HizV0MuOVk3TKKBLn7f4YTLOqqSCQIUAc+fMc79uaZYwVu5nNFZRjFQmI1Y
IrCe3EzDIhhmzn1SXbwWGJPRVaq6gS2cYg0z1zAHVoCliLnc79gXfh06Bg0rxv7u
uOcgigTntKhKLpoM/U4lQ9q+lKoQdr2SlsZrgmb4/0sbX+z4xGB0HQMNl/We8yaV
j7M/yEX4FObwsXeqKe7elqD7dsROYFEPSIUTXzm7+R7MKl5lclgCFqdf675K7fxJ
zl/ujOMHo6m77ZyvEC6Xzx2pW1ZKhY3Nt4IiqNqHF1YyX0YYV/NlK7QsHqceiIJl
LXVvnCfUkpnOOyVMMW315nMUtxJmyJdLSjGI6u689C8FUkgSQptlKNUn/mydsNr2
w+kNHeGgBeEdcgBAr816oeLuAnDePbV2i/LxQF/H0hPp8eXHyUbOxO3t46L+Cot4
Y005FOhP8PFxZJrx1MzYEWdFAiNAroesBmn2rwnJmQtU8OLQ4mZNizmMKdXpt/2W
bmSmFvQUnroFRawK6Nk+r02pDNTw0oLaqkBX24qtozXsB9OC3zldv1C1+JyoAi1l
qRt7knTeq0QzSOwBXcn4Xo0Tpm1zVpKgjvp5kCF2hEY6CyRM/WCGz6bQjQllg791
xdCHM+XNBElxLQGV+McQQQTJgijk5yqKBxilCcv6dMDpkyA7uAKsN2QxgmR139vK
5h/zFvxgsGqUBTPoFQCpBoMIjHpK3VkOnTKeKE3OpJR0ntTWhB2w7I3wcJfxEHlc
+x7jpe+0R3q7tU/ZzIW97bYxhMFACfJpAbqp5M8k18dFRuKvSQ9G1ZWvrycJ0+ql
AolJGr2YfgJQ5YoloQw+Zr2c8X3P52qs+/qIJ7cCdZ6TPq4nhfqSbY/PTLkJdCkt
79PevId8CaWKhVMClN7H1ItQ/x1THmV8p0GzKZguyAwzEfDib0FM52SCuYRuhKGV
Bkq3X+KTYXvc0jwtOXKVuyXQJwETAmhvGi9QpGzVsZGJMAc0lRmCA7fSFXFeBpJl
yRy8ntXChk6TCbDgN54DdPE0LG3mn97TwzVHZKE4EA4dCESNjoydiiC9vW9lr67m
GgdXdZT4Sooe0VqGa+DSuUWEQxpu7zlA4NGCSySan9pcc/f2MsvEeuWXrHQnLW1J
/uQl98rvH/8oe/ubYvlhYA0inHmhcRo+7KS1Vi0RuocLH7EvW0Y7HG/dq6V/QiEH
3L+kZX+SZtxLEKZtlON2HoJziPHkVsptgEogZxpMSQZ6SroHE0s9Q36ksXKyEDj4
nDvZmor+UPXu+AcQNtQi+6EIyrik4h8+aMJI4q51s7OnswB7c9oJNJHpt0gx2hcR
/t96ysj7JhKCbRI6h+QTURDMcEIFF0dwG/sZu1Da2HstG+Nw4+C6apTZFvq1BTqQ
fDD+6Kvx23t9Jt0IiZoPVlQuGanW9BVcUWwtr3yrwwgS6JILFuYsaFzt3BLZVm/e
hkpRqRKCnmSn2zKrmIEY7VWl/ksRzAKp0gVpMvy6oxxEwljHxDdwDYYu6xQy8u5e
mEpPd2ATvTJL/nF3sJFGyJiisTtUyLu3Dhj7JxZlzvU1ckpHfueS/X42qktRPv7Q
Y4Tax8Km+7J8UckL1HaqeNFD0uvFoK5+Hm8LufnYECaLKiWhkv2uc7EuVPAecaI0
+hZNIkI+QWL83N8OingLPfrRn5dMKq9rm/6vAalo8PmWK0d0yAxHTAWzPBIBKbSy
sRZmt/+iQVdw4G6DQFGo+7arORaDMYlD3g1lvQBtCxIL+ZjRlvR31KScBnFKXOdR
6uCHsJ61HVGZLx2BgZUD3EeophcagCecXg3psuIkOQl//+3STjdmlnpq47alvUlh
p3igTNxRZ6Acw0JsudQMoHwj7gajOUx+tGnDuJRT9TjC6ubYUHUrDS/BsQ9ZJADA
rGfIKchlSqaI9rTymMo3A0Hbw0XK27/ecW0vj9ca3o9IBXZEhc0rOqszB4jp0jLU
kBiqJIcTmC9wB/Ttf0SCnCCZEmIkO+ph/KTvJBk2aWVsYGtqU0cMyKUsbOglEOXW
BFtiXt8l4RKpFG2YQAGLcDCq0cDajBHMyh55tqvgPOfyoETWSmI5HENI2AgVMDn8
Is7I9SPwIixb6Bwp7/upwZQFlOe99Lj4ICo0WyCdSQfmPl/+Af8PGtMFKDrHjT/m
uyaPVGRY/mWwQqRtgOlaiVsB2oACxPqCpAKgKi79NOuBiTLY7q773NEaa63RtNyV
jL48pA3HyCspwqQ9ViQvhUkoltBDmDEf/f4AIFi0BcBVsafBjN1xODcjrPYnteLk
WE/NzMYrSvVKcZnjhRTWHDtV/OJ/+1LREEWsc9MUNn3Rm8pc7STQqBzZB/kk2D1g
jUOYXuhRXvuVptdpUt0HGFHVL8HyiRGCGFWr30NFIdSqtpwoPaqOG4sP9IXiYwLL
4rrhGntmvjMZecbG71MSZ3AWidras6XdBDxRE6ImmzGgARdgFtOPqpkNlX+z7tne
sQMiRljDxSoWDS4MppaXZvn8kuQLo21IcJVEEh5Ko9ry8xh57hTfJZS8PNjiivlj
32KC3TwVH6bot5GbIOpJSpj3LwlTdw9d4tAEgW4OIm6mjEIvLcOnjuideeHijfib
LRQDlRI92NCAf6oIWl0JSDL/5DdvBgIFVXy68dFVVrIh4AAbtS7lqGXS02MtI+qQ
ldei+bqKpqiqJN6L8FZNPT4+3QTFAvEvIa3eBcIQSnQ7pjQflw+4/ftnCjTXgzod
AJ0+Y+LdEiE/NEuLkgZU/6yw/yB2crXpcVjKit0UI5Niow7mSvmcTQy5mViOx4eE
T1SOuhNIz1G4L15MkBv0qfmRGb36GL8M0S5OTs6T4Pi0bf/pZzaohlG68G5Ib/S/
6iPnEmKotWn9FcGK2MVU0r1LNNRPGP7dyLvXAeYd8KT0K/SrnMkZ25NNxqF/Cw6q
sqQ88OCYHIG94nrPO4SltHhLPscnFpwgG+9BmnmOOM4HrycTKPcWXdcUNpLgwus9
3Zj8novQEGulelUJhvoM6bAZwDfv4p7WZUQ3KwTowu46ZQbDohOChRRSkQEvmGGq
zftNPJyJbrVQU2Nyb2554AtfYcSwWmSCMq3AbMwKIlOoVu4rIlj9Sra7wS8bIuvj
m+gjsIh71J2yxXHEY+rxwsyTkBwXcwh44RNt2robycZW1j1QvG0lpKIqEB7fJz9l
JsMMswF1MSDK2dcgqvbidV3wy2It7k2tVDENGlAERoQkiotxph6RzjP6Ku5OQsQk
eHnTq4QMgzjHddzW9I53vZ/bS02D+N549mHwTnfXufh+Rh+xHoXKBezsOo1HgVxy
WiuOoY7TC60qc1elrPJCloBJCDZaJQy+2tmEnO284zUVXJQ4Uu64WOQ9EbhUDyg5
Ac9SetoeR+dTyH0QEvdXcVwNqpV5FhJxfnSemT/nWvERRden5qdFk1OH43hY0UGo
Ossu1yuva+ydBqcqmW6Ed8Zx4v+KSHYCZfoh36F6bFXcJEi1rcuO+jHY/xrhqktx
ibxcWgfQNbkEAO4PKkYIm2y/3YWkh7D9A/HqmtJLiZpDBi231RAADYttAgmQBeJg
c3eXwmkJLfQua1KYIoqzIIk3Pw5zCb08n8f2eujGfhteL2vEUO/zIPdnvG78P380
PTUF56tplLLkrKbVBhEhO7Bhs+Rf9xDofT/fVJehKUw9C4Pb4Ug/pu5h35oK+fZC
ZFHvoBoDb9qEKE4CXvdf/M22vwSZ+CqrsAIc6E2n8RppBWwy+swDBmyn2l8p4udX
gC9fpZojAZR4gZWe9kc41iiSjue7YB70nNLNQqlOxrEBYv2xq9Dz7xlKrlqSjzN6
SnJxpqzqHV1X/Ip3JAD7Tda2TvnXup7B9ChhorV6Wa410NlPpu6hasODmby1yr4f
J/p/K7+c/O7321y5gMLF38mybzPxX7d9XNMIl5fHhl82chOTUthzNxOJjh2frU7Q
iPy30WGYbSX2BAs8NGdCtvQ247I+9rB/jVJ0sN8smHXEjRAt9REkOiicvw1pAxec
Bqh7F1YHDpBYArz0UnBwY/MeWaid8gpg5TFXr6ig/VPJDzVnfaUH6i43+b3lqWWv
BaSB2myiL23UQrW7IT8Ve8zVX1PI89MoS+RWLWpWVkp2hOOX1Yr8nLMjN5wZAw7h
uhMYnQEPOaiJv465ngevM9joLkqbvvW8CRc2RKto3uB8un5odMZaOfKGDkiXJLk4
NN9r/vCRIjTLL+gJAIIab4G9cZD5AgGjJEL1ltPWdZWS9rlE/b1fXlSO96ljGHrm
5DBbJxsA1XG2EmDJgo3LccQwcKi3BdiPbTojcXh7sLSGsf1Fca3HEq0uRRbl339t
plRiVRaKMvGmyy0y7nkk3LHJEVZFXLKpkRmsBQX2vusuSz0K/PwhPB2k9jpg9ZI6
m9Vy8JajVUuux0QkW7cvh45C7LoL62lCRggkH4TuA806PCMG5RZQhXRKtfKb1uxX
24nLNi5NRDEzQpDzFKYD67QuRJaE1SRyh2fSbNa+bZTHqvMfeuMhbX5dwyVfp6UF
/FDrJtHQOz8WzZ8uL86JlhUPjnm9ILOCJ03k4QrCTUyHHHyo0oSJbn9Cgsb5Fajg
2Saxbc6L9TBjWMHymLTfs/iGBitq/l+V30mpLNSAShMK51eGc4CbcdhvsiJvxncp
VHatlClYpbIRheBMP2eMzVQp1siuwBOtRQPY93+KeFSFFG2dT3MAoVBoJ+tyoMFB
E+46OzWb8m2IWCq5LVStbNqC+x+EUI7B+m45sQTjeW7Iq2hJJmTdAWcUntaX6UZM
GKJBu630n27NVM2oZaMkJP0zxqhVoehrHns5kbCpHpEeExgmlxnI89kkbcNXBona
vJJqxRp/Fkjjly0LAzpPmGQWAYymn8MCPhT7dTU+9WTAfCWky9JKKljvc9De+ecc
H/XW8cPUOu/m22wNW/kFyoQ3IZxFgvvdspIR5TUKSdp93I34gUEk6QBXHYlWZ1Ls
byMBkPLHe3uP81GcdjpJUCDJZvIYNG12x+HTug5I6r4yqYB3UH9jN9hlwGIxAF/b
pTTFrHnRxL1I2rtpJG2SBLkfu5HF+JhZLn1WnMDqE1N5vLq7pV8DoqdNdV4L7LLt
m8b2ZB6cg173jCFI0zhjoFjbKDGI/2KraR4hHla1o8rj0y+x7ZjmZBXtsFHcqrFC
VE0olVHfYVLQHaDFDnr3ZoX2ZQq6qaJRP/4+JHJLi0odNfAL+xV4uUygVrmXBj6J
RZAkcwBHyp8eEK1rjhEez1C/lrSZOZWIcJTOONifhBIgv6K9BSfbQqwpYzMFGflU
ql8n6w7yXIesG/CQblt/wrz8chKGjN1BwM1zBiKIBzYA4OsX/oEVikgPM7zpnY/d
mcC+1RaDVi0MNNd7QhyzgceLn0ofN3bT+bxKjayS8LIvOg4hh1Xh2lPTmywwDlcE
9Uz9cLSPvZfY0tk2HRth3QkCq1qLCJSnIGzFJ9OGkCDfBiejJ7Gz/OvoHGJ4kZag
p03fl+mrRDvYTLcKppjOB40/rXt1r7kOf6fF2yEUfBpWmaEnaNsi3ali56yt3wKg
CTBEpUqm4V3eeSflq2J2mLW2LWODJ37Ro2WogWYyE0JWn5m82epfGQbQkN3d6tQG
ntVsMor6U93f7nd3IeGpGwaXHYU78XJ5fr5zerV4joCej4gt0+cZ9IxpY8Du1XlV
XaaHpNarIMdQAnp4Kv5IVzf+r6s63EUchldzhg+263ZXK3qfoxdkb6aQlwrQO0tH
54w2CoGLvIHh6TARSp0ranIGLLBBzNt8eoC8KNEKJjD14fFm/DzNBo1ZytiUPDUB
HLdFi1lwhhAyuLYYwvJWbafpWBbholn863L7BatK0PEWDVmk4XgbkYw4Sd1mBwXx
twYtsM7rIcdkYPXNfcGqb94Qyu6H3AklFpOgQh0UaCO4NnNWyrnrFeOdz/N5p1Q2
Sj93Czk96IPdcfjNSCeguJYLupeQS86IliBQIHbyFuQ5/5q4jZ7VxYU8H+MYb0Ah
dqv3ppX+2nMs5o4tMri9UxNM95lO6HIDSDUZDALPQ/ZyN3dZ72eOlPUAxM1R2ZJ4
fotYhOe81ErAu31AStJflywbVGSluWNMqy/nEKQfsllyjRiuQ0gN6QFhvM8C4Pq4
bIJIJVfBo/W8yAZ+SoLtdSnLVTutL4TUnSy7UWyNltSP7ZoNTnEexvuZIpeV3Zik
piHEAT+7S2dV1fyoos7hAX4YH/H67+1fR8emxTzq3dSkJ6j+phkWep+X2wyDzdPy
MUHum1ft/kGmerWZ5YtCxIX2VvnH9JHValHcw8vz1JR7QtDzMpuI+9bF/PDnNxXx
rOLRYz00n+ouVijZC/7XZarv5E/qu1K07+28kYVV8inRA2vyKnQUNtdnlbVIhh0B
P4De7bYQ3AeIRMlqnVn+J6eWIBwi5u6Rw2v5bI/lcczJyCR5nEOldKsUpf42L8on
56tWcA8y9FktRcZPVmdINfo21lF3/zWafuCkfxuhOu1Y0FjPH8xlP7u2KOvrXUdv
El2aGaHnbGBPNTx1VtroiM8GeL5bB4wHPDi6Tygv6JuFsSV67arktArNHNbgNSAm
7qsNYBJKfUTCbz6H/kOkhsTZV4JdTRwuBGQmIAZa0h0IEffAJ1KP+iHMsRq6tILB
0hD/BqxoTr1VsFgMBN+/+RuHdpSvH3yH4Nv7ZbrGPBgS3fwQ7ustf9lzsil1EaVX
XkMlAgdvHAc2f9ZyllzrrWhPnTO2avWtvIwl2WTFXW0jCFTOhv2tXCyDfbn+QrLf
eCHZE1ajPyNLj/gkgR2XUfVoygP52Hya27vO+/ASZ/196N9xpK8uzdme0eAu/x8A
p0CVGvK4J8DiYjEncxPnSBeb00kQb6NIu2d1DVwmbYSnj5Ki3OO2DLBRk2byxQLi
PKa1/IMEQEcF3zx83PF4UeMto6MHpWXfimdjQZzBIcMM7jdGqZZc4VyfqEzvB6lb
zZAxXEz3uCQ3ySkdwVSeAQDrTov+GE2Nwj9fh9ZlLXv9RyVDDoCrWwTv8IMd9XeO
PMPUHf5O6FO7t4k99uTu/9N0l52ZXKEMOkp2H4XjIk7LO9ZW4pxsJLFqXU/R+DFy
zta7x0VMku0CVktCGukfDR+eVLi6g471T/k4TChvjJ6zmjhvcCdgWm3EaDsCZilZ
76qKLBjXbo0LnjP5nQD7oNo63D6mNdaoUdA3byougQ4rSpAVqQgAWwy5D/TQ2ibo
a+wYqaQHziGG0sot2DLNx+eYZK+tMqDLyeghRCtNwByjX43EO0aGT5PdTTvXl+hl
2W2KZ16QikkCFtmNzpDeNDrVyjQYnK424G8Oq8Eo6kcGQbSYXKsJGNevV/83tD4v
OLgydYVfZyPaA/4wsZDfpHnE9Cyshv46Oire5iVfV4HOajXEW3tvSIoRvDJRJ6EX
VEId4dQlht4HYDeFGgl18JpNySA3N/R4RN79bw+1CM043kpc62HaazejDNaA2jKB
K3FDatZBglHWn+TuVnm2Z5dHRf1NWR6d37T9xJbzQQIss89DPcBJp25EfVKJpxqL
9VWrE8x1ez1ukChFArOCqKfxFt6kdsBfOk3JHGVu+7gh3CV3zwRP7b1OdetPWT1M
FtRIciJU3nDoaLGe9rOdxAS277vM1flVYS1oTDBlv7j+cJofdxmInnPvHdTELdUV
ov8g7BuVkgizfIleD5289nHGeWpTk8oo6GKRStFX7SH6fih8n5b9qFw5GOHZuYzw
y8TZ0mYAMsAXWkdMb8QTNQVUbtX73HTFnHsb+2DIPjMpGO4hRUm/jnNBYHGpJGoq
dRI8XjF7Dto9VHUEg5Hb0Slr3+fFTG2TgAJ51M/JwANXWOxEQHQyTn8Sde6mL4Nc
n51wswPpbCq5lWbne4GfXU/Wpgo3JWg3QdVPcPZYgXMWdcm3Po7Ic6tBmsekMDvq
SUv72cgx0vFrJnSfDBWnRyt+2nha+jIcXNBhGMBWOmpLVIhnLIjctfoGkbK9jNY8
g5daEpZlAZ4cEY0HecybNUFzXdVdjd9pvSb+zyUt5gXl7LSnBWWYlbjRMfz4LbWC
3lhsI9+8uniN152cuqFmeDTaE1VyhDkw8+eqCi2FSOsKd9RooPzMfL280UEG3XFT
YCBjBJoJXuCtLr18InHM7CvEsyAZikcTNGKpK25NJG5VzYgzm8CLuutufLK1Nmh3
1+YUPP8oRbEQYSEKhlG4RhDjOBPQytLBPHIGSyNjBz11KSXiMoo59hadv9dXETgF
H4CCubSth62HKcuqaFEyBvOmJtMNPdIZawfKtTUh9r+Gku2bKR1XZJgtLsZbCb8r
Gill3DCmHGM2ZALPLuY4YUufphhlP0J3SRCqV6w3n78mlW2N7Yr9+zrsufFQOG6E
10hekrQ/1wk+PY0B+JVffS7HK1sM5TOt+HTvYs22ygrWT8UdFcd8PHs7SRyjr2is
sAICnLaJRMvt0Cevw4C4CGKLOkofnygC/tqyDCtccb1qCRCx9fK0Wtby5YqZPfil
mVVRaiFCfBUvKKMKfg5B35m3Lg03eyiarcTK8Kmm+pJRji1g3BdORb/3SkZtg/8u
1J6WnUbUFEFyp3k7rxYNwt9lVS5VYmwqBcJ6M3t3AwYu0QZNB9vzcCXOfCUEB/cB
+BEUgZoTFMn622aHp95K5fWcMUpphVjm8U3eeuyh9UF47udbmUbYUDzjfHxjgg8H
PdAl3beyzKxG65vW6+JOHqtTAEBxGdWBQTs9kDzamUKxaed6IqMLUhRr2rpFCEp5
iW1Tw3KX6sL1aVpn2o1vbo0LJ9UB0+S3/vgEIMjKs90uxvvkNeZNZ06Phyk1Rbzl
UjZ50z4Xt40uCPMBvqt46OMQwZlqk3xeu64Qd3RW1f9CQFBJrvOcsgEPb8Cknw0I
W7pzqmarGK4S5f+tElGHFKFtfzCt+zuLPIERt0ZDFN4njcVEB3ppbDju3wcjfKp+
tDFvMa7q6F5xG/gLx90QB5QoHyX8P+eI88DIYb1HTIeHxk6aug6wZ20+D4dDEl4a
j+va3wCTD0lqNWjEhHLE2NPHyc7MbJjaNLC2wwbku6WaN6j8Uo6g804ehI4/Ah6j
R1fRlIzv0ATFk5XhHyu0RjweGUOd94xJ4EtVX/8msqDJoW1mdXEhTWQ8+hwHPQNa
41b+h+LMgAov3Nsq4NHB0yLANLVaEspaCD+2wt253ZZ+XleEkQc4kv///vQbq4ND
6vQ8Q07jQICfMlA8LeSkuPK/mV1zyNfQsrCydj+brU5w5AmK2RHcthXanJle2EEd
QO6bBnJoiDLdSbwoKRd2zDyumsAeJFaBl5DTAV9kDlA1q2coedW6FBxmYhLGcxle
j9vd6AFxcQ/fpZIf0S2Ho4jgta1LAynCABLN1PYlUYEaaGumdw6w/kypVJLWSUfR
AjOkFm3IcLzl5/qX5pGVE4MAjmukGSE6S1obw4a7VYRBMFHF+GoTSML0OT6ARdsm
VRAjNFWX1Iu5Ez7JfYSiJGUNkk285c21SJL2eNTPvy2N9gceT+N0fAfk44ynSDa1
LWZlADyu6EVsNAcmIFouB44CMcScg0+wFh5wD2fe3rXwVHYQtNNYtvTXJjNTHFEU
9wOCcatr+8lWMzrCFscCW4g1YCgRglGZrqu0kZzc4ipnAyj1nu/eUXDLmhM6zDaF
XetpmvRCXrWy1Ov+GUdn2bueE2AbwWKF96fD/EP8GhNQtRW5NlaigdxesuEawQ/W
2bCnfSW1TsTn5Id73yHrUBxhdeYHGWKqNbvAM6loqLXKkp17K3Xet11djS9zg0YR
SK5BEXIYSFOSyts42RU6SsSKjRPGrwdtBuXxFSFEK+kvyS7Y3LdKXf+lLgLmef8L
01RsNnweqCn/t6E+Nj9Qhn4H+emfq79g+dsZNHiBxnJoARjb4hxjlaXPrnxtCL95
rSJXptYxdA70CYdqpNcWFEda8yQIEgvu104d3rLl5rDN9iNyNrIv2u0WWMd7LE0N
GVRvPs7PJXvg5u5O1+xazod1PAHteNDF16Gyx+80BPlp5TRAePgFWzdiKlX+eb1t
QCZUB5ICNDlnW9diP5THyMy35m2qFIICOxAugWArQgVaE4C7uO+GjXOmRAFfP/oP
F8b1LRelGiPIpbjXNrYYmBUkXcl84PjlsAyt/cM814VccTUPKCb/CHNS+t8Ctxok
vfGyGC7hs3LwC7Vqk0E+WjNj/ecDsGWv8T/NAUvXxyMP8cY04DyFbvNq7lb7OCeT
0je9EcKcXV90AjcrGP84PyLxgX9Roru0pGr0SYoPg3s9ylPk46+1l+39mnVW0bh8
GRpEWebDsWZhxAFM39ZfBTB8G9BlPV4kfqbehgVv8hRyvFGeenTLq63Fk44sRgLS
/V/UIcx19Z9zIm/cK2b24AKKYwwddTtjgsxD3vlRtr968yeBD0U9+QL5mE+VZrEY
T5+dtX9LewM4Df2LzStXYBReYMAW0qNg1qj42RWWmf4BSyKDQWO95vp67djkW0dj
VLJEmtdPOS0FAGlEFT4DzqXE03itOCKm0MQUvz5OCGDjSpHZlX0vqAxtam5j/ChN
pGIOv3DY7cZmyXsg36bCms8RwO5YuzadXG7LqkmIgMz9o17uqVT9jGsKNoCE35WA
MUPFUPE4vCIDjY8FpnK3MrWk1N3GVkEJqsRro8O8A5V0+yRzGbhpE63Adv6T8Hzw
JgIhH48W4yGQE7fRzHlV9NPYlikBVwUTLWwM6yqo+bCNqIHyCDfFaxDaz1byPPX5
6B6cgbLBpjKfhqKzuM/fmsMvraddcuehdFip0iSB61hsLxHSnr8ndtA4PrRNuFLj
k54bqYKrZczEuHs+yHnrk1ePUZI9IpGSenZ6/xDlxgwOuCFY3KrCBnk98dv3cv9h
ad1vD5hB8C48b39Is3IxcC7VxI0DThtr8f0n4jdOXs1UwrCH+MjRlEN1ST2c3sBb
EosMGloMQ0xtyXVnwJZyPTnCTv1mj73x9nRSejw6LF+0OedYcePUuRwelV06+/P7
WCdFfsVN6EXAA0AmXoVnsRXr0liPYjwsQyz2o0l5iowDHdqAmJiWD6LNlYuuWLIo
Y15sXUYusSGBALneariavUGydCf/3xVxWF6R0dxLTA5q6VgnxFm6zQ3BViu66g6F
1KHPOsdV5NjJOC0wjsyJn/hnMLNapckX6DSEagpBlrsmtmqjTKP1hbuXwzY1ee0i
PT1MQ2sgnFqTsYR99RN5Gj8LXokg5LRHOxoRYu8gCrxJEyrdF8LaawYL8pFHD9Lj
Cz2hBLrPFEw7zp9KViOIY27liTuZohIZrrY7YWWepR7+oLn1IfmVjGB/wjXfn7gI
O0Y8muy9bhevDPhQh8tLTMtQIBrQiLVC2XlEnR1TWvH1f5V5OJRv9sz2b0bTV607
AMjfjY3xXZBsmv1r3yB4LndnH3C/Nbdg3vEk6XfuOU7btKFJRtv0hDEFnJYbLuMm
KHW1sFpStkoXhXkp7wSK2zGAlskTlYYm1KXOA22nXtavvpTFU+mAhW2vcEQ367b+
6czNWyAUPYUx2iomeuLc/DKeYZNpKfdKEKEGBQwnwHuoJyA0CAIZJ5NhJ14K8JbF
3Y8+BRvhOvmOlHCMD0TMttg/Qx6YLd8sHZuNodXZLgWf7DflA2QlyXfGW4lnLeLy
DuUG5DZtM5VscIBfqD4BblUJ+OuopZ2+VCaax3XKZewIrfRffV4Os0DM/rLD+y9e
WWEv1eEbCKyr+rDOYkk/D/61oAo/HkVQI9eeoWOtGuYBdp42yNjN1tsaE8//qGMH
A9vOFUmQkvAAJq5qYLnH+V888MMh0sY7OnBTtLo8AxTur9ibcqLnCIT0SnIXvwcz
0oPRNg62DPk9EJ557zduJtr4lHhNEYmqIPQw/xq3re1b6kNeJpgjty1CLBK1cIff
71dgGB8DaZEWqgZDx/s/yGglhjURsQvxTppKZ9f+JyoN5cjqn1XH9mjXmxTQ2JW4
6SnWEqVhtm0IJSG6jKlR5mukqvfi/z4dPMZkfSzhjwBZpiUE0WPiMTBhW/PYNhcc
DSh+/PbuZhLtnjT0PZNlyBg970Ux0u2AxoX1+OzwiaAJh2ln38ZbQPSxdKUQ6MPT
vilWV6iimqp6p/d1YMQ8I+iPak6srv4futlm5Zj/4O1qbbaSYUFGNiH9hHG9mH3C
2h6ezvDw7Reu2knh5HTkYtvosyaFzmCWoj/DBKgR7UubwSr7QWt17UId38hp1Wp0
fN61I8owhtBEt3Go+xCATm/KRbwy/L5FURJvjP/3s/AJRSamo9VTzX5JapeKG6XT
PtVpBcg+5TDy1MmwG53j7bRAs982UY+SEKj+UjeliJmX4uYDlNmrIRnFuAtkpjI8
RqOTfAHs4JHhyM1bsC8npcI0dK5FMfMyQCrwUqjny7fMA90Rn+anzLLYilo7/6aZ
avLFXplhYXNkFDCwzS/v+piGiopWyzdpIAEGBIKZl7UMUreS1cxj6A86NdUNYYbD
yRJzb9Ko2Y+V4GtFfFq2Pt67qY/kG8H1Gg79uMKUAD67qHT3XzpgRB4fQSTFU5he
3SwyFCVxIWmuzP/thLHo/DXHGDIe6UugMmTQMuzFO8DYMaHvq83OaQw5hH371hlf
fSaJj1cwZ3Cm9DeJmTOa3Z0ocK84p+QdzO22ztRLOcN1bkpTXoDffTgaHV3rWG/G
G8GU2NtrKhfEVm/4XYVlpCuxJMEYLhv9i187WThFH0gsVCTGP6nRQ8O6smB2aVG4
qCUw85t+xcyKkE1HPXYAY4pd7V+fv8EOug+DfxgsuKIo/mS2OpgUtn9Zus4n71nZ
FDnj7e3btVEzUpdV0tA3+fiub9ZiLfdrW7qyPcs1aTvSPYqu6m8c1j5mQwE2CI/G
bqFeafqnciiWOqmyGN/5cswPwQGKgzHNRvY4fe+rR+rx1APNZnXGyrRXtGNTQBWx
x0JfTCJ5RNaezgvuLlJEd2SQDyP2+GGpGp8xViD9ziDwa2rqDZmThtixv0CjQrds
UFeUS2NQ1AJYV5eWjd+ioBaM4oE3OxwLVzSJs3RAr3biLbVkzEyeW8xHxK93vbfT
v8dnCWLn5DSQZ0F6qk21uWmXXWC5WagL/5IS3jYktWXO8G39sRiIo0nYd+UXfDip
dyy90RUnuD6UA+ZXEzPXk49U+AzqBRT47mxZHwf41SyJ6LM/WcRZfH1caqwlAmJY
KB6EeApx9P5GjF9sYYVIoDxZNAnRZczCsGHNriUOGh00WgDS7DMGGHHYyTlxeCNn
2lFmUsazkbbx3r26FZPzaa4zPgmBgG2F8rCKzY1mSMtDHVcTaUWDyjO3dqwZ6dma
fbOMfuV1geRWcs54/qyhR2RBnXXmNyjMkW8KIyGiak085XNo3LyIYJ4z5H/0guYg
TZRIKTQZPT5mOQk5mHLm0tJFS1BVDOpf2CISrgkWnzq+KXFGz1utQ6pEW9sggle7
IHvz5vWYrbGH1BrxCNqhio/qrDu6BagyYeFek5G0XPcOvxh8opeqrwEis48BOFxL
HMXVxHspySVABJ/11xo1o0AG6pZpI8RJCfG+o015nZ4+xGiyVmEg2feT98/yNMkr
nkafFMS3udSQad/eMaKlWljQ6wh3+eULvwq99PVtSIa/8qNNH/cEAbMHWVxEW1OZ
sDakz2GhmpiuMSkD+yNzQQLlSHWNM1TH3maqKMagTGgwA7R3o8pYhTspMPmFL8cU
jq47rA+HiBp8FyCyAluR7ShW2QEb7igseZpCqJDRdCzFEAdzEE+F1kyZ0BFqxmG5
JY6WmrRtDvqgRmDAXv1bOuV6/ETrrq/GL1oWFGhQZQDJKIK6SrMEpl5Vxb6nZ4FX
3TQIQtEdi+w5M/LaEJA78WMpKY/h2muEgno/TAewxnh5BaBCtihJyclzS2hG+vVV
dETX81+rGgzcrexI7/RY6mrene+WbSewln83f4bXceGT3I2uDH+4WyzJnhwFD4b4
OQjJ6g4pRM7uzsI0nSSeQFHcnHS8M5joNKK0KXzP1g+o2d4U6FSl/nGYz6/V0I+A
D6+g7LhmGPs3ltYOmCT7fUO2TMelZaZCZao53zEttMgfH3j5MvZbaYaMaWjKq0jz
7xUm/WYy4FGd4D9ceBdV/8+ibZEEgiXjO1+rtz5qJXv5Ths6L7CehAyD6j92qHGC
cf4fPGj9lHRw6DIY3SK+x1NrrGGMz/jdnEsCD6g3JiMY0o8dJV6S8RurICws1mKj
Nke6Fx9mOgUc13a2lAM1Ji3tLU4CHfEXjC41LJ8tswSq0Z/TnhHb/epRhZl9Upps
OAzCqFU+M7s3ByDJrEkBsOli2zoDjyHZhR15lvuK+8zxXpDIeH8QBd7FM6LvEm28
BQp1y/4j4s9flwHwsBUwcUPq9SGI1lRCmmQB/B0h4vxLH8V6uOFydLqANHNGc/gV
0/3sTAvR46rjWBDiL0Am8uaKG7+s4n6YiX474nHhriEtJ6jq1WnmHmpvixMEeBl+
xMXa+jRFvWXJ5pRaIbRH4dvO0ik0kSC89p3+YyQ/x/cs0xbIOKfsniVucKhWQug+
tsW+jDt6rVK40kFghhag9meibYIgVX8Q5mjqacOewwwzFSafdat+hxbOAl6sNV4X
1AAT/iGrGO8wlB34s4+MYGsz29AA2hw58dafYQPTHrlOQA+80DNxdAyp/5ZUIkj5
REC2rCaMaiuuHdnSiy5yEWQxRjkT0dd6IBRUAk3oTLEmoKTEvW9u4qzpPdaSwuW3
L/Hxxwbybc3z5z8f8F9wpvAF72r9uLtTgMFCaQa4yAAE9O2f5IfVvNaJChTIFbL0
Wc+D51GRzOMRA26t+MLGFm0V3SmpNAFkLWhTpwOCrqw4pBidVp7DOrNgC6R4hoiU
jPOg2XeNu47ys3OEFDnYjFmGmT+rs4+FrqlEooyoUd0waMnvFWQhld20FqWB7SBV
0KwH8qbYg/xVqbpJelJYvjBC9a8gm/LVnkhjm0noQdu1iayAtM17iNgIgJgkJicE
wNqm/P40blFYXtfvs3+8t2iOA+gbfxSATH07fy1yZspY44C8JkHfr5Tses1nGToI
LDX84hS6SSjZ8G55eyft1O52lzlWqsmL27H9yh4bgtYjZnC8YxbamLiqTU5b292U
IDmUHCJ6G0FfNwzoFagoX0ZFE4Y2lTIzbKjvV0hyq0kAWpo0IhocR6zSTuErUOx0
bzqshXBdWqfeYtUqEpZ6J1bzRKzjQ3HVteM1sHWRZtoQYHrPN1MKdbRA9VKfPgKe
3DPaNtjIcpPgTLpwDWyuOaHmjHAehgYiivg3+zrC16LFxcqK5ZT8lvOU3cGS14X2
DLMhbMFNRBn7UAdkatM+ff9qUpQ+fFSck+1kObZElVdw8F8fAPeh+nt/cB0kmIIX
DoiMPBsUH2ighiYy7wsI7XHPSNmZMFPdzIcZm7aSsCsuiz1n7LEx6nEFyM+ZA8NW
lRSMoaTj0BKFlquiW2UiM+t7zvqEr9VmCAv8kZMuhCSoYc2v3v2Jm8C8jUKKD0kt
EBU/i3UfLow6+DpS9MHwEWkMF6NJPAl3Uk4+LGrxk3rQj6z/OwRN8nDuUnDqRSwW
HJsKKXNbfFjVJ9qwkPGz4h2YBxr+bpJAdS5W0+00B/HMIhYf5Ir0pLfsjO3vyKXO
pPgBSvLr2toBJfxBMVo0OLOm9hIYjOfvvnA3+utWadULpMX9UI/DAlFjuRVQJ8HI
/mA+UdabPTcRCfRYn0Igkhc/NogUKiHdocooZc6vrbCgQoPQkvATGVbwxlnrMT1v
lISazETELG5Y4lyLRDoxQKqyDpxEK9ALlX8b3pwmP0NeKmBfRu1uibRv4lSjay5k
JusSEVsssr/j1qJYhlVRjl7xyxZ23h8htd8yPUmTvyx9Ds7xGulDjHee00kvnZhw
t0Ar5APbp9adxBxHdKA+PFgctVoUH3jpK46opnMCxth4vQTbddJdxAWM7maolPr+
fvspb2BcQ9CnBSCDP2ZpTZf9f9k7+EjePnsguqETxRF7Mb5mKEQr64+SbcFH5Jto
IY8hVWQ9SbhLHv+cfm7SxlOH/X6pnQ1Tm3dRb5cHHEWnY1ZMrqFTmhrH3Brn/j50
NeFqVGsVMFSfZra30VxhBPkrLu19E+WFQ4x37RQyHZvZTgG06SCcm4d0tOOG1OVw
1CNabASMlGhDWXA8SHbbNWbQ/QRbL6OJRzvKYlgoNaoXxrg6GKR9u3uPY7NXQz0M
Ix2gZWxmtTXmoj38PUbDynQ4jj0ZYxw8XhsBS89Ywa4ZFLzh/gyiRAVOKmGwChGu
7/mjjvQ6qRDh6dLLaHVlQdxjAnapTYKyhVoL29DykIfMtx1QrxLVpiSEsMXlODcK
DoxivdzprDdl3YbXuXYlLa5HqjeKP4cyAxnWyFVGYGRhj/gYiX0CN+jCRgsdu7Im
1Ujafp3Y3NGgikbeNh9Z8WdjzoII2gIeZqL2wz/huNAl0+0iIy5f9DREKtG8sc+0
wCXCWUWk8/1wu5wGUv0FyZUvJESyaQD8l7/0bFIkrCD3KK2ol9kk0rBmwt81Sfva
3QN5hi+1Ct6o6ari2E47eKQoRLSOyFV/Nd5s4zaReU9stRLBUobfMK/V/61l862J
uZFHKEo6rd/wgw3vZKqKWVhXUlgzUm5DcqTHcmkhxfVWGOxHEh1kpfFzjyKAJ1Iu
SxxJmM8FbFHDUnfDqCQ6UUICIYu8k7nkITDWF/ODIpuSDqkMsYFNx3adDwVQFKLX
1SCtXfeEpH+UnTQbBD9/QO8Ey7ILDGyhvUZSe6lvCv5pV47HPhgO8Kws8c8a8gOn
gFGzTCxtL9mhCWFhv0FtRbdD8d+vpo+JktmM/BcsjsLvLtgqDNOuq3Wtsi2lr7CP
Dfp0Mdu54h6Q5pG7ayqqDP5wR/2kyipdgg01felN7g+Kql5U9lnHcBBpB6DFMv26
jgC3NG4GV2QHnkuSHgYJcDE27lRedh3Vck/bYsUd1Wv+YXX9ltT1OTxm1nCchDxv
tuLChR80nfm/1dacAESEExx3ZayNqX78sGZxWglO1OeZqeosZH0R+Z72kCz598ye
S1ZwVgEooBAT5zA1iq6wIiHtPndNhU9gE9bUPAQkgCPmNkl0NvlkEoPZBiw+qcQg
KkBGVjbyuwnRjAlo82BNJlvSHvFzKnyYTtxcVKgCVoxAvuGTJpgYk/mmOXc632fI
M209vagF0ee/oTBEo5P3IwgpNgr/xXDcYmuIAkiz7dYNu4NS4bkiKBUM7v/kf4dK
iYWPHNXGcEz6U/3JMLE90WCyTmdQf2o1YRI8qFwWrcXPpyL9Xr3nslSTaHiK/kc+
//RH8YbbbedjSY6VVlDjRSY95lTV3PlS2lGfTU24xvtytG9xkQOWHhZxB4lJSH0e
nUy8V34PIGS/Od23lBHiqX9UIucQ98teg1QVfVOsRG/0G7X+bfroExCQ6uGdeVKu
ggsX4EcFTLfJXgnkE0xq+P876AVH1y7tOhuitQ4wQPKaJxjNCYmIJmDd95zxhNas
UsJ5l2z5LUrxLb/TL+Ij+6jBvd+zsK/O864gAnlrSlaltR+E5S2apVAdh7lNjuPa
i33W6cKomdN2pkdC74ouZ6n9QWxkcakUastWqiaMTyxPTDBVl+ZZ1Cn5cgijtGGP
fDmv4rqfEwv53TCcUnaHQV3l7nFpLycJo4KildyyIxu6YzOV2VAEqfL17Cro2jSP
D8mZG5cn2u4wPp6z6CkoJPsYd3HKcPEbXGQjZavRg+d51bFZF6zVqDRh/fXlw17x
mPYrZheBRAqBmoYri797B2rk5CC0DD77vl6nVUDsNcsmxAOQQinVFGFfbbGBFIRV
qdK/jJc40jYhuU79lK+x1TY4W0Cr4btNYECDXwb7kI8dCTsGJlD2zDcWXiTZqr0i
fpahl/s3AolsBu+KTi/NeJeuIPMqK7T5FfxfcBZzQFZttLSkyRFHJwkzG9gXrr6/
UHjSbt3Q+dF2IdwHAXtXVAjKlPy9/OiGnnHaLiDsMhw6Ltsz7ARvwitBz3i8p1a7
jgrRhi1e0ogBaFkMazocr6AbKKTvM9PmBC/pccax61eHXIFD/N2PfLSXOKEUjg2E
BWTN17aLzqOaRL+5iwLJuXpuwDoBL9aDUltXUZPZR2bNPwuomrAbbVqDIilYm8g4
PX5ZInhl4tF4byJMWstpxIxjpf3OY5YQEKWVEgGZpdRLgSQPIS/MNIGH5QCx46AB
KoE5m8x/VsdMIpP5sWQ6o60duMk2gHehjq9qH3occlxOz76mXJoLtuLqz113T3bJ
+qal8T2br4Q8y0TxvEXZEr5WJTynIGB7JSGj7sD9XmnZ0ey6mimOXfVzo93zi+ec
GDYCCYGrZQkTntZyiSaW4pMG4l/cbpQN/nzDHJgE3MuYABcP0K9Nj/lXUOK9Lp9q
dLkCaxsBZ2AK4LtOp+1X9BzNic6imwh+1sOHeUUSjmh/2QD0oj8ik2Is4MLGqNKe
9U4ng3Sxkii52TKT++UaxoAhLHaznQu6lTYH8NThCi7qqTzcBLJR6cK+44vPH/AN
VUlgERpyXK+ChYAFpL3gknwuJsoIwdP0TZGFScPcD/vioc0EFTpUGJcctgMKTlzf
Z/NYBIDG+YACXYmMnfN6YwN4ccv6UKGo9jpf7xTsSwAssK0RFa3eJiu9L7ClaFGF
O7wqbcDpJqq/JZ1hMzxDwbJwfp5PzfgQBQfPOcv4AiCSlOaX6evB3vwAtobsJk9H
D/fvapguxENUvhstTGazuTOyCkuEUOedUn4zziUuMXP2s1xMkNosXIjyVt9swQxu
8gQeF4+/YegKs+/005pssEsR1YNLZ3nWeoVW9vqWqrb32T5ABHfPxryvwp8RMkKZ
v4fWplit6tF1PvTQcnr4ZMHX/eejklcVhSZ7tPKhB3zQ5vQXDpMiK6MRWd6lLnjL
CI8Balhyd1NQ7s/b7arjzeBm6yaSvblSL620xJRLlK0rzrTz/TsvPbPQ3XoVfKnQ
A78iDZuq5CXTjHvnZFTWnGWDrGA5KKPVXnQ7YqH4L8obaYt1iD2c4ptupA+4aLCd
dfpBkyFrFwNth2PEbBIAShbl4U4LClUenM3DyqYTHenCVZDIqtfhusUJe5gaR/O8
1Jt/gB7Mm1a3a+6oJVmDyqcibU8UyaERMJnxVvnEv4YIEhRNahzFYerO30XlIchm
7IUiTERYTtPH3wIyQqrDQFpXyR7sJmu4XwR4OkO+9/ThaVcqExDdKVGM9u62VPfO
lE4yEvxvofLCkGlr6FUSc0JTWD7itQvBvQMdKy81OoFjie+ATTTrUCDWgtMM9AhC
EZFsj3wwOe6GkDbAiNApASg9X3OyrXLojJZSRPCZwJZH1skMrJMQitNDgJdVJ9Vr
zx7Q9s3TTkTn00w6Zqi1ceyP7HuZx5or9hrXUY5X/DtMZe8Ev9ic1bXQ6D9DLZuX
cwIOSeqHia+ueHslhYVPfxFtTnd3XnpBTXlgLKGdt2T9bU3jjRIJAv9zZkpQ1TcG
Zcg37Zguk7RaqnTiz//2Srv4Y9UTtou43WPPQ73r+bFaYa/avlAMEJazbUruFUuK
PJec0gOoqr0RGiINRI1sdUKPrP81lP2aclSeX0RzQprPuDbUNEWcF312eHf+c8r2
BW2auNVCzk1UADPGtvbPnS+RZhF03qlQKe9zH18dszZ2W4WD5l0YWpjIQ0VsfxgK
W3CR1VBw1ldDYiB4un2LB5bNt5qN/uHDpsoONiaJ6abGL73kKjQT1qldjEA8jBx7
oa4QKg/oFZ/RRok6YI/o5JkvoCu/oWmCoYK5+CHOK40GcUVS8DNIFWnOMrllS8bZ
c7sSdrVIkJTjCyJ4AUQv3RwW2gg4H2vSogOHqfKf5gYt+PkB12XD2HCUFlnMW3Vk
e2h698mtdxnFXFR8jp0R+BbqMe/r43+gsZbCQhoKu3G2K8EL4tk4lSPwPl1lGGao
y+fEjOPWkNarcf8Qy7ZATwciBPigJmVvFPMMTxxUCg3xbYHLE2iH8hhLOBjhP8wa
VH9fuUqTnEF8uFi+nOUzHJW6FKKBhsgpZ++tp9CJw9+ERabVCPCfZSsYH01R4TPy
YB4TxVDEog85LzbWCjbvrAUuXwLaTGxSfFv60DUflDZcvJ/3JZRY9qu0SY8RpjBP
3aysP+bknBGZmeZmhag13npSoCc6xBvtzd2aYKVCbwam+8QvkyHZMtQAB4rMxbno
5LzmFF/HLiKFkoQDrv7+YoRWpJFItce4nT8Q4GN1eaJoGVcMKG2vVpn4wKMRXQx9
9+/98WqgYBOdqy0+A3Yb6RFGsjM9SysBDdbSs6cAUbwSVCkdScQYl9jCO28sBMMY
apDQfQuXKbZ+Bx7dt0GW7Xw0ti3N4wnWT2Hf3Csj9IEOBwLSAh2NbwgyzCrfyIm6
XxGCPyGmcvJUNsSu27kIjpylOVe5Z34AS5uFTPo0WWFWLYNQz7SbVfAiu4WVmX1b
BSC0IcHs8f7l4qEqGL4BiMuR5/bN66ZAXrfjwWhsw4b1bRbrjsES3WkpBxnyTVFn
EpaQDFdM6LK2qZkmgcgghwkN9CYRXpJYKkZpeDBS33R2GqFn2bmTpAEnKdPSE42V
O4bkvrtc1kqTmWECu8FZ/ttaYo+w9O63hZ9mwMYZMPsqiN26ZGkHBwoHaCrc8+Jz
xRD0hJ9zgggu3ZuVlRh+kCTKz6Bv6eGSorVkTehqs2YepzjwtQDg6Nt2svsaS1j3
RV8xoMXSrs30lYWE0TSL/Touarp4ebz9+NPUEpkHfIQg17WSMj9aXPyEXPSNj4q0
KqVOLYZhOsgIHsUSDcfRjiIJC1rsRKF88U+3Cw+1itaO3UmPWszU+SkJ9FelN3Qt
ZxZjRY8vufFJbwz86O6PbIaZCUE8781c6AKVgfl0rzvSV/XRv7FFR+CJ5BqFfk77
VBvqMj7MQeljjn15VLIdLXtSU9GLTIuYrqSnJiWcyQDhOM6Mua5p8HmQ0yaRhCmu
h8rBAWgyDIT1WghIxTsSK3tjpaRx6tUriKZLnZJ6BS2ZIxKs+o+b8x+7LWUeFtTW
OcXdAkDGkF9IhTSzQAPaQLGRrxYZPm1E49PfcdxNAwh2lk9VcA70KU+8yzFsvdme
I8+eCW2WP7m7gyvzbUyg/UTaHYbX4PK/EOz2EkM2DHzukIbJFSqjXVzJVRNRX8xN
wNM8SNlfnrSgxuhXGeUkfW0EZA0/z0gXmr+eMEVn08fzOnq2YxgfXiaQw4mf11/q
jZdzbvcTosCKwqIGXA0rgQu1+YflzplKhssuYQUAqZOWvXPl20Y7IrbKbr2vbgxB
eAV+2gk1rrpi+Mo7qRIVkC5kwbl27+eWzhPnqOdmXVoLfVnFvfD8yC+/3RMK423u
mc4iCM7fJ9+BPssBYl3Xl8kQqwgSJ63oSbOVi8kt77RUBQOutGNsUqxYl7UAX7hU
c2quqTdBblnsFH3HscKJaTRoeQ+v9WFndt1J55nqb/tRE1zy8U+4l6PkO8b+CNBc
2scKZz87iY+ZxksVFr0wTrBEPjCJQxUP1xxwD84Jz6ls/R/IXurSOuvgKOCVyA3z
uWeaovZ5QX/uFyHzowpJZTzlEbAy9ro4U9a5mb958sNCwLoG6d7ejX7LOfKATkim
JFTBOpMkeN0hf13I8F3XQ3/lGUTMwSOeZfju+d2U2z76O5knyyFFzWuBnaATheHS
vHmRe/pMMwh9n3pj+dPGuYfVbvnFnFeh4PVqdXtYEj5O+k776ihJNnQCursV7Xga
wQlNSwCzmj780XysCsQW2k1ch3kFsgvoUGL5rg6OHMFv8puC/TnSRg/u2ATMV3MI
C+0UXXi6KVPiKNTLjTm6wORx49a1cmjRzmtI7teRijAFms+sH8CuX9nt//LgbEsn
BhO3Hfjr2pABRka1dCAtA7GclUdBnI/4lfKqxjgRu6dSLSS0EEjLJNRMNrN2IptS
PyuKULCrVGnWeY4K0VFDJd+UFQck/hHnllv69drFY3sfh473jfI0jwLIn/FKZFo8
umlmWX/fcraLro/fvNmfyJButTZuZvcqVWgXZYXS9y2XdQuhXpgH1QcglDn6mwC/
/uFNx7mxpLuj24/TtxclyHHnADj2OCRChJxs1eRYB5Anlhkhaxz8DMDnbB+B3Ixk
BeztxaAKyThv6n5Tgvb+PmsB4mmiTPld8Po0dho3tspAZ0WE64cvj9PhLAhn4VZm
+sye/xDedeEDe8GS3kcXC22D5pc6aiGZYsA2mTXFxlhgs9HpJCJSoOtD5fzwhl6S
/fTZeTpaVPhQ/yUIp0vlmJFyQg1jyO4wfyGPEpTOHOqvL9sKdxXgpnU6FKwr6fHh
qTgq7U4cYM1jtFNxfFY4KBRsbsZZrr88wVY+4Ob7mSWrubJurRmsF5WW4UKXTBD7
0xo0lafdwZ9SOweQ0ulJWQXYEGoPYJx5Rq63aD7lztNXJIGVY890MY4miMLFiLM5
FJr3d1dSELtPx3ksZpBGhTTwhdco/B4FW3loY5bKzX61H040OdBw5ZTZmNSiA3OI
qYrVleiLoUkWXkoGi+t0NcdJQCIehGQA5TMVd0DaH4E4ZhppwrDCoA1JKnpgHfYP
+tYS5MczjjESnIIrIajn7s6bEHYbEeHVpcJ5DjiJMT4/qxvNTx5i1EPdfgfG+hlL
2yIavkaZkfZokx2W7CUyizVHv//sLOSdcGV2UCt6jzp1zSMHdYt6p1R+igliziH/
AaJWzpvE9BemsTmrKhO6zGIDe2Mg+YUomjtT9wVex6krh0RgwwRMntpJbx2bm02R
dFacJOX+zk+I9XZsFCrH/I2ab+MowoWxn83uwZ1uvcwkS2azKiM6D1/AZzXqpt8K
A/TGDlXNrVhBWB81k4OEqWfAZ/DmQKFIqsrOD75SkwdkkdC1fDBOmPQSngrA3HmZ
js/L1H/7Ifds7quT6xNndXKmGd4BSnSAYzLcMOb0EYIJ9dsINtnyBbJ0OXCoFl+g
GkNQODeMKfBYiOZ6ZAzdy0uEkKHYUoC/KFgcHZCcCpbLy4hR4XURsB4rct0uWVx4
dvbaSPtUDSlTjJCBXI0FvDngwsjWt5fbeYTujfO9oKF2NS6EullVipzOTrR2bz7i
Kf7OpJdEvKicGn8nrm0UKWWgaLZEzzIwSfnRLAqx7quo5wFk0ewuim7po5iK3/Mn
gLvuZlAit2AnTV13QGj+gXQrF8Z0NrIuW3BDheWwB9sTrtaA4LjyCj08cW2rWdzS
DoEm7phxtQP2nTCCXOh1Pw72PPl2DZ7ASTNpQ3xPk8ma9aF8aCNYjLAGWsVSN2l4
IK7amqs5noh6qM3c821DEWOOTYc5ts8NOJTwV57yXTQtsfhWh1xCRbi1PTWKXuBZ
7WW/5AUEKujVRL9SS5GF1ncXIDJ3jBsbg9oIdlfHNM8ZgP7hXQquRJRA9t2VSotR
Xx9OfgMRsQA4Z4OEXjD9X4hxPXZdZXAYZODOM542ApENZHKDC9Dz3NDMj569YJdQ
V/BX56pSXoh7DYctA1J8fIFyese1bpf//WW9+fCdq3QEkGqrsi1qohiIQ9G1UEmp
LLY25YgdxoN1VWYGshVXrikGfnxJATg7sc0Wly5y/OyxFwW78ObAyiwWNdVJdO1y
4J8f678lbN+OLETNyLis//V3R7zIItt3Ed7UZb0TxCVMe5/i/0vomOJ2+gqcpQAd
5Tdwm4hKThnEavO2YTIpp83lzeIx86B7GhuASirkt6vbNZm6jptZ2rfQwy9dMvL3
GQJMLwjAZjTANUUjGrokNwISNMM1IhXtj9A8Fe6SMs4+DjfrV6bkmxY1sSdRiwS1
AqZ1yAeuylQSKoVKEvPLpTheuIrV9SkS3lfy3TAhWRu91DYxE/Vg/KsJcxZBkb8A
Kpz+XqC2sfxgas3lbQnY7U4LtpYfa9RLkDxYGimlH5i+rksOMGi0CIXtkSLsS7cT
IV9eNyYBT8BYpo0MHVbOmGO+uNne3RvKA/bKS656urJmvn+U3qFAtNAXkFSS/bAX
Nb5pPPwbMnrGGu/iAmkqP8SsCZdpPSqw0qLrgNHh6OQYR+VoYkw2JFxGL0NFA9aG
3vYKcsXZAJVT+0nAJeWxvZFgmjL3KPHTXuZ1OVyrSGClWeqEmLWyivNX7avjs5nI
HO4WmZ56n+iEMDKZnq/qRJv0GCtscFwJNFefV7Smm5zeYJkg6x3q/YULSK6+/Guw
1sWgh1HXyMFmsLdQXvLkm7MrpsDpUMvvG/YE0hJtWsoqK8LUAIb4v5S5iw8TZ8zC
rBt8RZPM+CtEhd+m/GHufJBsrk9gN3ueA5lki4tSMYFvlaPpxun0KLCIjb6KIGx3
Df1pcSRbjpi5uyBL1CwXHTP40EDiwI6qNCujGFYePNKd8rwDZBXquVzcuepEztdD
cZf8DieXVHyTsH4QOzTWyjIgcK6BSmUv68YXhE656u5IBAPqpnU30AIS85i1npej
jdJTFmFWQx4tXNj3XRQh29oM+KLGMvmYr1Nd7YlZ1v6Qyf2eZUgNN/qQdTENJEY7
HT19bD9ORFsa8NxQ77ajMLX0k7wnW44KxwoaMHl4D4DEU981A4T7OsD4ssRhdV74
gRCJ16nVbDutMfazy7QKAyOiTN3cs0FMVeNKahT35xDeEIYR1CZwLbnYmr6LgXaz
XlDop/FEg/mwPRYNVQZw8f3wu1//bigBlyXU5HkpFhj66DJ7lOEmJ5BqA7dt1xOW
wD8lTl3VrIW5ZQOsZM1aUZfx11nRcFY8XoPDS7XRsmcU2dS9QwEvgx+yCd9vBuMs
6vYI1C83f4v5k4DzbYd33NCf83fVgy0qm1FvOU+rB0RZ+vvoNCrL2gQX0iAQSKWw
wTl8K3EqZEnZhN5eIDvr41Flsgo83HtM0qq2xaI+kSxFdC/LeJj37z9XQrWf54ev
j/ua4hKsOW4KhqpzZvTrjhD9Q6xF7J3KJhPmLOJpnc2kUQQa59GPp4pqrjIkBb3B
oP5uc8Og2l9xnzSxBjvQxrWH9yfIMb+sUXwsc187OaxceHohDnECz99nPu5t55ht
ty/F40HlLLLwQQeQ8pvy+kDH444WO7zY5xANwEOQgBvVmZOrURcG1JRwAVK2WRB2
jIro3bg6siYVXmU909Y4Hyji89DPkO/LR6FVJ2P65dyyum+Dk8LSpgKISj4OhGdq
RyzZ1Bneg1U6baEqu3zpdPvfH1sTRCTVdumxhiPFACdCle+Po6KTHBwy8+H2hBe4
h1yHfGpAj8zETbtwRvit8quHZjNXiKcW0e+F/duhncXM6RhRgHUdygpRxcb6za9I
AEAwpFqVw4NjWgnKl4Bww2fZ808nPBiFKFv+nO5Tg54eoUigMSqHLf5z/HyCe1lj
kuol4VxTDErl42XO8S80RmVISfnXfBtSJRTmmrN/W7I7hnuVC6/oEMZkzBts623a
Phgk3q219o78plsQ7CeQIa4foLT30WtfnwqYeY+rm6tHXvK/G+VmCGYDEFrtKExS
/BKH/3QSvKWXOQ563vaGjicEnvJFb+QTMNA9P7O99N+j4nYzNGLpWWOoGG/4vgJK
dszzjReRQZtwQUFZRrpN6pO22FvVg588ejWY+UycPQEPY04tcKTxiLLOKnwsu3W9
rn1nsPt3cl6uFJXuHpThXM1aKAPPbMII32uCn50+to8rYxVzn+jUoLjRm4YbFYzF
59IK+UDrp+XX+5/UGNXMQ/MvJA9dsynkVcaP0LuL+I8gxZBpm7Xi8aFRuSryGled
weSWxYUxGsvh++XBJuzSRrD1gioNWQnxr4oz3lkck/7bXToO9N5+nd0N5f0aUhRM
dZmLqOUBJ9lJOkyzW+D1CyW1JCEU6aDlQMXD2jqZTl+hR1PXlN6GtVz6W8iQfzkO
ecxlF4kFIBOxhbXD5xNAttRCvYdM4R6kmkYVjvGWt7U2KR7RLsX8y5JT79o3DE0U
7mBfc2cJKilbIZI563LPeUkZJ4LprXbBFCu9nAlO8A2OSp1alEqHvfyVJpmouNE0
CCuzoDxhpa7JVyKzUm7nNUxnhw+piODcjzGO95wztaE9TWau2BMaEdr5A0mkrfPp
cL3+ljoWz3AWY4PIJ6r2ATc/wTI2sPMTgdP+E3gJdlFrqXE2byvTEsC3UX3TYMiF
dEU/MvSP56ggRhFglmCwILquUcFGKIgh90BQtPg9/oyX5XW9Boi0ZxsYkAu9lc7a
0i2rWypUTeXRREfEnc932HR1B3GsX9NJb7RKk6Ys6hb4ntOHsPt0ZG28I1a0Cch1
egonPzO3m5Z9gafZoPjDSXEzTZ8SWaV4L9jayvIHL8AXeimWa/ghe+hCaaDT1Q7J
Z3KqUgpQUihV+wx0L6IcodOyirNFp5amJR11HJyizooV6AcmUWbd/uhEkhSy4cGD
kini6/CJis7HHsH0eAiNEXNZxqvJZtvT3W7g8A0mG4e/pIpxK43SN/BvVtfIke8s
f/5EyPEbLuU9NZrBZ1jBjN0Db1qS3otP4pqEad3Td1hhnfGbcpl5VE6sgkbx7ACY
HWjGNm7rI8Qht8YHPaP5yvTfB/FoZ78XSKglmtTIPzf/DCbKbNuWZyasFuGkNtax
H6Zj0+GJ43IRltafWxF90YR3el57oYUY6iHphy23Cg13rZgSdxzVovRJ+3c7j7ei
gXIhHzKd9/OVVa4L/x0+sriPrgHdHyrmwCOBN4AttiMPsOfDk1hPw27+98bpoURU
fdDZoqQLPHU6gLCVJGaPliavilHZ5QsRrCX8t08BIWY+8U4BZ9OWz2WNiAKuo3q4
yzapZOzFMkmK3fUtFHWTNDBCGYP+SBHg5OaPdit+VL/bj08CqWBBjlgoWZAoo9B3
66ddrm3HTCDWKatqNloyVhh7qoEkWTK4ZOYDvnhjBXeTyoDhHnUBlKezb547m6UC
BvMRRezgIrRUAuQJWrPp3056co4Z+pBTATZX0+vfgeUaU5A0f1S3UCm/jH2Ti1Lo
ISPNZTCyCWUSbwrFR8rI+BfiHKihWGP4aEn/JB7DU7PmDdjt+mgNiplsQ8TuZBfw
TRcvn07LVmWgi7LEJkYCyWqKDAAFsQVfUPs7cNztIE5EFyOCMeLPC0jS9/dB4oW7
YaKG3fZvRoHqYVyQe0AfZuBbA0fxmtr0FxJMjZeRs8zpJ3KOFG458/vMxfusvuzW
bsOeYLIp5U2AVl1rRhWwIT1Iw9jChjb8G0C4ysLHhE2QztiAifC333QM8OMfBMe9
T2mwCZTQZgFzJTBCVWOLUqFa2wmrMs/BckUxC7PSO5BR/2M4g2JjHg28UZ9dhMw5
EgzIlM6mFgj6P1/OS0HgYwWIFzOgpYpMEIqogoMee0YgKCCSrD09OllBUxV1nPSj
dcRO5F/5jmJdcYLaDgX/CqxPQAu6AbsSNxQ6cuIqppHCqEnmTH4vofBWFf21o2Gb
K+fY6wQzxgTcThmh57OGfJwUh/w4hsebv1JIDsF20Gc+m6CfEHWYeiXorITi/dwG
WAOH7mZu9122ipfFt2CD58Ycu0gLnGuF4l1oHjmpdzGN3x6Ce+EnLSKoeyejMyU1
JqUJSmekuQctrAYOboqQ2PoafBQAB1IEgnpaDqYpbTaFUcivsnBsGDW/hjyaPV9E
XJK4M9Edn7GoJby8wtTiFXlvzCIPCfVHBIYpAnDV/zV6tYvIWbeTSdqlDDjFMNcN
t9X6cv/vAPWdg5ipMTIn3indn21K3XR6AxZ2vBXTo3pjRuQdIM+wDrSr5jnt7Ztj
m3bkBDchZLHKYqKNw73G9Cr4IS/QRKCP9TLFnGJgyS3jeipq+qQwppkuSAtzxRfj
+QeAd8S9jOi5Yj5DVm6Hs0CY30mzInnASG13qVFPxxl15QQ/j14zPfpXHurmHGOb
YPAJdwwpPZl9EwmhY/9udThByPFK7SUWuTd55g2mpjqQa3ZpWxBuBA2iurD/e8MZ
Np1gLWxxWuiQbyP+bZM3unezBaPcA5ywQQymN1vOQAt5MGqN/TTP+8AB0tmn0Uxi
jyejYZiCv3+oA0JlDjRtKtJZZ/9D08C50h54IyHBxCFOim9KgIeS/co3eUgk3UKL
ChBXMH44XLSAsujNxlgau+RjZhgf1TFLnmy9J493iKMVcJGd2yvO3yqEQR9MGjHU
xWBDpuNE9aiZuFxz1CvWwHnDXTMY+qwGu+ltdoY9iH3SpBllk1JHhSi3otoQNeEB
5pjvPxmPVXHlF2IJ7rGx1kVNsaBs8iEuXp1nV5Cdv47sKMijkRdPX7WMEbYF2Nc/
DOFCDhx7oUrIsxnUk/8iFvz6VblNaXOkXv0jOL9ixb7wbiDaIdCOv0VO5vOt9z4r
8UQqzNnLfb4SE2L1IcOFIW7sxGO6Abe3gRtr3VmlBy/0Bk3ALBNIgY6ZYP7u+4gU
/XA8TJoSWzWLG+gfb7mXulINp2pf7z2icrlOOJ+JdkyR/3nwWBgXHf3qfXblUg78
vIygwWw2DJM8zBdsJORVm4/3qCRwfHK75yWnov0kh/QdtAi5kpLh8WTB6vKTXKkw
LC1TQBMKT/fUjYS4Da4smH/qffq+RrtHDZYJdvt2Iq0Gl53V6PIoqEYSG3LX0dgA
YEehvIlMC/6Zl2PBsCcj1IEhlEIJN10Xwt29IvijDakeHyqeF+J3Trs1iL7wePFS
3+Xm9Q3kPobkLMrOxUDQuU0jyKns+tmkHpqvg/ulWQdKzNvK12Odhxo5EkHIDk68
NP3jOzKaVoOgTJBJWv9aUAawcktcfCWV5RZ48NJdf4nGg12+XmdYGiTRINaphpUd
lNDXd2kmRBd5/nQeVQnIPJ8EsT6ArAwsgM0U1FtPVkklLkbDVOFD/HYUldeTHvzD
+CLhJdNxmnDIHfIsYD5/tg5TezZobH7olzfzGNw2qCAZve/eSA0wQxjVCI/7B/jh
2I3QCNPdFzWnrTvg5rPMAvtwOTbDyhSO2ZRFeTC+AAuv4bZNi86bO8k7mdyXC5Ux
7dTVNr2aRfHFPC5z/bvg8xyjrxbPlJO9kA/15LBhoQLi25dXV4ycChR1VY18cDxx
hoRfjiPSHD91Zof2l1jxlR7p/860Ygvdmyp/ymUZpquU1833VPo9R8zlYH7XGPAh
a1zzbNrQDIQaHkDCO1i9ktMmhHAuq3gVMW2/wrTNam7NkAW7T7CmxLfM0dvl1LIY
HIfDxD5cRs8QwYS4YvrZHc4rGS8xk9HQjGxNHOFxZh0MdeRGuoENfQPBohRJ9G5Y
sFk5KPlC1A8XZJdpy7NOOjtYj8NcldzQ8oCm/2MsD6ADNhoB0PPR0lHM8POfcCg0
xD9tGAWMQ01k4wYODcieocI5dQuf6mBJxTSOt7ifjbELoJH30vF6ScirUa9AK5zi
EOHIzP5FkvtntLPNgrz8pcCxRaHjebbtopcMWWZGiXBY94pUvWwmW1nI2BtTuGIm
mt4JS74D0cXNZpPDos9n/9FdssO+qImTAh/T6QXCCZ5iRGObOgqev6MPIfeLsU5D
6PLZsNk8E2/8yMtkPxz3DejspNrh47lwP35DWIixRCIRkxlmB4YroR8+HP56y751
NpIN3V9HHAtcHhVnXYFX4eXQtgdVuHfRuAWTQ2lUJ4CrI3V/ZkGdYq/zArw1aIS7
h4a8kSKi2aPoBcXEmCJ2U2Ckq5hnkUNg5vZl+9sAnbIvBXOsmMdea9b229c6Lz8o
eyx5I6SotBMmEhFw+s/7xdnCtJtQguVzBfLX4KaYTNEV2njzTDAoOBIZ4ZtJqiD9
Vf9i7PIE/X6KyEyT7xSvvhQryAWNMiuox19VllMnJiNAkpARbOKde+rPWMTrzCGC
QNv6o+XxzPO3nCvJTaAgkt82iDRNR0kgXZtmuWvYh3ZU2tzcY9/pSF7MQ5rSjp2r
YGRflXa0WcxHxx49OApD0tsTuhXtRAFY+djstq+X7K652YZVmgMcgCYs+Qp1z0JH
MNxKoR1uqRt8euIF3MQKtC21CTUbnVIW9yppsm7HcWwjTyJyGAn8xsZUeuQyPW2v
0DBMvB9jpN0grMYNS0Wk1akvPIFj0yWNdMYXJzR1yyoRWkdpBQ20nS4q9Upl0tq0
a9YegjZfRmHAae+PmNUkGcZr83f8uECs2POSeis954O2BGadAg0NAyZysfX/k6qS
mIPs9jAmUpr7W5W6nkdOuk1Sm0SQZNa24DYRB02U1it8PsCynhlqXeN8IVGszF7k
Mp/IRGkz3ihfJvwn31sjW+IKCRoJ/3I2KFpjA3sglW/dViYrccPR5+R4LZYyigMU
Tnvh/s50xWIktLm8juyiFSL4F0Y6UzQ1PsPC/7BZyrRcGOyQBeTReB545ArmsISb
DCs3wP/pJvHXqi4WB1jeIm/Ers2OQ3iYhpHUpIwrHw/tXd3SboZwfsn0Q/9PzHJm
BvA6t/RCc6VM9oFbgfoaSOv3+SX43h0csgPl/+jFbsIEIkz2nlROyjSv+Q0KX7YE
Tm88SAyMJZMO5KH84qIB1FhImRj1LHyZOtV/Gt23rkSgKi0+rzia+G89eQc2W3pC
NvRd4EPvMVFG/YVxwv/L/ebLsWqCMdPXv2jMxXzIicBWsyAagcu0/pdROQP+JXlu
ehS4qMuUkeggFw/NTQPpdIrRN14qmaJjqSBOhi4YTWjqpZIGS/7MFtd+FQGdb1Qc
G2v6wvnLgP0zGoYIZ/bz3umets934HsAHAgeNLhSRrt1T+ZWNib+6I48w5K31WVU
/L029YUZAm2y4HbJu9IkkIHpreDbsCAXYrj23e6T8825EXVVV4jyf4Vr8g+Ijrn1
7lUWxYS5oczl2gjFHw3on73k4jK6pfZtsVRvmB/nwvWbH8nzvDID1DSVffcTAl5C
KrFe8q0QytTc7PsMO0F8juCAPEW8Ngcuj7xDBblyXRmsZUA0BcZ3mdt0Na1OOH3b
Gda/f2miNSEuQuZO//qukpdeA5eYeAYmaZltTDaMoqOy5GxLTqdUU9xe5Rpt+vDi
v0PrGSWbWuvBQIpPGe7jHN0UV7CAc8DhPV/CrPLOrjhroR/A6hBoOtNA5SRI5/+s
gFFX3vAP+UcniP85DQSx8QWO/PfMfYuiCymT0p7in/aPFyeOg0mViABwdyFseTl8
u0zyd+FP4fpxgpnkj/qPEvyYeMVTKhHgXrPGn9rppvejs/CtBwfdYmEV68Xzrghd
Uzbunzq+tcDweNCs07ADrJ7jCnuYxXYKSYl93zdsTo0h+/GB6WxAf5YqMvD3U/U7
SO/ZcCyJECWeWH2YpfA8haEECNZeZvXQj/6/8g/rJ9J4GQcDSO8dGmARV/ArYPRq
HLc26uYFSOtuk3UOPmjcERT80L5LHXjme9YYqzTSBAOs/0EzXVpHvh2s1c3J7jrj
knFLrdsUB97A+p/YEgfSvCbhUDyh6LuRfX3gFpB152iCuJL/JW86z6Ptg+5Sc5LL
pwESK7IzRTUie38PbVYS/hT9guNecurFNpGe6CnpV0WONw8OkfHkQCTqY1qV89mz
omKwRHngmi6v/S4uLLD5FhKjHDH7qQI1CMcVILfxmCxqpCr04Wdpv4VQXxEBV5gf
8Y37tPZBjQstfJkoN9T9nFwCzR84gSYoYw08p+o6W2bpwwmfZYcs6xsimyleTksi
q885dP5QWEDi+qL/qowECyspvz9Q4adZqPlS+8uZ4xuakfilKWw4yu4CMKKROAr5
GlwnDcrABZo1Xpe0KAbbDPdAqwsqh/pLK1Fq5GDXejNPi1KoXXi2AFmG93sqT28j
87tVmk8YJqJnUWORgWChtKk/1C3I7/J/ZF/wn8nefSkF6uSiPgX0T9ZlHoMZuvUE
3pxT0UtiXA7VZNUmF8O3MqT0gotTrtPNiY2niUbgnEzrcHKqJSdQPDeIW9TnGO6/
XZZCeN64IWuZAX2LAuUudP2Td2ytddfcsIwgfLdDyDfLoLIAg2I0uIFYvhMQsNCv
teqJhzWnWgRCh2RnSV9a6Se++REafS057+Q8EnxVi8pjUUBg1kL3HamGDAU1QA3v
UH3ne9RBEMkYx5PusFLyYMItjYVp2kpCHqO880UXHCskb56PzipSr/y6FNhTwR4w
yriE0fLT+Sh28Do2wiMU3wshr6THjFBTMn5x5KD/YDJ7syOYCTdZGWBVLspu0SPi
myU6geNG36qDEBNbZ1lWFJDc14JEk24BFZ2G70j1ZFIGmtZUPby96KtUReIKoQID
SXRxwIdeoq7Pw6uKv3hZnC0Xxl/+DtC1PZfHH9c1yFGUHLpHpI2fWh2weet3URz2
FnNhYpb0kABVsPYLHkO7W7AmPHkQX53D7BNMD3AlmksmcTTziOEgH7DBF2AO6N+o
rWeCZ7SjimIULvG32v4t2zyq9ll9298Wb62xvRWhkRLWd8rG9aQBZhEJ0ZLuSEGj
G5tAz7Zk6EP4lXrCMNp3zadVMUuRrSxSX8hVrkSMTZH/EOn18uEmWA9OiwVWAs+s
EwY9CJLx/kpPQNEU0qVsUt3bOwwJ/a8abo4Kursesozm/DgFrZrE1Ui9FsLR/SEf
CxMnGCCM97iTztrOKwYZPnrawFg8Km76fB1ZOJea8Mk6JkxjbWDwC+Ihjc0Ntev/
M2o5NgcXFj/Lb8VMEDqnpvo2xrgQNbowipS178T+TR2/50sDJZivsxCCte3UBF5W
4HCnjQY7jYG7Z8COF7XNDAAJvH955/ZwVg5I8NT+zxkgdC2bsvEJ3VryPOdsT4TA
ZBCL+PTNdAv/ydcZZKgWhrIEJ5VnPuZKYY18JrIv14VI1IytFte6cl4TLFqcz0TL
K1MBwOSZnFcWlyXfE50mAWfp09HMBLz9+V5sDKo1JmFFHH56pUw5qAnlZclxaZb6
pGtPJWQfiPBnZ4zGoHZ/PxiT6WAqI0SMN2q0Ftev3Do3cz9wv4E1FgzXxg9jyElh
/MdzjSA78aHdORO/l+0TQVpEdEFWLsxowLP6iCYdrg56wwbK13ezAbAZpQehItaT
vP46UM2pprjmcc7n3V9U/mRHaKHZJ5B/VcUslXOpkVDqE8A6j9AEL26ymGeW10l/
4gbf0nNTYQojciDv/UDs5uaVSyMnLxrtqkVBiIqHNk+MnjIbJUnCP0P/7RjbjO4N
N7c9Ja0sCKDRurWwYor3zNbK0jpD30nwzoDHdjv+BNyeCOwyHjbf+jIKrNoZGDpD
xitKi8xOZMJ2eeRlkss2ZNv0EGpyipfVjosX/Cw4Hy6/rUPHSiwEKSGMVyhl0P+r
sd6uQi5eNPs1zF4FzA04xcSydXV8V0wO4GRCuPeqvpI49aPSxcrotdoiuV9D4ZgU
3KhtUFVLGDdGdELje2zuAq9ZDKu63uJ7JIqbJRUK+zXKmpgL3EPY5wITeVZkQUMK
wNTYSDYJ2wYXYKHo+RjPIp5mouvvlDJO9ksns/vDazo80GRthLu88/gqZB08GGWm
J2XFo126Et3JJ+sheR8Zya6rx+n7zeAaRy8mQvLAY3mPaJzT10/ogeztdhtdqPEc
K5VDseZ98x/0OkPJc1P3AWaCd3dtb6zvAOnosDXybr8NOuGCnX9tac/Rxjrc2znk
ov7ZHB3VNMHhSSseT0OIJ00gLw+fQFlg+K4dcK+Nqc32YByheXvqb8OhMSmF7YEr
IPRo1LEDiJS3nv1vvFh9UC+gyjp/iFPN0+lUb+/Q7Kv9Bk2/DevhdjV0f1EMuU/Q
C3lJDYYoDoD9KDPeU+mbJb5Ico1g8t5i5KAle0+kC/aBFFuOcroSay9Sg3fazCgv
HFJ2E8YVK2V1KE1aUBV2uwDWHZ6WhvvjvrjqAV33cvrgQLBk65HsLvMspyoVsRFI
qxBQwd1m/Vpxl+w/KcYHF3flRrW5ykLz4XTCmLH0jdiFnofDOg2+MQzSAWOYuSOU
7Iogn9gSj52HIWjE5FvPBVCZt9Sr0aqrPvoFGatI1Y0YnCf0L6SPx9Zi826bKRD0
1dyTEla1Rd5GV1S43IPnXBUTuwsZD+I+4f+v2Eq51VCXW+eFEp+CaWNdhoP26eD3
Hm+J6rhxd2y3V94K6EXXOt9/jLB1fbEiIAgKbDxED7h7dMLdPj8W6Ki1UVs9hqwj
K8k2Ld/eAgw/W/3BdSRcj/NLztpzm77qxGodJJBxaQD945RmXJfDeiO1bbTe5cNG
qpF/8dQJgRzod52zdQhwGNmjsbqLVq6BAit2+6n5W2xWsoyjq1qGWisgeXNPSLFC
WA+9RnNd4MzxHnfhruN8bOjl8xDPJ/Fc4qpj9nbTb3Cl6KFQQemliSohbAqtmG5S
GZ6DOYHjlduCPmta0tspDaGyW9hhPDVGAFeCd+L95fdMqQur4zUUYMgOR2IHFx+p
fNEtAKq+ISkrCdoRI02oVOXWtGHy/XDDVr3o3GQh/J1u6t3wbYkYcTlWH+RqapfF
hNh1oA1qCXLIN50dizBOsu9qoxNaNqmR7fMaf2U7IXlTP9z9S0FpeY6r9Szn/Jt/
jPTYJB7uLdR0KH2TdyNso5oAWI1SVhE27tb7TVFmdNhabVn8m4Y2DyplkPsBvyNE
mNkFlznNcfsEYzPShvSoEOcA/466L1dIlEX1a0X8VcvDhXKzxNRC6P40FXunPrwu
on7kE/9qJLdisTtQhA4u6p6X0zLkIBQrF2BJkHoilNcpG9rX9FQe2j0Y1suE8bT1
Xp+anyr8NTJqNbC5P49sVTUPrUgb+a0A30sBKLOZNrxgkl/nXlN0JO7sMCGMH5LP
dPx3LhAvs/7rre0aHeCtvC/tXocD3qX3TyQ8LsTTN3BJfVcPVGOxg6TTIpfmjRJQ
JVKze4BoyEQe0ShX56/PW3GjqN4x80FhzS1Us7gvLhMupTDbbKBICOcSeQC8+II+
2tSWG9yiC/tNlR9o1kuUfUI7p5LkOWFVnKXy4gx32RHVg7zvqGjiUL5ShHwpdGpA
3ZP59IUH1XuXV+QTwYWMFs+RFTL62WQFuT4ir1Hu5Rg9wMVdDAAbbCO5WiR9GNRP
lfObKC2KTHmeaGIGXP4vc85YNROJFm6tzMjPqxfr7SjjBkqWV9R/GTyOWavncB/N
5YtrcGipG5KDRCaKdvTReqyeGeijd5jW0aK6vdXKZ/IFmd18GWe+zIpZy7S7KEUu
PBSlmHnprUGewoNdC8+b9egEkKbjjM3BPGGJyqC8i36HOyAVi9BpT5k9Wwl0mQ2r
aC18lzRA/Im6ovQ04mFRJvmTB/1sHJ+IHcoukeJ5vWpj8ZjEp4fvD0+tg/0ylvjK
R1dZNic7LuSycoqKiV9gBsUNt/EofmNcNy3qi7ST8ol1GIINOZn0XrvWPYYgC7Z8
f3VDmfOBjRaxIZD/O6UEOE4ZTbtNHRhTG83maSSpwOPYCg1AS8xdJ9eAKRROrNcu
/LjfgO4arllttOh3UJiWy80sAlMKH/qcDjRa4PWBra0m0AxXi4iLyVqaOOcK24Es
WgUhLX/E8B6v3FP4i/2ngwDgl/Grm+Xy3DBKgp1OsenKnbXBuE2f7tgUOpHNb7EN
1hvLlfaNQQmO0GGzQYn/EUahHBGsIp/Gn5nSCKhZrGwNU7dlS+d8ZAXshZ+N9Klz
HZoDYLa3qxRTsnHeA/KR9cCTVo/mPMpd1EQIBmLbrJ/Hph/5Phc+IoEkv0L4sy9Y
ujJHcKEnIbP5veY7iGai4nU2AH8Or41koQpXTPrQOiz8gZPXnLt7DaIBOpW5t/QP
Nq+vlNb4XHtSJIgBjdGU8WuzOL89kmkUG4ccebOu1mq7EsgU3gYD462NvisbijrS
dSmfiMxX02Cx8L8PB59nQOx5GHtAFj08CMcuWcjZZFy4R7+fq6raxk0tki0vSwfp
3JPmkZcVnHTNXDwTJtdWaRs2exgjvdaqkEgLwOrQzYVp0jllphbC8/AtXslY/SlK
QsapzgZJAJBgvl9Vj+EhPLXgQ3uakxleJ0AZB7Ma8sn4bnDKreN0GHR9EaX4wj9q
COVqaTXz4wcvhGC6h5KlqSpmCQN3uKqW/PxAVTDbVS/Ee7FCtJITKrxw9P8mrjhe
rDYbvlIE9NqVbcpV4hI5sWlOyUkDA3Rvk023+YlALFZC4UbsZXIPJ2Sh0TkPCatN
aHODzhUW4umdEFOBlBPB8ASdi/On0NpsAfB/EUxBawlLaasa0UE4UIeHpIlIShxY
IN8aJbk2hlEnvTvn2cTEdnnNuduSXuH36Iy8pJGht1pk3BmkedKZumngytlM+eXE
uEFgJfdd5dtFsnB0aZE0eVwQb1JL66H7Iek690LD+Hw52s8K/NFxhTXXUYceRUf/
k/2yfxahPgPPPPPH6fAGmNNEhQz21IDt6j6uJPQWzVcv9mYiNIpHqu9b5rFrnvGQ
IgTxxVEIrh1OpsbF/QvcLpAAQrb5hIouXD1UW/dgN70JxgGiNk1ocuVIynh7fmae
7NI4sMjolk1fNlDwHwBEXl5RVkv3NvFmM1q+ylawGAm5DewbQaKva2unNuQSmEua
4RhIDmZj8kiIhwzl7Je8ATkfEkp14oWP+BCJHcQxMltG37MKksgjRPN5O8DvHAGg
P+4WyxlBCdHpaVEWpAkpMeYb1rKj/U/sVyuCZBzKhcLSn1dhd6RJ4VUcba45cegZ
505UibjNGUYc6yEMLZbc7EZbwWc6AlhC24KffkoaipjORK5/qmCibKwpFZi2aM1O
VAMp++sU4ckmzNA4cMV4mlCDzG/3Qhn3nLYiYEKwXb+w4NwFi6GesU/lHCknGJFW
0vmhYuZnbOC3WTRTQAfJxEPHBcEzhUv8tZpklHvZGGuPmmJNxkWMKnfd/vMEeFQC
dWR0atPGKaDQoaW26vgX+qMp5EcJg4Qsj5SS654kkxcrIoCG39MOMfl0saoNxP7T
Jpnthz66Y4jEKkTV/F7l2P/m4yQHMixDaL7IsjUeBP0FJQsnLGdZ6SEBhQbRDoav
O4q+brxRJLcE9JuUliUCIGqFr+eE6lNURXqv3lN882vHmhnOWPxcD9preGlhC/Hc
wVAkhdke7jkRDu93yMEpCyFdfxIEQOFSjsRnD58Kz8XQivtocL1J3EiRpF57lTol
WCKkg2ZcBcDMV5yYy04KGNPUvya+6iGfo5QVQF2ogpNMDkgJGU6+/zFZBu5JOxGG
vaV/U8RAGuRD9I6A+0CHpA/IbA3fRsrvt5R3+3R5CPCVoQX8vSyl4v5r3UhmPMog
81/Hp1VvMYmGxqaN447pKr4dTR+SzfXulieZZH9XHwLwJ+5aOpXG5ZPN5G0u4dT+
GlewcdjkHVy5la09cVCbe0ljoYT8sIodAbdB/LSgny3+CMjZaj39vdpe8W5lQnLg
TfKtITg2g/mmG8+Lp3YSltkQ7Wr8yms2iqdhAsy0r9Oy8qVBpTFjtAM/IloPpLQF
EyxHf9MJpJg8dbhmFBcefthEKdytW98R6fds0El0HCspGLz6A0TBUOc6G18oMO96
J6WDc5SNxJb50T9SdQuwfMCoagOb4XwUG5DHz0u1nXx8OtoXWMm9rxVQfQxcGXsN
u1vDggNa4W94hGWVpsfn8xHGvib0ijLNAVuvcZhV+SM7fji6JTcepy6zWXtJEqFc
A6MUR6BugrQdw8grXrSY+C1ghfT9ObEH+qkvLjlVk0bkMV8S3SPgd3sHhd8UT2qC
ezX40hJ8U4KLYfQbQ7FgQTHnPO1PTQs4Gkopb40LMZ2PAPh66Vm0M/1J2fBBD9cv
jaOt7ouJGg9KB0X11Nn6RK4eSl8RTIucs9ma7igBpswkFvH83e8+kEf7HF0RhXse
dcHRH37a8R2m6s2SKCNj9iLWCFdop1aziry5QK9QdG1LO2/lUkbPLNBYNFVQA2NN
d1vdwkmHjkVNXn/ayU2jyZIleU4gx1nYQSEJPYqB1DwRO4A1frokW1Yx21oCNPlv
0/RA5rXsKgrbRcO88K08vS9VPrPc3wnFFqfiN/LhfW4IhuIyOKEx4lyUIt2mbsDb
bwo5nR9sAk7s3LORKLMI0gVKJRiZ4hcShBj8JhyZJgRrQg8GqCDge1qYX1ievlN7
0dDwMzNlSa2lH1YOMM69eOB5JnTolRmhTY9M+GPesjksACAc9ADUZnY89mbXf4gc
kaDZGqlzczbHB9p7beYLaeWZPVbIKykl07xDbtzNLMHa9nKI+AbasARRut+kIMfZ
/6J+c21pwj8Jfch59TY2/rt/dmK7HWaIXuf1HQRKXRBC1xMLc+KdNx4zE5//ANVS
Y1g8srEvkPg6ZTRAiREgI++WqzeQdm0DicBoaI4dwFZfhXc29EhGyKs5P1OOxKbu
OJZVtCwHR+525lBJmih8Nnsf7j1Ym1hDkgVbyGD0t8/lko2+Ffe3EKhUg/Ubuo9Q
naaxXn6+HwcTQc2nBGzmktX9DOBwClGDpoBA3P22svSBsOMvmD+OW5RyyVRaj8jQ
jswSdqSyd9Ku/9ajTtrGD/kHTCq4cCW6wj4nAGwK2qo+FmxObQBe7syG9jX1WAyM
cEMuQ+4UYFs7DUOwsNMO0k7rF3MPvo1Za5r40sstcQcbcSpKl/wVeuVmPkuzih3a
Mmu3qYfd1aZt/ZqLikYfmrmXpiT7lasr1dJhVz+cH+mDKHdZ+OyCftJUTaFwVzNW
DamS0CE9Zw59NN4OOfRT65bzfWm25dHN8ill7WC0NdMwmx96DtNWlY0MMZDy29dZ
hqO9g+WCGlHzwU9CAqInaJYQ4YnxrlcVSDR1IedlD9iUCkflRgnFzHDCTWrsvlGr
/n2bBZOyB7xwqRTOes6R2k+Jv7vHym9fXolOhHdi8uEsaOAvsdeyr+opUdvIEt96
AmemO78sPzZC6Fah30gXJGpTXiQL1OALb46E6xZDiAZKVw8uck57VvdV5j7cqfZP
34HnWzbKz1a9r+iOTRM68OzaZkLKlj9Mzzqkj4fyNM7TKzwlrJTOFkjSzzVnHDsv
PlKba6YVfWlRP3uOkZG9CvYDkQnUJvHZlHeiElXnPNqlEsl5fEuDDuB83AmJpq8w
Joq1GEHd2GXE4cP2HPm8lOzin/qYCDYerwaiVrympOfP+v+bDJXd71Lu79eBFfwP
DC+Ty+TE6iR8Jc1bq0ZvhUs8GtggGm4aqD9SDsxcyJvG7/Eh5idgwFKX8e4sXAjt
2iJa8fJGA0wL5e0qXi5pqpaAWwnWa9kVVcglbxxnZJ9lVbZQ3DAqyLP4NUrJfJ+u
aGnOjq3p888hcvf1XdI98AGkEYRD9R2v4JmBpESNtCxS6Ph/zm4D7a7y3mulCSt3
vtgy7thCw7Z/VCYy4kPMx3LascIOM5jL9t4Y1AOyCdnV4yzHDdBxCkzX/hnA4D3h
6nAhGmxF/0Gyf9jBrCm/iYFC1AufKGHCymrqaXeu+G+e9kpeJUnRBG5iJxOWV0OF
jgzylhSzE0UNjAqF9+0oNtuWi42j2z8X5hKZFNGsTEgZfCxHy6LfFdel1Kljw7T0
RcQvdr+tKyyz/Pg+5+fnAT0gHDujgSrMJPpnWe4YSgJmhFHa6oae34UgIcJnTADP
kDT/cJ6KsCDqVPHMr9dVNRllpD7/4VzJAcboT1Woq2gqiLnwsi0lDW/ZPwdQX+zy
qDK7nl/wboZe8S01J4zYciMxX9Ysjw0wjXXB7nZj8d9x8c9zGP+FQJK8nl/Xe2zR
/jSoB68IMvLQdmyn+SlAa8d/MR9z49bYEgFV+ZryvhlwNVMKJolxfNsqSlrJzjqy
axERBj/CHmDwYWZqAVlK3SAYylJjd0fJphTtrnLgX1WMNsm0Epdc4oohoEhmDx8X
uVS6WYPKElb240EBSjrzNhPvp/Lxp5gG51pcEVLHoSuMiiAePycmIoQJfTinCWqk
O1htVvAdZouApvJziHVfRrMObr8XQOwE9PPsPndfc6P2U50ztAeoS3isPVVWRLI7
wUddSrq8NdqfHSqDe2632XN0HtjxQGtnQVkCoiNk4qTMz8QxWFJV+uFXJfj8wDfn
LiCVd44t5zI2InGDeOq70DhxMVeerv4aJgfgH9O1AyQ4Lp7/eqUZJltU1UzjYJBR
maq+WIpTFhEPFAimodCWmAqb9hYHzpIf3os8XjOEaRRjmMj6ua6UHB0Gm7JaG7YX
3ymTIBndNaPsKJ99bIgG+193RWLAl+cjF2HzQrpxGCwNeGBAk9sToxB1H7oPYM0R
3UaRRE1FuVfa2RxlKlTm/icrRESUd4shlC4NUxAac9hgD4mOfsgrM1IH8jLlD7Y2
qcfQ8b3BrdbBkJIIjSc/gt36tRjED46Fq+dLo7pN0aADBxg/pnuy4rsEsT5VOJGK
8iw9eAXlqR7VkZAwXdAjT6DmXbobbMjTPCqEtXHCDaQONrkO3V1IJi+zp+Ch71Cy
RAIqvhQamJYqtNhUtI2SUt62ngmkShvsNWsxOmCE/eQWaEncYuxw8jGSUZtddW3B
BKZhbEEj80Ookyx+6PTqLXzCkB0p8TAQjcPvKPXekvq+gAETHYrRlzJyWWAHbn0Y
aWSzFAvz55iAaWf8+KFQ08D+8vrQnSA/S6l1MePwprHYwxSD7fLSF6J969BHbH7P
7EEIZcZCVHsynvJTU0vrVe6emn+aREA4HG03SaRmKScwfi2KcgrsUE7lACW6yNf9
jFPTkHiWJT9coW3vKpa8tFh6hfcmvDCZqFwioO55qbDVhA7IpF2vGBbyKDWkT5+l
8u8rdpkfucXh64DTKe+8kbM0t88h1YgjbcFTmUE90z0ehNTY0vG7IXxUeKEEPJQ9
4AjHxk0lV+O1QfiDrdJucIuYmMQFfuUrrG1sEfh0qIdr5GQ8eaVRt0XTLoaLoi7U
8Ipu709CzyVy+oj+6v7PTioSXc4OPnkIjqz250eZfuq5JYKIDoJPyMNUMkalB6cl
MQZ9xYKGc9ahvPYZpyN0mFdwNc9woa86yuEks1BXLHb657dmo3quagihD3DEoObN
52wk3xNmYeFdR7MBHL0zCt/XTjmIr/Qg7rztPrBHhbZkYH7dLUOsqiAjLwBN8cDj
wvsG7kg+kIvrY2txu4HWNaacICrKTQDgVY3hnG28Ug6kd3v2ZgdHSFWAB8dll39d
B1FT8kAjSVOnx5OAcJ12JwBSyt1RlZh1u5w6Lkx3swqywEz06NSCKFDBGF3FCJbM
51tZRL4RXfr73C/Of8DoSl0eDAg1n6VqwF2yvpseaZ4ttJ9dWYT0Qs4nPPh6FdgF
TzEJKC6wS/IT0nFtY6dw+wzns75aBW+J/HrNVn7pxNZE9n6b3Z1RBYog10z6hdLq
sHKBYUT502JY0c0Z6v0OkmDr0AV0WIP5DVJarsdmx3xRUEtbzDWJeKU9l0p9x8Te
SaqtA1CnQfdTIsOqZgSmKs5IG65i5LDOzIWBcNewshXzqsl1j7cM91D4FDswP9Iw
Vzr1F6LQ5usqA/qdULxJo2eqrLTEcRARPUbLdTUO3/vHIrUd3ie9ISugqrMK9BX+
iAtZlopOjB5rYtjoI5jFxuSHmHuKdAfT4PlxgnhVrRSYUUkgZbz6MwCXbYqm7WAp
GzB8hlbGiqD2uCbMdqWG4aXzrwZxE3gWvoR1O6Y4XIKPKQ0b7VpTTdFu4TLx08Ry
5F9M7FbZrQ649lOt5b/9DEg38RsZYSh3OLHao5OpkFAqg7MS2zYh3YnpfHMA/As2
18MSJRe/XS4+ljTjMXhNtm/6WgU33JBjnFhovdBRIFPwIgHmnP1a3Dyfq4p6C64S
xZ+Meg7PwdXpqh9EOKwDiALD8nMWqwY2U/n3x48j+bQ4g6okJ4sURwQkXfEO3uql
i0vuIJuQeh+My1axFcZ2/EkWaMz3z0WDGxOu72h5KSipfm0jGzcMGhPT1XnImqIC
1LNoxQQ+0Mg/oDerx02QaoJ2Y6hA0WbS6xZNdk38E04Vvlpdy4ifqbgq4x4Gf75k
4ZEeRojbi5cQJHrQhSxTSCjUd8ob/hLu0VSEB8NhJCAXWY0CPdKhM/dCJ1uQv6QV
uRFDkgIxu/x6CviBwKy+DJtiB7o5lP5pYi60F2UmLV8dtuizxJVB1GTKNTwLj9+d
sIQE2HimQSiM2HLrlAvLxwsp7PSq8yDRmus1PmziE7NqqZrYauoDo4tHR6gtIMdm
T6OV/Ft5MuAxNWNwibJ0azT2EGs9r8eOUTZ2V1qZOoFb0wo8T8tJD5Q9/maae7t8
DzRpdeOoaNoS4KEqsxkX3eTB1GlwlM5AwmbX/dFFMKLDaP16yEH7SeRCP8lTp9w/
HbkdbCYmTPm5VoM+xC8a/BhOtT63FJcx75tvO4R1PCpczh45n05ZM1SBeJ3HM/KQ
qG0/61ddMiVbO3Fq+2hqXmo3Ujb6lIdOa86MUshvhH47IQmxahVsJWeoIaLiQcge
wMwG2WZlBXdiv4bMbwXYaUOKDziqvb4OIe73Gc4NxXdTcVfeqv7xp01DmeK9+vP4
fJhD7/2hdwFWrnrP/ilaQpmUAfTTJVr+jEDbSQT0YldIlLh216Rdhz8W138T3ZBJ
zQE1R4hOLXjlhJnKM9y0wSDYzWpZ7AvTtr44FPISis2WUumDz1TR0iTzEyrSqYE/
yojj95O8pbTVtwpxSDGm/E+NQy8ZC6u2Di173GZ46Jx8IUCPjYPfLynvE60CLRMq
K7nclO8B4j6+4KQ+oa9Y1A5IrHXkUsJXvJAhzQ2EQEJFeeRJRo0AtPdM6hcJMmYD
0DUajGlnp2iGoSk45OtFxWs/8eG2QeInf3L7yFpZ5MH6Gl7mkiungE1A7Ql7T+D1
KAmdZ3dWCf1r8saFah13gsWc1PI9U94I93qcGw+l5iBzlo2XTaHG7KPNyq9p7d0l
eC+WV9JHsk4Ow0rvU7oKNjWtCryuL+W0aGw2k/GtOWOLX++BsNCx8a6An4pLEr01
Tc/Mn6K18WwbgX6KCaqplgnaETMdcGi+5aFBi4dOujZdGz5ZNBWaikqHfJ4hYjHt
JaIB6Y4a5t0O+jZQswbWvQhZhsHr+LLXEx7QbmCulVe7AMXdD8jM2DJPpDSBBNfO
7DWC5S7NiB8wI88fVi38gLOMhH1i4eHnxxkx3edzS8Q44bsj5mIG4zwfd5u/mSHK
p7S5qWaFgvb35nP0ks0JtGBQDGkpc2YVNqZ9uzgOcBZmHogWyg2WtoWg089KGuoR
8SVTwWzeRgzYs6IdBxDItHGFdCNkZ9lTYmMwOhaXQNsJuDa//gV1eK8Rzn1ARtba
MSbGXS8XNHm6Zs1NhmDT+06qJjowxBHkxYFCP3L6zs12t53uy1/gOLN21sLjySdh
2CJgcclTyQVubPidzlfPHTA0OeC++SasDMunLreRfExIEbmc4dfNt5EHvIVT8dqP
SksA51zlG/UINkXC671/I8SASMXcBtfHrY2ADw+oVhJUghAJ2OkUUaHYlXg7Lo+i
4yd2KW7/NqD7KR0MJYAXZ24JO+knKcqjb3lTBGaGYr4SE460fuGsdVWj2awOoY3r
Xe/ipYE9p4Ev/nwx0dy2apufLbNV7Sp1t/raBzLLMyq27YC+isLTg8mtGCOo2tnY
sTUm6JCMVF/VvvRWfKbtrqmjRLiP3jvRMwu8Z5+Yaj1upfCLG44/aeeBCdGEp7Ol
Ei33kfsVtQt05j3WQNpTJI5z97knVadsiotYODR5aEEnsKXKBkk25d0Il8yE9PPL
12s/RtknW40x6nSMtgFKRhl/8E/IeCClPqyxYu1FE46LU1VfBVU5cys/neKmqcPn
jSodcPGA748QC9F4lo5D7/Yp2LWtoc5PjxC6XIzVibML7jqqgPcd7U9j4SCEo1jK
XbvpjjSu4eQYrUY/CALFAG3Oh4c4825lsFQcHY0s05qO0mRy7k8LVbXSrcvwkIV5
w8iOVux2ubfcyyO+EQq4yiCsYeF72mNSkVI3QYtrUraRTHOl0hzPLfa9i5vOpMDM
pfNlxhm2PkFzb6V3kFVTUSNXYWmGwLmXgnRA0LefkA2W90m2qDL2pwitbIqhnoUD
a4naGyMT3OKpg68FQJmLk2jefwfNa6vDnR7gmurgYza2nfJsuc9IR5blVxvbSKu7
a64U252keIpP5ISQieRnKOS8VWlh7nRI8l3aGdjDTbUXUpsaywHV6nAWtsKnpYRg
53sUZpl6g06IXyP0rIiQo4S4Ynpgx4GO59QTbA/5Ux/CtFnX7Pxl1U+obO+SDL12
UfHvymC6wl1Z9EFy24Klyr6RVttNjymrzkBlm/o4wa9I8EY3MAclEMJT/6Yg0UiR
WYuVjf6wffqCb8g/G9Aqyb9gZII1XM3fQaxhCM+6bQA96GHp/O6DBaqBR2zSBwJk
Q97abF0XLwMa0CFjB14U7RtPBPicwxxQNqOVqZujtR+B7oSLJmLXArNR0XdKSGN3
1wYLcjycBXWRCSpy9+HQBv18mVxXg5SDWDsUOV+uFu5+fkq8f7OCgJrz+tdUgxzp
xMMdR79s79bXZI6ItC0eyWNkpkBZ8Eaek3CgnYHcPGuA8P54wxuH5lnHFbuqdqcg
FfLq20ahpRnWytqK/C0+7PspbxAStpIKYreetnhmasrOUa59g7bdtkvDQ0PrRQgy
qDhqJp8DTCPsWiSEMxG9teqZ7HfeAACV47HODoLPXv2Xunr3ou+z8wNrd7BXaKaI
AASp/8MNm7BWdbhyjKkIzGYBG+TL1FsLs3Pn2ZX7dqKEBEJC8fdJErISGoxt/Pgo
YTL1Ktg0U5QNX/gkdWvTgsJykQHkXntdYlH8sZkhecoN2F6fMOt/jh1dx6Dt/YBP
vw8RdRxsOsjcyD8WHu7Swz46WzuSBXhhp2uCUHDoSyw8z8OaCfNwr3ysSV7YqQOY
dD0EJ7+W5REAqlVFMKpPGVIjZ282rDMn1HvD0PixNuOoZM6wgnyg4Niya/4Do9QI
pyKw6cMChIpFTo4LsPWsgTFoiB2VZPV0DuZtrOmaONZNoGDGVR5VxTeRfSoGZxCB
bZvqzNLvXMcSkrHpzqedYDjhEBdr8eZebet63KmjuNurN1P0V0ejTxsFMsUySVn3
Hv/8oUp8y9YXsvhMi4bxI/ma0MJMhkfRgQJ08w6GdadARiAQTQEya8DyDB2MahKN
OcH9eFvZ3MkbhM1vtWTNqCIZH0ytqbkaqWOPGlGuINnXzic9oTslLs+/xNwoKqNP
VJQQQFIrsMB0LlySGhYBql/kCJTtTmCMCcWDFmtbHgqfVHzn0sGzTgVwuT+PEpHy
vjkjULxcoqyy2/ItbOVCNPD7lOhBjdI6XP+t4vQFVmopr6ilOL1AqT+qurIIVsWX
kPoxuBeDzxFxIBjShtGfD6Gk3hmCuT+LyYBPJPD6TxyivvU7twHlaiDlDoAIlWOt
8QOrRIV12G8GDpQCICvMQsUeItY/Sbmv2KmZsfmVsawtYwZjRJ3h700Qe2F+6b/F
qCBh6i5HOCDfM0RW6vRt8p8gWIzj4DmeEGtrnjWG8JrqtWt6DUAPhYbMPAKXRlhg
UmbpHSYS4jHYA+cYXn9fqBDjqwb3gcWafuuIGr0Su8imS7qdx3BqL8KZvD+oF/hy
Nsn7VjRH+45+YIwl7GOo2oHid44LINvD6mwaNknahdPWV76ib5igZsykqXcvkG0y
Gu9lm7sPfPGHxtCaAAtKokOCb+U9ylPLUEP76dTuTqgU28jEQ8hvFf+s7TvIwnH5
Vivuix68g6mcNNZQBFmSTu1QrQ4uSYpGJfVnwfyOwioahlTlifFNDXYRG9a3JJOb
o0gbbAoCOtUKFmktaKkrCYEPgwRFNvuynOXNFD+WEda15LVBnc4ldolJLxdsj3yi
y+n8IoAXx8C7U6qqOHQNrRFzKxDhq52s/mrijBJc14PnA3R0paphXwn0Jv0keho4
NuMtgffn2KNIR+IpDmfkNIQCOOoic/zAXRBOoQOpOQTpQDQzgmLMiy7hmpakxAT6
q9NWfetTgn0XV6fqBZLAx079c1yeKfcCB7RKu7p/Kv7V2Yg0RDD9AwjAiXHU+C9+
ymxfEvkFYUq6VkcaDW6NYy+2A7IIVHHUnfbmtpgOBnXza61u8XXDHkIict8epoqh
UWDkpzhHrjEUp3qkZD2pr5LvPQB8WP/DCqlswzGnl37HmcnpxwHYrU4HNO159Rwa
RsMpS1olC7W5lBiA5nGjt8uRxY+2J07DdMqeI97h7vRnlHc+grclflKEVTw6gRAa
K5tQdbs64nSDkpVYtT8EqXMg+1n+0SEtFByy0/wwnlc2a0EPTzOMYJSLOQEPPDFp
YT6NhPe49raXjss70f3lvsVBUnbuKyt46Eod/Moet+AU1GT4FwYfpgBm8cINaO2U
hbAf0yFaTc8tUI73goMfdDCyKKZuD65LXL0qcqlnz2fMPUcsglNljBgP2Mg2nDtC
WxAysMiMmA10U3b3dbWNZLNyTTY7UsxUkTcAxluuqH+NxlSs52b+NZxxMhKn9lUZ
gU9CSrb4PHuJBCxr0tacVbUEv1zFV2EmPpEelT6ymdsqEFDOOJ0cDXA2MX4jyQ13
B5dFKWkoSLrX5zV9gn59roiBTqeVym8qfkMGKK8cXKbKl/9zUcMKQQqjUj5C010Y
cMJVdQA0lIWkdMRXKabiOtz8SoipTfs0zQVsLVDdcGJE0l3O17IuLudXehLrikET
nBTOLlfhx6EQg6keSxAlW9w9qJb15yr5tWaqw55aXWSAcsDAD8BzW6NTrGr5XviW
c7WZr424vhQ+z7RrNcEw7NKWhYKXAW6/8nwhiVl30CKgx/HBOXdxUD+AA56CL8kr
sdA1MXsRBAe2FgeGBokVrz7lLRW5Km05Tm5/hNin2E1d0+mmzw7r8b1q73X/cu+t
SXXofpNxGDXxew8YlqCo1QEKf2b1ilZipCn+dNojqIIpuj/Jpj+fie5DiUb4+HUQ
ZTfq15e8NjZIwE1ghai18P3MWap928Lwud4IDmcr2hSi7Ao2zKX+iQ5QG4BeY0HY
UX0q6O5ZzM5eRtbaQQc4Z7PyoIQJ3h/ISlLnWi/wl3BNs+pchd39siDwVf6Cz93i
PlL/zyP9CEvpOZzz0VAEZYTvwpMDikK1LHTSn2K2hND66u3Kdr/EM1nksSGTAFRH
lf9K82JSD+7GlB8rCyLy69aV6rNvwGbIq7i+zDF/9OQey4UGubogm22WTQFZdoW4
jtuKZzVHJuxlq+I53TvtjsRFbFTWIwIlKHfKvcS7YeOMA6UPyS1vpC2L8UAE0Bzu
B0z2SCc/njK7cKInrJmSb90I8qYMF7r2fLQ0wICQz0dSpBeZfbWFAqUFW4HE+DUA
dP9jlbwT/RFXkmMsunkZzupExyiFV7shuva57S7r4x4Wlx4TvWguKHq3TrvswllN
WTBGWGjwWPv3v/+i3Ab+73UDTQegzj6x2WL3T+ZDzHSxENtmNyHzNNia7gVCvW00
sEltIKL63ObCZ+UuJGaFM+iX9s3HUcmyt9oc5Kl1y/zMWPi3KdbNM937YjI6OMYi
QDIAAR+6L/Sz4djB/3Be6b/EzJMAIF9Sx6sH+ncZP/+4UoIuZw9mwuqt0DWVYAkt
StIq5r60o0EXvHKQacVSIhwC7CdRAOG84eqbssSetK0FjUfcHGpv/36pIUm9nKjM
wW+MLJR1Vd3dqAKPzUxkHIhGzY0Oy8zHwImPDdnpSg8GWXQU3XvaVBt+afBWPkQz
ZWkLkGNdCnZDTJqIk+4XvgpiSEa02vcMU2WaJDq5k7KQB/zqfauuZIbV0O9k8yqb
LnElCW2uHuZSJUm1Z5pHe6xiw3oVD9rIOoDnXzcXySoOg8aMMb7Er9GIP1skUgua
lS9AfWrTTh/IUbI3GcQPhc3uhWdXrDMBRjMS/EUMgF/Ao9sIkUAUxoJuqs8BwvWE
lQdD8DwwPyuS4S3Zg3OyPUWTmK633KS1bW5gbKCdGOquYLc0ohCxvKr1o5olYxJf
AuLt61O44liZSsyo9XA4dma1EHRQPGol0Hi1ayw7Mbz6Fy99NYv7iAIxtF+qHnfW
nK9FDp9mD6iuSzD9iwQph2aAgLX4ZxuBCdqXZFu/vl3lc18nzPTFalbK206rYvuw
3AI8qkHQlzWqHXQyOxHHq8gpYrRIFZODFUADfbt26RHmUtS1Etk1EzmQap/cg/pW
CeFqWHdT1H0b9954WGZjCTwQdKDTJAU6R1dyIXoWmlgtGONJErW8yfelTqleMUMu
iRp8rxnIvZ7MY+JzIrddXD7P44meWVI3DwVQP9A9cAM5grTqrl3RyXKIlPkx+RrX
f7HKPGi97E2Nd7HmMzRR42Nep9z//49aHDb99fvjM9sFNQ077snEFy4XTqk78O/3
WpkAE4mu46cVV/SSTEy0njgfGkE7+oHTSs9hANPAYchw9AkK9os1Sd3A++QEhSgV
POuQGxe1MiDjA8U+Dc9tW5QLWWiUzu1ShgwpDpaA6pqLmbX1XiidtKJhLigwvuph
GTfZfhj+1pDHrBkuzQvdkIgxnkX941hb3ZZRBxS0biVygPA4ZBxUd87zgsR1OUds
CMpItXvVhZd4+HQZXGk2Kd2JhQdzmo90k++F3g4/9OGmOMygI9jH3H+DCNGDwYS2
yQq5c9BA+1mDdKKhOkfht8ZttSPJWz7yevx/hT4v5YCTktm0HvfYgO+NiXBoorGY
qn+tcVzkhBcIXIGrZS8dgY4R5OwZK+e1F6+APc7OpM/i8FFBoZjLD1aTcFHm2nkC
box6N+DyuEy75KnE2vd4f1c2gFgOeVINxP40XRuGjEHxiCwm7DD8mGWs+917GEVw
vhjZpPxZSYGG4YkJg7Re8gZ1S/dHFRElZ5WUn1Nv3WXz5QC/SOGFDNEW0bqh8rEN
97+OEl7j6uqkr4zvMIaNX/K1Uuz4y7nLPPnC0S+sJ0ZezCiCD1dHXcIByJdjhXn6
YJq1pPySw5RDT7vOdMXL6tMtAtEVosyhBPRqrzmtdDCcyRtdqFPFZcXNQd423Iq/
cGMyLx9jeT8rBn8YVtJsoBnpGpAFhgf/uEkAGFJ52t2PihoK94h0+qLg6vZJmnF5
chbk17N0TQIWwVlotAHWVEsdII+la8VpasmUwv2nQJsDZjuxvvfLF78alz5pmPfG
UneQnGQ3ahLsyRHEUDpkOiCvkAtwx8nGyEjgX0SyB6+LOLKlilKd6i/4TxAMDBRl
HKHPh/PEwOqSI25bC7/eNVOzgvI+uiciW0+ug3nMdf6PSvcyLU7fA8EYdt9KeObW
z2Ops2Nr2dlxGkHaoktNyfx9DSvxzp2AIScnW5cq9/JlFdMlhpsu9W5FOQzM6o4n
zXozELdjegbVHPUIjiFI+FYcJuYN6oE0Ed3b0yKKHnt+e1U/aTs2rVKj3/uZSnNk
hzPwVF3N1fa5Zf9njiwQ1XuKpsQSiMHK+K/RaHB5hPNKi3/qfby2qRbpRHraTwh+
uEnzI5CV1EqmXS7vA4kvRwUrZce4c/+2pzHh9xCIjSxgMwWUTAs8i92Wx7eGufkU
L+VpznKvFlGtSXDGUcPCtS+Hv3cf1KhtU1+LtcFDuIXO6vIWh1Y70wf0+rLRa2vu
o6icXTEi1C7dHbu9VQJIs2jNhSmt8vaKiduT9LKpq6jEGPh08DkAS0AiGONS7Bxo
pKcNI4QtVb3dwRRb2+o5aQCEGY3b5yQSi8WORnOImlse4hA0ZtMQg8HTJ7ZptNhK
BwrJ318pBi4ybh90sDbJ0r5t/GsZQRHOxNjzIos1rCVrFYsatscMad4PgJzlNVf8
ESJyMXQG46nRFZKXSdvfxCD1anpiWZoGZk5hhzQ8HUQuDUS9+KqBAlpAsOtOjpaV
+7fDenjojMkbZK6nGemZEWN7mxzF4LYVQRDhx7H+/esUAyvlzsI3Aa3zfOxbpET7
tz+tIvXbu0zdBKxY5/jRXm9DHX6g214oGBYuBe2eT1I0jANzOpoXc4q+M8eM0men
ud2WMhPMLfrluPPVRBPdvVw545VBfbkzPhgzT5M0TA6ByzzK2h2802fWdWuy2DWT
7mx1hgF8Q6DurzfqxISbwQYkIXFaia0g2naJ8LyUql9UlHQIgS8uvlAe8o5JanaQ
orXdubZbYsBOwnzDILqEiYP/IQcoTes3O1DCwhjTA31URLIHZdy9PyfFsPjrVa69
dgSCZInMDiKtLGZGwmxUh5irb866kKLw6RswtqlB8LvUH1g2fBXPbYWp8FIzLeog
QUdM2eplkXi3dGMpvazyg9rtQCYe7tKoCZILpLsCJylC7op40FWWqzyLybuTqUlo
K3hR2eabRNKSIHstvUJHR4EqLuSR9OvCYQG6iI2XWrSANVPPFJVs8KfbDLOKKS1v
dmFAN7Ky54ZO+Ts7tCjm0JceFsUjl+M4NEMMhwMRhTlozyXaZtxd/GjapQ1sHu6D
Wx1lmYqcyIfe3F1LFbWi4oE24IwzVu4sIDtsX0wV8YvO4aJyIZPaVqpjU7gqk9FX
zI8s4avPzKuc6UYqm5/00RNyVcKOJjp2YYKC1fT3bOjJpp+m3cMgWZp8p3M61/1j
RiJNPQgvjqs2u9Re6VjrgUI7Ipo9Tx8R8oBoLpzFCkPheXVKnGcY+JRCObISmetk
xNBfU6EMM1OJKaE2rdjCErBKS8D6QsHGb2BdjH47EIFMDU/P0Fkda9Z8u3aSIiAi
DXra6xDFcGZ8wnq1ixg7UiyI4cw8gb0D+vk09AfooxNJNzgiy6npoxyIN2JCVuYp
7yvVsNARDbKHJhxo0OiNYS2yOCWQAsYp9JzIcdrUghLxC9vZYsMPXyhhAdfMDw4+
iwaqlJKX84gwZFbz1JzksYcST0WTT24Aqpzl+9hlmdShW9yA3RRbwJ9U9XiT9fR4
nYqAOPaOswJKtS8mU+JAgqdSKu+/CBmdkyMhHhHe8fcnc0jySfkKbT/kDLXDe81w
HVPotYr8iX4i7PlsTaHBm4DkWbLF6U8/p6L/a+FefaIXaiVVoJF+EyAUJLmnZh8u
z1pnG8/YZrwQkvs7jv0Erbp3gRhmczCY8gTprEBv3RVMnzRP1wXyeF/P17UaSkeD
fwASeQzQDHWMVCf7Cxnpi8yE7852BE6FZhYODIHg5hchG79xtWi2iD4Al2g4Szdr
u+vVpwdpMftLCjjXVMGhSy/rGEw8OZj+5x4Mv3QpKP+i0HucUAg6f2c5aYdStMzQ
1/Bbg/IoQc2NuRMxOQ/iXrzVfdLS8Ccc4ZH+4ANoMSlJVdvENQhvNEEVdnbWVbnI
fPgBl2QbIeA6q5tDdFayenBNEoWvMre0ne0gkrnFvzT5S3faMp+NSXj0RAR3tf9U
rK1j4urxtxoycPGwR6Z8vfOgnosHah0TEAucTNuznvwSvrdoV97mswGFbELhuXIF
4I5quuZ1mOrZ593gf+rhFUzmX/z9+i+T6bEu8c3pvjcZFrGlyYBGap4yUfrUW2Rx
XXDQfm9ADXcjpykqG6D85YFIyQta4s62ufU5Lxy4C+n7xYpAzMLIQokyboDs1v6S
o9FmhmYKOooriOedQ50SvbJxf8aR+IdBO4PQot4fgOXOrOzwEz2owtY9YKyhcGm9
GPtXWv8YwqIpHl34LtH7VM9WDMsrypnlyS0IITuzcR/AoZUg3V1crt+izTSoF1pf
OhN4qJjq4c2b27B/Bpc2Q6vru4wWaod2Ax4d+TV2i5+KLkIyUa9iwqSITJRikrd1
a+GH3cg3tkov5w/s1YXDvIbPaGa7Fvis7iet8OaJAL9jXDWhd3BjIy5ZL2aklL/q
nlCMOct3RCKafn1Tla/8LG0ZlTtJ9KRRZf9zrCAcAhVW+wKCENdErVu5a80P46Fc
u4jsbJTdKHSMP6c6ygRBnl3NCloZ2vZ4io7M2XoyEEvilF3YEBJAazFtZ/opya8y
dHSvUY0rraUPGEFotMfeJ989yJVVwRMf8zp+Q9UwW/z6Ei05YvBbGvw0fzzPjz9k
5anLas5YLn+c7sj2oScPcd3KLCa7nmdQd31na03cb66nIFUg/aDdtsc6rJ3YLMkJ
7VlxXac7Z4HgVF7nQpnzNz4jlnWYuH/bIDNthTSoR0hGDF4BSVvCi/8EuELcjV0h
E8gnQzgkOyWMBCwnc26T7Wc4UMXE0MpnqNbDsbQLjvF0EmKm1hputjYOgxjjonuL
FYRgjgJjYWa4g70tZ1+T7DQaeTwXswXRH025hGiSAzXwrgLRdLORHaJP3ZCNhYhe
Js/eJ+C9jYBgvmPIUYP/6oRvRGUJ6SfvLwoSP5LkeIg7C+ASirqM1DSG3fuhG5Xp
m+21MBMTpJ/YvbG2aiKN3onZsHh5nwXrQjnUCrwCJDjqwofQcvjHUcR45Q9tjJ+F
yDTq3qWAo+HBZZ/tSRc8hCDGCYArqijldMDqwTZ06sxQgdJJz5yngN1t/a17lhw0
Tt7Z/iYWNEfbMrUfIKqlN1HAs5RxZ4ivnLLXhRG5X18bOMxAqwdas/DJxKhjjOfn
lqnmrk1unrselGrlSvprUbdhbnKxRLKWrB+zp7v7tv8iNl6e8+uJe9m9U4ewfG2+
tHkWjQaRmewQV6Lroy0Yet6EpQ8MMXdgCvwV5AadyZY2VbszCOkx2ZzDuaE69CTf
IJswAZEk6+criczsh5f/i3gJUtA4S4rDnv8ehvpPv3JmuUQFEUTbliRBu/etLT88
00Udc6Cr7HHvz9I5vNOraT1ZznHZUHaNNaAUL0MHyJH3xD5YrWv7kRbAnN6NHX/H
EOOU9GrTjAP9NIZuaqJAyaqSqHlIjlxgeKTzjQnM5m6YwseDo5QGPleoRxaBOyse
Z5NKwoSbL18slF/WwvH2wHX+UE/7FQ2Qe7IAs/yBCNwnw2SbICUjdSc9lJjXX1LM
cI5eYoxCpbApTIuO2ufZgMQ1CLJtA2zzh4IFlQZUQPYvkk7VmM1pyZmDv/EphuAo
jfwio6dRAYRZMYqk6UbjxoZqRpG/uXdJaN2dIiT90p3T/90FRqdM4aNJr43cCoDZ
32ZWkg6XF7GXqMPx6xHcR9ywEMwPxg6nAHEM9M6JPmBm7dIP5t9rkxwlQ7o06zCa
IA3d72o2KFVop32Qjf5LG1L3H6Vx5rXnYLXxUOO1f1FqIeSAy13YHxJy43d/KHb5
ipA8ck9uCGk8KQGXSmyHJ+MHOTPpSSjHBSFqKM+vP5PzPW05qFoQ41O4sJJd8j/P
wOSzlyeKeiGrrqtFUN7X1UU3LuxPAluKlKAdEQMtt97V6SBiRYKk0Wj7WbwfpQNF
6znw/buL7MYF8reJt7e5dozKHhPCWrYE8vFaU/kJ/SnQCkmHnXihUQc5NIvxhZyN
r0i9QYbsi/TJrnfQGLr526j9/vGysQ4zJcC5wFtMQxbNcuBwZzWvmY04u1XT5Uz5
7v8VfNGNFxFsesGcJTN3B72j/ffTb/5ynEctgw793BeqwRkTtzWjReQseqpehVfh
0k1+7PajboLNeq9ofDvxV/Rd3F6ufgqK9eBC8Q1Y18W8obJjl77f9Jz5pciZ0yJ3
kXFoi4GXSXSYzAHj2znp8pofZ/xmqQaE752nAgdvdsTFvPRaJvEzBNj3cygOp6yq
hxwOMn3ehs8erU70n8zRglio5zNy7aYFWU6cz+84qrEQloUgBAyeVXro7PdpF6P6
KkNCbHGzYDJ4TT6q+CX1xsbRxYq9OHGGuErpEuPCLdx5MZEFVpwrnBFCkq7qRWfS
GrKfmdB2bEWvkpCyY5Ao4FG1Igmmo/tsQSIuYpS5376UPJsDPDB3Oeojj3/QuOpT
y6ygFPTwfsaSZKAbJ+UDocmDKxiHo0Y72nXhRNl6juxsg1JYwgIVNyxt1ZqA4eCu
UUW7e5IsEH8GZqfttEkLJZctFCV9RiuBu0EjgKK21pHT8JUbDwEV7zUNEJGCH4vP
GbKNC6K1YRyKY5R76jBAXrG0/9u9Z8a8uwRx5zeMXicqKCCsjvzACltcKJANi4pW
8CtqdyGDsf9oZPU5RfALtF1ZQ00iaFdM/XxD8U7tGzWI5LvfVOxbghAY2vGEuIcK
l8hN8yaJ1JnbcOUwzcKJwm/UK3HPI2A775Q0/FeJhBOQ1NI6iGP+F2xGgiVC8hvA
YiZ633zncHMe1AQL0Qx92dIoclIVme9VMN4XvZYecyA9sy7jlqISYhgqhpSna4M0
BWl2VdgqgqLSO3P4o0V0/7foBBk7ML1rMxzyiBLZ13VuhOJ+67wjAFVs/P6QvZEY
Nmd21spajd8u2r0uzku9ZkzAv0LJ6m00Hl4foTqMeerYoPQ1ZG9HYNqXRNVH3vWt
288141mwSAOF0ektTiIgFbNKXA5FO4BawtrMLExhjFqbtPEYiMxJKTCXraQDGL58
nL8QTDd3RCPS7Og3kWSKurFqiek+2NQRQ0cIfvVdng21Z1FOtAnVaUQfiWwFQVZ2
Rwkl5hfHL7cOdhvV7fL50WkHNp3uY34kVNfo2nNBqCFw8+OX7pA/0rLgb3GyW9Fe
/65abIhHqVmz1I2WfXfF60N/fmmSXba2NCjs9IYevJtr7q3v9dG+L0GE2QAhzQaz
EBaQZIA+foz2i/VkL88oXOmC3CXJgbWZmwmo55jMw0vX4l0c7KV94V2XQARu74Dj
HvqMPO1fPqgTEBXMRplBlS7mgCCSObmosnPCwu7Q3g/fusYD8w3WHRc1lyPtdCZU
t0VMRUVAlYerRE5cZMtWukuMbjTW1JD2HCiIl2lgdrmqvq00nTSqJ2Y+EIxiiSaD
KG4CxOJHoiKNFlrQdJnnFXO8UO8n2qx8CasrpAyRXVKSsXmhvg4UYDxOSmXuQlNE
L8n6yESAXhZVDR8pUUXRdDUEV53oFOe5ZaYiJLHQI9nJMvXc3Uuaml/5yLOf0DXL
pmvz4ctxsFJUPDzXgoezNueYeLO0N/8/3Yxcu27/j7X8O9k8CfOfOAX+s5jmzmkB
HW9VYMT18l+q2mTUW4PyQ7YI8pAFq3CAn+rvU6eQXW9vhZK27KhAeqpeT7JQWaOF
Aj4ltvFbjpQp0UcF67q3IUgFYc+/aO7jNctqMaY8KlF7k97k9HhGvzwktqQ7ntLT
i2xfjlYyfDER9YfGlIuMNgrk3+PJEDFiuiKTtOqdT8WW6W9btwdg35AfEaTngzxA
kSex5mteJpE7uvLCCR/GN+ja3lHcgeEWrLDaHajdfr7R7GChL3XomgRVgfWJLmIH
CbpM8UiOOs+rPseycjLxPZ6pSQe0BbNGxv22Dh6iWvmkHrzf0vxU1FfPCrXMKgU5
Imy7WUSG6e1rljSmqamkULpTv3iHp6vp8osp74lW9TuI7ITgqqD2OWBvq25vXURC
Ybc9jrkr6MFcUR6YEEksC3+H/cK7yI5sOdWGl2X6ZHMfxezHuPM2OExDJsD42J/w
ESJrGz6vJcrXRjA/UU+NlR4vlC/IGNS8c7hmBlAHkWWot5JOA662mNrXEO4FMxRn
pHVdWdCSr99RQ4SH3L3/oPTManhK+XVBlXEt3jdAWnOBnfPtrsG/pciO8uMwI++1
51Khk0hgzDezisTQXTkcoNqAMQJrfCEM3rOww0KmWlayGnywNuJ50vao1g5wH+QL
7WzN4VPeICxKTAlwcsbZHPbCk+6MtbsOzRMtZ+qrJMoR1kdXztW1Lio35cKMVYQY
QdDvlLdjLZHUfweZONelSAJRkrNnb62ax9bY47DjolRAgZRMq2cG+JTlBuqkYbNL
KILYl76gUtpSWagaSP7hJwwVuboaNzOBE3fiC0+8NqIM3CsHgIfrD8o/3lqBUAsq
vyNNyKF83UOJe0QHF1/BVaEmFhklRbjCNKyQxnn5ID5VNoYynuGWdOxOi31AQm3h
OzRJ1bma9TdxvVyTZ7T7Tun5x8GpM/dt1Msrq+zZo4YdoLnmo603Zw8ISgqJoenK
JI+zpVtdLWvpjAMW6wPMSU/ifmwXGLu38h1P94O6Nqc/52KjoZ9kzB9JyEPu7egJ
YM+jbsmTYJyN2k1IVpBttIQhHTojw8kPijnIXuSVLG9vc/unqvMJH/AwQuTALdOG
5grXeMv58XDCY71k8y5Ei0rg/bOxDNFPVNK1cbyVThM46l+AgP0d8X9psmeh7IqF
I7hO3Z3uO5BybAO7DQsW7VE1GQ+sVvkY4AzubkLCwlwJqg3btfaY4OGiU4PRzxSw
+AkWoukHHIsjHkDLmK/vmlih6MKs2spM4ZQCq24TQds9JCrh7DdoJqRGcodzRsXc
1+60Hbo2PNEMko0dVldroov0Jd4xw9QzPZottWfSzshjhxW/TrU5otPb6akvIJFK
OHWGmFNGavAWAAZNPoTs5CyDf7BRd3OZ+CIp+wQ+cpd19pBUBRO9WFVHIZ6FJdgq
jvECpIkFjNu6Wsf+KdrHZ0EGXdJ/XxczUpO14e2vFtXNIYred56KzCAKrJPe3cFd
g/zwMlLernkVErpGia1tzmfRmAYXYsyCnBGoP7Xuq8dxDYnFlo7OpVrCgzGw9fdy
+0mhqvyL1OuhEWAVoBuoMBSNTgV2UdCACbIDC3HwrxygFYU81XLW3dclorPWvx/b
osTLCeQTszWtRQf5Eke98M51yG5hWfVVIKdnpUMFimLcAt31YUQlb44FdRSoKUgY
5nw+RYq6olDQyOV50IKvsV7OBioyMCRp8oY5saCb0z8pmVoyJgLBTo0bGWFBVT5d
pybzAANGNwN337mqgjKp2uqAnGQGwv4UHiwAaDIF5jIKtx32zWwZT1YioD8U7b/B
2jT6v68aYp6ah30k/tdzVL4VtClFvVl7bGPWI7P3XJ2VnRqBt878ybcHuwJJcJLm
vLo2EnaVJmRFM09J23Wj1mS9E4Htn1eieWiSx9at2CNk0SE6bWEAwZ4LzP6+LzRR
UsTW09PGKSGbO6qvbASLt6jviCT6UieOT/Y8m7O5jObKUdcxGqe4aF3p/DqgRRBV
taLL5ifil3TYkKTvOvphegCh+DF2fjMGKNF7lmozN6Cy1/AUki03Qp3Camn5J2mD
e4kAM/hEvxUwcS8ud43g2wpsPBNuAo51LGxR2MVMzpHrOEBEsXIqegz4TbcMM9CO
HCJAARNd86LM+zO42n1hYhZ1dmc+2+R8Oo4UTEgbBiogmQeshLkksKPXSClRG/Lc
EG7Qm+Wi4f3Tgwly0zoQYL57MS3N57QEV/nwKfdVeoyAceKJueFgun9pKd4W9xPf
Ho8LnBJB9SU3Q0XA2ROL47GVxxg75BvVlBOPfwWyGum7fvT3n0n1qGv01dMOVQU9
qntcE3Tn76W6S8fjPFyL3obJbq4iy4qMNrF2F4qjdpxuTWS8ZdD2AtXvi5T/V51J
Kw2TJOXQp4wvp6ch66V1ZgALSIosliMDQvYa+x5L9WB5K3+EGXmh6Q43TTW/B/Rb
5FqbA00ENjH2K7Az4oe1bBRBv+/RWtGjeBVJZzYezP1ZT3kHb+9/QsK3E3g9SaOy
1zyT2YjWIWh2MlOVE5mNGi5R7CQlZ6tLNxEWRE9w7ib5JdtyDxbyypiFYP49VITt
IPbqujfJjM0KIKl+A/UWG7y/6fMooDMWRqhy+Nt7KhJpwZfC7Em0Z/r4TboAFU9V
PsVLnCO5/ky6UR6vXQWFfXK6sdpt78dOy8kGEndSjKD0uNhUvwTvjOLCRGjHD82Q
qqg8ztJjgAOBX8DPU+sW0JsejrkJQrfXjkTuGzcj8uvtG3lSzAGfdXRq6mjZnwXe
VbzciOwwSxnMe64ItZZLko8yVQuILbRCHRHwTmhjhfDxJXPGUuSCmF1AGvnEvxnH
ZBGv6YjKFvEIgZkLCyZeC6znrJXrk3xMCXIHPHlQflOvAA30vxyiGpnoJ3EPPPmJ
ztmxj0KEBMjLyiuEzZe0NJ95qv49JlJkvPXIW06qa04ng4z5VSfuXLNATu9pnX+m
fdA7YtBnB1A4Bo7mwmGZ9wl3C2zi5Me3Heo3e3qGOFcz70g4aCBuccJQRll82jf7
T/46jVHssxfEJsWy8NffcxovC5T9y7N7N1P14Hix/e7ugqM2d4O79C7v+vAMKY/O
SSiwZKcZKwk4RJP8tk2Xka0/80G/Mi9oxwml9KgAf/VJOJuelKz/wKMG3cV3bFpK
VpXM1YGg7e1YQ41SUSU+TI63xyPG1777zC9F2NdZhpEDclFbRxCpGU01iy9f9WWm
Pfk6G8Imlz8juYjIAK1ncvixzY+/uVFZXWBAqTh2VmdmZrxhDaWR1QUNmX6s36M9
gZtklKeGlDgC8YgFcUaOClB9//Zv6euksTEGVQ+tRbtkduGvxfCgB08LUpQjmI0r
iRrHtSIxq2wLx4/eey+1jWeiWvKTGJZgzLSuabVyLkP0rHVO6FRDXkD6YXGIlUTw
M8L5rL/4JPFslH67r7T6B2muUb1/O8zt7Hq1CfyKi/q2uzxaI4RmZrPocpC+HP4I
hXlFskGdUxLcvA+MVAkPmKaLruMI3Fp752MRsJ4SdAzRAu4VYequS+855dSgm42n
NX3jZpVrEFOJMtaUJG17OWPQIYH5xJUA4EjsHQcBf+1955AX3FHl5cqEBB5vUFou
1rXpKIDqYb1x1oZSmig69hkqP8lcaOH0en9cKp+HP6d6+8u5zu9v+nvK5sTojvCI
iKcdWg6Ik8WHnsTNWsmJiSjtBBnH4tamI/WX1y3+/tLDVuLBwFneigrMXvbwkU8p
v7wtnIpeQfRelACuv59SjhSOJWdu6HKkUg5rsZYGM0CvjQBrEknyKBNdJFD7BIoi
eznyQpOUml5k0uP9eVUznRBDva7Cpd0fTDt5Ar3ES9JRT0j0AtNDyHxF9xUVgXgQ
wYsVxwiudfqBCVcNo+ZUHyosgVAb0p2Q7QcpHIYOBtqx3O7I2aqw/UExGfjBlkrm
K4jvHif+je1EvielLmzRMvHjOHLxTGG0ViU3Gp6IWYSjHbNSOhDRezpSCSxhA/qm
4uK70hJS4rTs4mC10Nv1dOa4oDGZ4ZUg2x4WCx52et5TGM3IRuHSGpq2P9lCauP2
wAmJIxIsZ3exTCya7uroY3mB8uQjEz1mQgSQQknxQz5kFaZrlOXz0We5SeSgCZS9
/V9en5Qm4u1iEhiwkFiSoAWoC1GpM/6CcDupwAWaa2LWKjJjnMv1ZQLyL9OYACV3
SjVzfL8EQ2rVZb7HhjcBAWUB6/3CFbVO6QGtugXLGI7LjP5fTqlGz5vpkAp2Is93
kT+dDShKpwTIQL53SkvQblgluPBEwSJ9QmMYNkocPWvlgNDJ5JI1LKvqVpmA66H4
wA/hx3rFSxM6OI+p2LK9MKj6w6mmjRm4RI4p1yCcKih4CmvFe0N1eBoYIgfOlBHO
4K7dEUIryfPiV5bmZBnWQzdK4eLHF3ohkWAeyeC2xkmQFyV6h1Pt6qsqezmXjvbT
KSu8EXm7di1SJwZguSp6IQakzyl81owccUvOLf+xrkP+G6B5RIa6mHTLO5/G0Vk6
Li0ucre7YPdD6PiNnZtdkwgCs+mxp49qCSAjQ60s/ebxLU6D4+vtZA3FTK9hkA4D
uCPy11/kiPXIxZeU5/v0YN+U0JzzIoUh0+rwBbRs03MM0EjUdNmmBPEYPMXCVzxK
Kmcq6C/q+StBqcifbdKpG/TPeAyvWumL7jvn8AsA6BlgsH+XCBuJKBTqjjcXv1LR
sPXd5AVUFto8kMjU+/zl2sN1+0nE9uQeeESBu06AHbGzdBZ5TLFefW8XiJsYMe6Q
K9v1ZGj3KKORYxgsPv55KnUhGzwuXVnpxXP248iZWndJgR8nG8Pxy3rrUHwbOgQE
RvV+wTuzyQoB96putgJf2AdU8XZxrrFTDhENzvhjlTHvB26lrhd8c+Hdl/y9do4o
Q7zJM7VNBJVYdYKCyxpdgsiDEnGotvMMkFp0My2eQnguJnhQ4KyuhYN95cLzqYx1
/zXw9ERpNiAFKPnrzA01bdnuSpMPO5ssUPjTM9hAO60Kl+DyO3ztKG70P6TRTQg9
zLQwQcfh0fZcMUd7iOqEN1OKNgTr0ZMipzcbG8xMdT2uQ79HJSzM51ajKqpj/F/H
lDAgELz6RBHhhGJF4hpmY2QemFjbCMo8R2tGE9F52uicoors78vfOtU/WK07Cp6B
Cm40YEM6ZxcsRKoCLsJWZeVL+aonZ/9Mmqz9jrbmPF/L/O+LgMOpvyFlguehSJl7
v9r2jW94sIRgl7dF3VQozi1VPvAfSSt0SWgJBIyQ59QgMZYTKDDCfEibDWVJJwho
e08xr2FAjOrejnZv6DAB5gncpeeH0jG7DVAALYnietk1x1GuJ8vTTZheCI+p5gzD
EJ7zBW+6YfqkCNkNwRXYWZsoAvCyK1FhQU9sx98ATj4gKRsoGcaEaV66u+40KziP
8zNH30ur/zQmWw9/Ia5EODzUZhaAcMFrU67xsNxi7cs5A4WI/hk9QV2ikcTs9r0g
8qlykDbv6jeEAreIIWyxbkRnWPAZtHfJwZdlAGrv2tdrXbjrq4bAkqi54HqFTqQ4
TA7wlY95t3uvfhsxDr0vfptQyejHbxFmIMxW4jKPqnwo/WhrN52j0Jgk473v43NR
iVu2zRUEpnw7DXFB4ytf5hGeXHn+XZF6MhOOa5p97vRBSrGrJmBnTt3IqY2f48Bw
s7+rIk7vR8otdI38+Q7GTV2O+XPlRkvUCLc1+U72FfPpIPqJz3d0S70ITerA4lTa
46r2Vsx9jlRtwIUYRHkk34hZ+LzaJ48CCIj6gu9Xtb+Ek9MbUMPOk9oqmPZTZt4W
6Ok0uTkZRCoK8j6gl0i0sF7DpoFzz2q17+lopF+UAVlADyv8fcAQUb4HCdd0Ftty
SnlTt38vpZcSsq3za4Cg2zgJ69aJ+WdKqbBNYZdWRXP6k5RB8Vkh5KGmtW5vgQe9
lPR1AsGn0hikmSdO+I5Qy0NM5z7WY1akeU9l0FBwslLDoZJqBDOi+EJQs3p78895
pA6xCVtMPGKnaWh+MHyyQbE/xgerKm3QMselogo9yX6RndJtqsCZZ8ImXsWmw9hH
+LLSJrHLPSk5DHaIjhHIXAOWpXI2viUCO/+rsNqTgqTOGVKPrGCERl2wxClaOwvr
RYUJsWXzG8dAL3bf8Am2dzxqa9QP4Ey7K+cgEd9nAACUfVbfjaPdo7k7X6XR9PKA
3/NRJnnVZMUZ89w6hwgDSmghHaC+GzF9xc7jghbwRQldQQYt/qCtqJVq1Ou3WHlb
ntQrs5vARN5zH74foM7TXzphgVHJIJFO6crfwZ9Dgqfu+9oqMYzH8kGhqlBittfj
GuEZ7STNfCXLX3ISm0eF1MELMZgjtpHEEJBYp+ATrqekL4VQ4XVgbtxU1aFnlwV7
HkAbKmR33lzbWc+TAJviuUfteGuQHwp4QTEr8TbMBUfrHFNVKQqYCZTzt9rCu8ds
kk/JlMzz8rLndIFNTUgVrE7CLJyqO/FaUSE2fPtN31j5f4o/qB2B3/HvDfBc2iRM
KU3RLFLPp7R+5v+NCGMU3NW7KjTvejUDlPiHzvEAiAld+Z1tMEGrkcVsP2nGF8GW
TW5Rr7DxljNXaLUc20eyrl2UmSz0cCgKqmBNn/U1iSeQ2b+YeNzYjqW13wOcnMsG
dn9ljxHrcQ/j531rRD2jtrZHZdNd3pauMrlFtT5lB4LQxXrUOyiDf51qx1KAMA67
G5RjlNajojEH+tnWJu7nwModZi4IedHe2SNk76QeszD9AL51WyUBIbgiHGk17iav
0AGUuvWIr7k5ObZPwcHe9mxeHRt957BatU+s2PtgcQcqG4pzOcCvaWk8VBTkVEOl
ILMEdjyIIN+ORMXk3SP73Cb7N8wgl0kS9WGQbFhPxkxAU81ZWOI2O1eplOUObYxP
a9d1Ip5WdE8AOJtJfjZRKDLCUAhV7i0gX+TwAVl0K8VFCQuoxbOoAMYZonNO/XrM
nYGaLz04sSAxOw/HvjnmKeygyrdNNBRhvrRc0os4GTYI0ggawAWmcCTLE2JfVgeE
VOO3jWgq+on9Hfrc7u8RHkT476rX33+YokE0yT+SRSpnIq9XE/UIdCg80t2hCNEY
wO2o05gFQbvNyAxW0B0lAZhEM8y9YH0Xf2jfp5dbkny3fmp2x13l+h6oK33lTvDy
lGw9guwIxeAkIjQN8Wjdh9cReqeQfspSg4z3LMo7gLlDHCI9ePUR3RGozxeNeNsR
FJI6qbX7Q7Nn6QVFV8ryMzPZtQhaiHQGaX7VA8s3HatmoNYKIn9pEhSUW0Cf2P24
XYHHAVWaK4R6uD/3jogzvxz11BRdkv5QrrHalFCnYOnB+P2VZoLOYNOBkBLsYcY7
6HnjkMdVJ18S+4Cj5QBTbLAtPTxMjngX6VRh4N1KtqABDMgtY27xsrvI7DaahvQd
IzV5ywHr785n0ra5o9FihiOzapQHZ1zcSVGPn2z1TCyAFs0YAIPfWrUCOCd21m0W
Lr2oNTG2SVFHvZJ1VVRase0SkzznEGqZM7EEhoJTdEQXbCbJyK3tfxHRRbxaDc4D
IZWwkFJ8sthaFEn0D298EPeUdKr1ejBVpRXl61Mq+C8K8egp8pFUBVshwei82SuS
4LM8cPfpC1sd1ZUGzk7vtIEQ3x67Q9GS+HB8DRbYQpH6lNmg0/Ptq9/LcWKd7szH
WXbPd3epzf0nBflbxzefRb74Ld4nM8uuQiYg9FB9/Nl8A0DRn3wtgvMOUcyv4wGJ
d8zr6illRmFbjsYfp3Gik8faCeRxNKvalITimC1hkBKNjIsIrj8P5vnufPB7vvxL
mWWxyLMV5ohhuD6xhH5l5aLMthXIzaaiTIEFiwsgqF0/G5+JqBZ0Lbg1r4h8NNUd
LNgb7cgGSzg3dDllhUGDKAxhMI+MpqWwlzmZraTlJkc6riS2RFttameOYS/NmVFn
JBHCsU6HEdHp4y4rtvJf3lUE3B3YsLEKEMjfDHhPsaWerPUwTEMDXdxV7WGHGU/W
pl6iXHhkEbq8eIi+UJ/VpiDuA12murPrFC9/JuN48knKCcQfCyJ8OQei+prdXrpp
0f1rhq3o3VyC6v1ulqMx/+R0Gm4Wik/hCL1AMDuXdirMfZtWTSi3aEXy+0XdXj0V
weQxhcvFEIFj0JON0/WpDQj8rf3WocjUHi8oGBKUBBglcFux4c1Y9cUWmjcoq9zA
CessCZWzSu/N1SfZkjmiZYZP+BV9/99HMPVU8XeL1x7QlgW4ccrELxbaOrH44ay/
ib5LR00czGQ62HHQvVs4xw+wMiF2VBJ5Nsal7cm+gfhB8QfwefejXr+IW09Qo6Xa
LAaYX65K7UHibG+n0AAmjuNWVPIb2lrcppdZoDsapZc1tt4pcwKZ/dJ0Fz28vv95
ZZmg7jKkujVVa77P8SqqAOZHcec6Q9MY2NOinjEGn9jeHT6/2Sm+IAw38VYjVy5s
aAD1a7RGZoTHAN0ph/4eBPJakZec0RM0BqOYo0793XuBDtK2KTK4U5Wswo6ozV2H
awL85CJO17a8fktlYN7YAoE6PAI8VCRsZzuTSMpda7u2VNQK7FWwwfiqvzD/xJL+
eOiO2RmzzgZ6Tw91D5GgVFYcksjgw6uufW8Vr2EBrPAJNfc2W5mV+T1ulagvfMbL
hxZi0RIpKjhAj11yIZFKolUOVvoqaU9Ejp0crDhwK8SwMBdBJcA0XgN3m9ftJKXT
Xx7XdelSbRrMebS/z6LbI8ZOjvvmg1qOLkDTf3AQEq84aE60j8bfIc1tZRpQsQ+i
nhGIGDT4vO3ucsXCxBlIdXNm7nmroxwZIgyyGopPXkFMqH3OW1d3f8T6Iwp50I1n
Keflnv7YEVDz+He+YetAXDKjpERlQsuIahV8gjHsXZNL7+efWcoWD/PPRmbUcDDX
kmFCcxcW88A/w5NISuZOQBoc/OOyUQ2seEkAkzPseTSYxYDt/VvtbT2sOVRwrn3p
rXSRGMG4englcvI2j8T4MDdqxT/H1iIQG90Fxvcmo7+m2EYgwOhzd5L+avoyDv/n
QjvHYbiWboaibwFg2O4oZLoYBMwrR97eRHew8X4xY3384jR7cQYKEDIKrO9NnYlT
od8bsjoIwV5aHPLh/3Nuz6/erbTmXZr1hEJhzl9EdWpDMryku9vOU7dwDdSa8Kd+
SNcyHeqXeGXbbZ5LYfkFrb0WTI/SHhYtHQNGlN9mt4B/qRSzmabNeR8couV3NA9h
ZY73BkNzqfqijO1pjniaAKuhF7XhUl+Js/zbxMFu4p5CWf5bV47dR9VXbBiAxkje
AcnDwNkF2Gzh3kBI7jZI1FsOeJhrMoztXBRHviqLwIBKb2neq07VPMkoZbzLI+0D
JTKMx4Z9+bGNKE170/5H7uzhHW9ZD9/zHf68sBy75PsIbgz7meUpY+zZbuVY49IF
/S9Yy7Y0ntsONXL7dMZLEy9sRt95nwCXZ5X5d6HKP6uQ5C+/lfT78/kX7Eck+gnE
aDX2We069ttWYxT4tS/UbvvYnaoCDdS4Crzbk4GCFrBSI22zfhttLmy3GXp3FAx4
Th5jgzGfrocyyQsAvDIVF5FYW32568PdLgN3VgoV1nkY7sJiqPoLqxljlkaPUBHb
RACevv4oJT2bLVw8nf7Iaz4eb/u7lU7kjEjWbG9x0z8gGPaFDXxPCeSSxUSIAMEF
3Fy8VB7gTsTyy19fM/URvVCj3bTkUPObT9xKnZb5auGxo10/9pcAmT/3vzlW8M2l
zpYWRbi4vJ/C4AwBGVFiaxVmbUcdNMlyIf2iIojlI/BupOi93tQCgBVEfAx90u1n
yzhl/KryPtKsUTlEDc+QMxnfoIQ6DFOVjgv/fABdka1/p9FAEpj+QwkkN5CLup8o
ZvwjdyEfxYqyugvjXHkQAv0tbllioBnVXP5tY8S1DWpOXeYrkaC4p0mpGSMbOFFK
8csG2jnD0UkGMPorI8/pNg1Mj3IPa1P21tlaLG7zBfx7cukdnZW2TVYdcODMmZuU
wsdiCc6VJGM+jYSGTlnh5D2bsJGynTNA4M57AZUJewDeQa04rdN0Q4tRqkVoiXtS
Hb6HwQXasHx6erXMCQffNOOqqa/oATpt0JcAn/YL0yEvP+xR3Oa09iAM72At/DhC
5FZ0+ztP3FZRfk2tjCw2L4ec0KaX5A/aw5KO2PpU/3z0TeFrTScl3Q7/HzZ42Jo3
zzJunih8YoY+TJKiyJCH9B92BML3ccgdKPC6/7lteDUPyDwGSbdZM4MmnvdazP/D
g8eJ68FltRAKdEtX7ym5+/pd6FH2gJuIZIeixkEr6m46CaDEA8kryJJU0NBhM1Q+
KagxmFu9UTmFJvXjoDWK9SjgpGIbwOYuVfOsiCETehjLVP6Vx1s5VE67B2AIE1Y5
NbCb4c3d3bDy7VH4Z58/nM2lFWwjkYgSLjkfmk/4xgYTaoyWsaK5q2y4xDQYesnD
9A9l5oyxi5cx24LaeNkpzXem5xZrZMpYU2LMQTCjG4XeP7gQcLe9O+tK75LJm2tP
/3Cs3X00NxWHXzv1VfmigGhTh8J0uyLiSQszcHu+OLSIBJd0BoROjpfVMY6ry4gG
afrqlC+rEOqfo4fNMyicvdcfmOlV0hUkQQi9STzX8t+uUEMgtIXVJ8VbRTGxXAGq
s/R8CYHHubjiAykvEZM7Uyuuvtwv3muHVaoQk3Xyhaf09B31aZbGR1K4qypep1+b
CWNDx26+0RfR6GUMegZ5dBLY7uLRcObwUM3s725v/hq5XTpadmJ3DwYs5yanplAJ
B+8sRkfl4FBlOV0RBLtg4wxqB8qvnGtxUmbbsLDDjKg9+W8VAAGIE0Pv6rvx3jP4
DIMDD3Z90k3NCLNjJBA4TFrt1m9KJBmIz/LaXH59aFpKmrQ2qS1GpfhwdcLMO+BU
nFsepuEVPJlhcIo9c+QJ9MwRzThJ+3CVO8pEE2BNIMgSRgADZ2FpbLrbjFmxQT9g
+wALo6LTs/7rOgl2erI99SeF9TEXEWz9bw2iKFvDptbfp7qMJ3WGouivnda7LESD
15jfBxBBPFH8FDJSGWLFuODk94/gCmEuutHsMQHS1/p1pOatcUYrxxsLs/4bpHyM
LB3RxkiB9wS4i0wwW4IQebjYfPWhWpdJv5Y4vtnzdIPlK6QbtexpoRwbjXG5/Wm9
dcOwNmaGXyObnrBC0cYPXlFIrC4CCMlwUgDTd7/TicZKlFj0BehReo5wPLBxtQ2Y
OLntHwhvxxMDZS45EEPR8s+BRDs4hdIAsFSk4/p6kthFaKlLJjykxWcVdEOsfTbu
wo9Tx1doD9PB75rGY0O39MRx1Q6tdHQM5yZKmmqOYXxFanBeGujclh0y2snC9e31
1wgvm2MYzpDncT0UCX3lenTtshlWB5/m0KZK7RMqW+E0KFkSMicKfOM35sCQFG64
HqhRaHGHKdPCp9ocXv/33vvyMoiRvPr1/3tacXpSptAo4FBjxRevOrMWQM28Y75b
emEx03xrkyJkMzEom/l2vnDNtLe3CFi1f3Kp30TSACOi4p3BGID1eJidYV3dwdVB
LWPVrsyWpFngLUQQ6UXBDst1Av0zXv/ehLSyjjsULA136TTCyyeRaO7BW9Fb0S+0
iEGh6OpbdnLtOAOQGEv3g4o0gIZwTkwTDZZZx8ECKA0bZLpUelgR5lHLECgmAe+u
Kf1V12Rv/ZEoLfgzmvk/xlXv6k3Dn5zuZyneYBNPGOWXuMQ7DqVj5Nuvr/pGb2fk
0xzKe2lHmuNlkXWyyJeg6F7KuyNrXoVRHeuceHWV8DX/Rq3La7B9yDS3P2qt5+yW
0j9UwH1GWdE0ouTVtJZkA4sKuUenlU0A9ysxq3peDVrW3e5aJeeomFOP7nG/0fRD
XFRXXHQ9BIxxL5W4NijGwWAb7iOe9atFs+zU1IB9pP9zhQKHcqj5nSw1y3EpEhXJ
R8J7KHZVVo4XqzZsHVhNERtY1MPZjd1Yz6X5sBNLcQTcop3BU77PPgIH79Qio37+
l5Y2//7p2nNk2JNLJGgpkxDNcq+ivUbqrVl/swzm/7H2ut+EtAN66CnN/chwthPW
/QN197t4BPI2+UGXZ94lySCnsenIShr77+X02MSI0UaM6TPpKZz0B831yuoWZVql
vwBzd+wrTL9UMBPsM5ukga2rclDWxmx1N3bNg9LyS43f/ut4CDmFmbXvgisWgLHF
/YbDIf1vP2leSxNh1WfAb54+zJfRzQ8yNT5QjgvmO39FY/TwXm5QZoCocz3mpwDw
KeFK2JHBSWRQsz3yq7YLYFBHs/4S7SWHPIhgBd1X2558smnRY/OaZVREJP5P8VCj
tYveTKHfgL5pOfXXVcQT2PgWtB0Us230JyB8KCP8iB4D5UWbsomt7pkjN+2TumqI
18RwUQdx48/yFH47OTYGGBddxPrQFhPHW0tJVVxKWFWgM5768zgfvVZBwabhk1OT
2WU+iKdY7uMuMyBAYzujg9L+xnAm0ls/WmGCKIB54lsP8/8EXb14vBSa4Hi4e+AO
/GjTmgQaYno8V/xLdJvaxekHc55udfPwiKBQboCjVQG127SUoimr4kI9NJWfbk/M
ysgloYMTImykvEPIN0ovuBm/N82heDhlJJ2reF90Ykhg/2pR3+v3SDqmnWAG2Z3W
hJ5SZjFPx+BRr+h7Xi6BhbDDdUQtM+iaIwc0ZfP2RbLOFrJIym5HbTGr0aR1F4Cq
ou01hSpKPBJxZXqQIaR0jsEANkm0AOdZ98V2dMH802+DT1D3XuaEbl3Eax6d404X
b/MmbyyKuYqKCGGiwnYr3zA8zfmcRRw1ZQAagoBZA8kIwKUmhVnFvltfi/k3qn8p
+/lqrJQ4e3VgL5H8z3PRIUpAzMloxlyQ8mipwvmehhU0Irqd2MRPAxP+6EyAvJAx
zGxuIWLgiTOQ2lzySoxuiq7GXiRnGxtYTPtVsnw4wSpkJ6Q0Df1QSznyVAjujbmV
FTtVpYKiyajvPSk2vqw3QvfoFOWQ8zSFCLGoX+XLN4SKUhuxlPwI+O+KsWLR2ICs
qEg5Q7ZWKPBCzgHYLTN9mEhDfZzy0M9ot8RXAtMH1RvR2rYptCjX6jzOdND+rkqW
iuV19eZMntDgIyOtbNiWKITfJl4cZcyhXM3L5mR3pGUA0Edz5QY4MVQKaoqokdp5
jPSk1NQeFXl+DBXTZkttM499bDXodIu9TalASmZfew2ndsFESPbOXX1PjaCxSbce
MVFB+sCgGxGMUciBoKUOGPoSKHM2+ewm5QZC50NUZHgO6GajS/lRsxWkAEJkfV/q
Ih/0vic5pt7vA5GxuzR1wg/EkM3MPHAnniXf+6csigBaNY3FBGAwRb40X4mUl9vd
VLVjYJ22m12K3ed+CccezQoHDu+a6Qn8jiZ+Kz8GLiz/F3ULTDqziI+IHN4QBRDZ
ileLsE0FkkBFWyaM4ESPtTy6ZHcOsP4T6wUqaJ+qLz+zvvO2S5XURurbXGzfMi1r
3SVA1rSCZvR0neyzJ+pgwLFe5IQaf296IM8BR/6ZL31FlyrthCdUdWD7r+DDRj3o
21elL507fUaNu2+0qon9CUL8Bk+w/1iKS6sJzHcnSPGCrorNmLalZX7Rp9HNmsDN
r9Mij3th+ux0dknPzX8N75QknyYIlBhAfnhEsqLcJqdCV+aid6NKppCGzI9lSbem
gUOx8Of1JCbWXzAPqqUPxcLYrTm8Jv7AksVzIhFbKCK20O6n4lAojJ2YZ6N/P5nw
FWvKhc9PCWCOYE4Pd3hnNxG/Csqt3/Qb0ZBg6NHJmjhsaUKUcqnG5D35n5WdmIUI
UhCRgX8d44bGNVEa5XIIJ3B8M7vw2aF7j5fKBY4mwofkL+gZ9R0yLZ+5Z74OrRPG
dDv4my5TEfNUu2O+arryPK86xQFqbrYOxe/fcyU5UJBNXiXW/dAANWDVxlH8QA01
93ZOUmu3qCU38Ng3Uj4ZcCsebcNy6EbZzCjKvFJ6TuwkF6se54BDC1RTRRRbkre+
nkd+ftIuWxS/3zU8gybXD4ABwfEgH9sNo5I7C2fa5vT1KS9OB+Pr8NH414TGF40/
+dD1eqmLwSQT25Bzy82q6c6WlxPkWeo4xsrn6PbDo01nYtxANyDFOXx+ft351xE4
8hXI8xP1e0Kn0RMzLulxjeckejgyO9Zk3d4yY7QDmlLNrL7qa1QdbD6oShwuwql5
SDjbz7tOYTbIrh4upAqnbqKDVJoNNH4q84jGEMCSs3OWhy0JHLvQVp0a5P69Eshn
dOMZSthB/VLh7VcKPk0BnzNW9Gew9AMeG1Uu8xguTrUCGZSDMbP9z6MqZMVZUTim
XYuhEvHVV5ud/ZlZdY/hoTmFQ7EEIQUZopmiYz/o5FAIToh3Y6JuJzwxBdgm8DDq
rvGCGusTr907jwAximtJ/uMK5cMM8/Kefx5vvCGFLpMKDCiBBgm70SHSBaWeUJ/Z
JAw6ELYBCBrAOEDnpi3bayY3IMZoWg62XUDfAsgUfuTHYi1ZJnfjTVkXMrpkQkdi
cTtsAExlo7sriSlLNfWKFseVqyNGeAvfZgENn54T6sGwkaWxJ8SGAZ9P076ZmwEk
uJwssdWLf9EnPTbgMkvY6u8iSaEC/9VQB+8n60u1ldoaS+1HLiSBh9Si1xbj5+SY
IBLCR0FDTld/H8p7zGTeFMa+7XBfJX8KNBl/OTcCd4y6ToIn17ovfe2BCy6vtgIy
K8pKTXo/QBq485hP3Kk6Fg+uH7WlykziXayBUjdGda/6FFTJv15raMQu9RiDCl4/
HlIOGz2Ue4lJ7bi44J1q4AsOeefZu11J+FEwvJmr5dyLnGfdZ4cDTWf3lYkxQI4X
dCceQHRZaKkMkKcrR+4wM/BvBkoO+giBTrUyZDWOwve59xp9mMKWJQwsdFjLJjaR
BNSQDzpm88G85dy0Nn2pkydMcZ2BQNLP2fYHHZtnFCbh4ZViQR/UvN41NdYgh54e
oHpUT9lTGEl84j6yB1dxqDhc9mBUvN+y/b1pdjluS8WcGmn1FvI7N4K2hvNi/B8V
C7Vf34RDrhoQlpEkBwLvmvuNAvrU3WgNa80XFF+deOSGIJbsjqSYmt6AhPgswqli
x517ZHtsxch8LFovPODD/8zK7feMMCL+JeupEergCcvRiMYY/MVFB0k5DjBb/gXY
t9+5rZd+1SooKfk/kZaVQIzNxfReWfR38F2f5IjC3d/gcuMfFEprX0xmfpENn9gY
tAW9RG+ihjKBf6/rJYKdwb0OGFAvVFU6SioiCoIoB3g1E4YSZpuYROyRLH6ozQPs
SK00qQIXtQYNckvcD8DalWic0OWBgrpxFQn4Nc/72pyurHAhNVGHtYSbAEjWws7r
Ja7hXfHsIJSCfhXpPwimDRDea8xyUOGtKdMWCMlJf4crkUeBs8wB4KuQvFImDiyf
VOVwh8iSYWVqKdpbMNAAPNsxYVRj1mEOLhEXmATJmD6dMSt1kMojBtoeVCie3p/a
1cTxTxpCFxj08Petfk5dvfjF2iC9wewizGFraXpGTyO/2r76dxYTLpBupCdk9lR8
Q4g+kJIxrr6Wa1tBzOYrVuC67Z3HzgW3OBORKV//wihGPuSCQD6nHMv8nxoclaKD
Hn28nrenyepLMnXXjfU0WhE9JfcfJUAv5XbsWdCn8gVuJ3BzCukyb4TSi5R8ksp/
h4iKBYegt23BrDC07vLv0gnAhhY+9UoM4fJT2o3M7DAy/OWxhC7o+lj4m9Tn17j3
mfOL0B1PAk4CXwxyDjkyUZh49RGNLZEiASWkfykkBXLfkCQR+NJYsDXqa0lxHxPe
HOKzenaWVTnWFSEU62vS2ybsS0ffWv54hSbdXV+9nPKsPUd+lw3q1c+puqt6bNoP
mWlpMDcw6X188iVg7VWWKRj1cpOfEfqY1x/gFuXsn4+BrQzbMUxmZoqRSTzN6bq2
YrlnRLKbdtBRRvYyDwKZb9uiXnBBRpRy+WW0Frjr0NEqQ7NK6Lh5EgErpDhVOLxW
UWumDYOOF+h8L/V4IaiMSg8usKXcL3goAjeHNJtQrJiGwB6G+mtgBG/9MM29lOOO
69J6oQGNANXeBuZE3lkbXW0bTaxjXeVgrGBfu1mXJG36mjcc4LeiueEHV1s6d1D2
FlzMEM0pdLFu1EJiDi7crkUKGRPOr1e9Ua8RsqQvULw3NbDihhYsF5Q/8k430EKX
poErbOzAzNLBs/xguCA9yd1YI7Xh4q6OHGxzlJdlfab3jd+sH68046Yz5/mBr3s0
pp9xQSRAygR4Yxmq1hyEuQQkdwyWLWsCbNQYnwNVCXoYh+DJlzOq53Kr4hyDDQTG
S/Tn8OdIjnX1kFxxq8/ExhjM9QZuCMng+Vx3G5TMfeCJUMedXlweVp/XprqAbamL
LMSdiTaXdJVVbHrd8XzUrQs1AuX8Sg9b3QakwmUNOBcDz8Mg7AYJ4QzidTKZz0R7
Rr9Wk2zh9OPT+lxb2xGPEshJR95UCpU3hby2Nd8BLgGMJI7WYCcy/DSn20/YcBlE
ztISZAKX72FAYBuLifeU2KznCqORQ/3EaUWnGzEqMrl6GB+/Io5XTzB4baRyG8cz
rsFAyyt/23RUruyw9YbUNc2atYRDv3uPnjpoNsAiSONrIHZM7D944y2JRubHm4BE
T/Yf2LX2xdbFVsCqiQ5JsAOObkVx1Ya3aTe83DhKq21WoZqFVtLIDvRLBmjnb/xB
If0BbWYpvrph31IP7d/v6OnZATcZSJ46jTyQZQHrMZjuZjlX75pnVuZpepjSPxWE
eFG/O0f1P0/8K+XjUdxK9dCj0juAT3TBxw6wIY7LTwn2Sho3e/CI1rpSL67ZGr57
H4qmJcL+F60kYTLHJL73IoBqmDr4z6pH8auV9GtXoI338V21HfysumK6jC3rpyFv
kVhImlwr2UWvhlajWLKg2j9bI3VFKjyqgTeAjPhrXX3Ev0XFUXECzAZ7axVb1wBG
nilgmN4SWSs6n6ZtkZ4qgHssfGBe7yE/nXE3aMbBq/GSm5Nq9KUwFTF1Ode1g+T1
msJzFtCRZ1JgGVotT2osJVk4l34U2GnY1mq6uodvDPidQX8tE9qPL4pkmCdtM3oh
NcMjxYT46DJJjneOBDBFsrDogUuVQR5XpwzA/FKyiREiQKL7Jq44QQfGO2XFWzSA
BSA8sQ4mgVeZxuXNayoNh3gxgH8iR8fqsrn2NMlncZaMWMs6w6eSworVLNOjtwbN
lZZ8IUcH09bAMDlWh2H3Pww5r0eFEisA8eH7wJTzccfQD7dv81w9QgAY7OdBjucw
ILCneLeWbPATUBW49bInZTvhyK/mGOUpEwFXvw0a5Zqb+CwTqgQ89ON+7YfnJt3C
eEBo7YTY5OM0rfSu/qlAQHpcakE08KB7xwZuMGPqQYRkl0JDMqrAFbMu/SH+NfsB
pKJQORT4/Sz1pWyMLgt34mhbwNhLKJSGHstyfx7intE6ERGx8yLpA75O2a05n29y
qRlhy0gHiLmvoeY44HjxRsN0zGdQ5ot1l0JTxbp+6eVsxd5ixZy3Mrmmw9KH5baf
knCqAZl96tz26air5wC/oeQvJ1lgwyDPEajSnfWZAaIXq7vIWr3ymtmwAMKdWHz8
z2aGKcIXVFAsijl08x/j5TAIQwW0ys7A8Il8oOu+lQ9twRme+VgXddv3DEHHsTXS
xo7hD2XMo2WxjI4rX8FOqZaVEDcofJhev0sMjUbpiH8qKQhVC2npjeFU/9+3o8Ua
6v6hYiq8WvISUT4hIvYMBXx8YoccBgYhXvs/xsP7yeSeCqpykAyLLSRxyGTxVEEj
LFlV1onfC+0nmHN47ZYzr84z0BWwjzKRRhRjIaMqw0QMC6VjLGE3cjSE1cbrVMJn
+loIo5eDVmN7G0qGdoavGXaxoSNoBjAZzK8Rxw7kWnVPY+29Uz9XgKkMP4gwpvwS
ne796Uf4Dp+d9SvKZdYcRaR1yy4xgNcnVSvWIvpUI/qdBZe3bv14+XLJfWDRaugG
eLOT9BGvR0RM99dAY6dayO+JRJOVwYAIeNyD4PQMweGz5g7h7JHonDy01dopspGr
vdvDzpmS9uobW9JezIwhT6R/T2lrk54sldTaeb8Hiw0OTEkiI63ZT1bXAimRidX8
ZEQCiN8zp0O5PVWY+RFF4DIYozseleAlin+LNehXsQMksXVRO5e7IDQqXXPYqRSx
7gLcFPPiCcIGDk9wQZUmzUaRR3SHd0LoY2waI4ePVMxIYgPKL9Xg5GldJ+0rS+2O
IH/0gBkWB7GbE2e+Z71nhRzuD9Q9WAlWql4RzoKZw2A2tA3HfjS/PodKjNhJWgTC
PvbwClWSAFB2+1qPGJFmAP61RGfSui4qCkYabjh+04O4DK8qOYc3zyL1Ma6UiX+C
LlWlVqYXv7DfBHL6DpKJyhgMAlMXnBkgSK9SPMEOqD9Pd1Ouhyws9jQCXZbG3Tet
q4A8FXcpj2ckF74RZpuONQzCTA+RsqcCbkSpQp9VI6wmQ6HMVN9ApLlxsLHHwWje
i8OVpo84KQRm19kb4XIq+wxkHLm2jEJZfh3UXkA2qRe7KNu3aEyVgsB+fBu+aWsf
MEHPvVwKb0RM71pUALEtcTqm+szl+6FLkFRyHM/VV7nOEvH18ztBGbaYIUAWAo9x
GlbhxgOCeUog2x6wlXbILHIoTr0PvI/3dlZKBe8wh+y/JbL7BAsr7VELMrGlK04v
XdZUnzi63t4hAxE32CVQjJl3WBVZn5aTlaEB/cCPBL4Md6FIPX+h2AswZBrJtpFV
TOc4NfUoRongPcRCxUtHms7jGLm5pdNyh/YV8Nk97EW02gJZlhmwzmtXC6p4h8Zh
NJveFZEi201Vu7rSCg0eoc01COkTrdeuqil0fdNFcyRwkR4FcSDjIIq6B8eJL+iH
q5eGZBtSCd/8wLexj5IPuANNR/M0OVUU1OxeF8O4bo/B4ZoJFFoSl3EcXVpKswGP
adoyH1u8gl3ckZ/1XoiugRav9fC8KklJ+GjZPIzL+mWF4JUbYYZVpkMMMe1gUkXD
xlBi6CsAi6YUsqLtf+eOLRvnygSwORn8Lz5ENQUG9Cj6JeKrnhLR70eA3nkVx/7R
FYWbbH3W7hnrkOALHGBCz93YWfaUUst9a2H5K/VqYpLH4TiBG2IadCdDUv08lVFl
fDLtGYLi70m4xk3kenD59RZ0VNm2NQAOcjHh05vkvwK6h2hM/1/P1NQMZcwkm3EF
o1sYntQWuZai2FeqsAS+r7w9lLGo7avJ6CaXgT6nqZavF8Zuvw+/XEBuqrhVCsbC
wuv/JFmPsWpUaJhFgVWGY30C1W/Lc4gp6CNjTS/kIgCN1QO2x4Q3w18kgyDDe+e1
TDPBeP4glabWzDwFpgW9QEjKoM2crLjF5HOIeDJI6N45QjezuFsxJYYNaFIzFX6u
51ZK7eNt2xiEgJJ7IlXpF4zjGPZR2pL/DGxXDfO5gEarYUsmMgYRWbx7JeG584gg
6z4gFXdDKhO3gPnaNj21r0Rrx8+TZuskcJdzO9/9rVGDNGVWSXtL3MUkAOLSg8yi
XJ8eeDQ2ztokigoyWK6QjnmPPI2zvz7fb3b+jHh5+7E4LyhRzX/OSML9dwQq9Yor
r3CbbCqm+liVo9F8iBA6sHIOPzIlMyGdNrBM9KemHyRVw6bQXeNpbdALCupImE45
h9bQvr3RjDJDwKeS3Vrrj+TGaWFK1mMc1TdNMBiXI8qLNx3tzs8OdvD5K25KT5JB
nuiQOeg6k56iZYHX50Vb54z/dhZtR5oUxc6wFFByVxjTUK2yFct+tVjlQ2jQLasu
Fuo89dDMoHh0HCIOp3ZCa2rXVsaD1rfz3/llgqxg3ToyIGcSGS6LZ0tq1O+NpcVK
CJI9CF9kousTSNrZrzvbJm/BZDNTL1Ql3fqOQTad5w4Om76ynGA4FDP5icODerHD
q141U8Jxbn95zvxnwjnNdB8gbVntktIzkRVbQ+55FaPi052jh6A3+sVopWmyOnZY
TfR/sVUMCM+5sDWzRt+GheuMWVUGSamNh/NnI7Ie8HEC6HnD8ip6VeW52ct7u4mQ
8DLLffweyotK5QC53oYoybhdPRlo1bNmrAccRwHNQPDUX7HeDgRapu2Pc2NaghyF
ReC+LJGQupDQ2G+aOy8h3eMijBOrKiGXq3GiiWiKyt4Fev1iKndTJoBR0BAJh6ZT
5/z86esHlPX1+10xrvcd6DAXvVzzQZikr3mmk+/lSwK0fjk8hh3TbpPO/Sgxjb0b
qDvnP5MXhKqyWLK1K48uAxcJMN5WEQPMezjqUajmMj1fTis511JpUYWTtRY86E4v
fhFYxDp2eVErV+wKwd8ojrRKBA1G4oaFbMvF2KeT+mI9Cn9NQPxhN6/vRKVZjMi/
RxB1Th6C8TYajgKhGveB00K+L2Q6m9Jr6MxMTxfVH7IDY/hBz5loySvFJz2X+/C2
xo9IdVUUp86C1lew39ixk3nG5EZJP0YOW5f2tXUBILLMfO31sowjj4yl0f/Os6ND
dHFBzLdRv0uiNBj9uS2Vv3fFX8bPNjFcOfLmZcfhx0wzbQ958YFg1J6iszSo3cni
rVXFAmNbl1kefaKGf0t3q4zuBSpentiEtsPwpegdC7kpOVKMofx8Lc5YJ4l/bSBr
yTF7uTCoPqlkg9u+8fJMZGzQtN5BTnLYEp2ckfkf6zedXkA5G4CamA3a/X5n7rKE
0Y9Mj9zmQKcXkkkXWaDobeZmdr25KYCW3U8l7Hq/rblSoMH6dYwaOG/ztYEb/Z0q
RgWy//v8b7qGN76fHYwvYSnk1IELYPghqLO1LhIso9TvPzxvaAbVNcfmxgvUEF1V
oKsh3E1nlLZcQFsY2ftJW2Sn/PiB4jtTWebKFi+dPh18XxV71hyLY3x1oXQrKn0K
tTP1dpfm6GFJR1/Xxuc+afNLhwMg6S4uXqjR6xiykBBHQaXZm6XBfTeAn6RvAdUQ
adGCCdIKsiyP8bMIN0CQE7FiaXpBxcyXqrQfGUDBfWH5OIx+BrBrBVGY9QjVrlW2
fl6z2yYuF+7PcbjYKL4kx+zTXZrpVENMVVv9Cj0fuPL6CJR5/3bwhrakxZJkvdFM
BQXWFsYr8tVQ9v9y678+0gDORfVAyFOxn23Pi20AJKa98cZnaNfHFiLgMtmRFLcH
72lk03/MczFybeO5nGsczqGVDhYzCNOXgc1cuBbsFwSQkbgwFl3G8rNI6RB7+i+l
jF81BQt+phWFSdG6yb82oF5IGVLe5pj3mD1BLv9d8p6ziDfFh8sL0iuVZgRdNFUa
rcyXLSTBx9xLkC0gDl+H7MOQR/DDwUuH+exoEe217LvGPaosvUUNgPnaG6E1tir6
p3ekzXhxpcdhg+2a9vrFegPk9Q0fTas1IEzRr/0xpm6KkfUbKCnKvqBFKo9Cvum5
36iJ7xGH5mlgei9YbwOzaGXLtD+WmNejN5pjPCVRQu/qBl6hAk3rl/rREwqm7t+I
su6bE9eTQVzAk+C0LYNy+oeNLxSvw7Suqt4G4zTj4j6ozfOp7/THpMF3tNN+uxH9
2bqdBObAuwYwiqdcLRl3W0eJ0F5Ga+afAsSsPNQbK/tVmMkyHeAwT5MgtBILo0vk
AC3wBu0POK7dEnAEMfP21+fsqR63ojzy3SOGaKNL/QFOhyFJqMwVvzViENvlLpL6
gbMRAeaXiTS/iMadV7wnA8BeKBIMUGJjKlE9y6MQOHuBzhugdgbIv3WOaW2DeKx+
kxUbDIF1vlVdvsV6Pah8KmM5ggW7tf9s4n5HkG09KG18wTprDNgDWkaN4agZrngW
JQsBMYivVSt5WnfHzFJaVeBQoU0g+lnjbYOGrN+lUie+E5lnq2U1KrEu1zwqfAAk
H5Aq5Bw8xxewy0x24OBq1unNZ00CKuP1QO+78s+xNjdS09uOO2WTVRGqwkofG2eq
6Z8EiuJ9pVqbvcKo6IfSMMQ4R6MdKFu6vS1J90R2rU1Rq6KlNtQEXcLnuO6oI2wv
GTkWWnenkFcSaMlc+3cw9Fj3Oh/RBuWMqZzEf7Q9T3iqnSw7EIbkCu/BcaroMuEB
1rhiVyrVdNy+e4o7VoXu4N7up04Xt0l1rn9zRhQB8UM07buForVbKdBiGnTygA9B
tJhbLlBryEcDYc23qqm6Ck44NQHm86m5S7lU4O1aF5HJyNXlt4BIGABfNVllBiUE
iMW2YyM175f585G7OJUnxcp6+nHCHIY1HxidkvQVa5Y1k2qnjXSKNrFKtXBbCfHi
v7VN8sRNoGA4L8qBU/C7Ewiyw48dc9fdHBFp3oTvN9+mNVNJuZm8CgkWRlycG5Cv
g94ve05hCQgSAiOPm3jpDQ+6U5pFoB8mnIgnt0d25Z7YNJ/dN0bjeb86V4nKJ1S1
6s+Mkya4wRZ/kymPO0BfL1t1j52saDG5Ea8PVX/3z7OSTSBLtQ6eQ1urRGGEK2Jz
5VdYHDkBCSR4yGip0v+YZ8Jv+3ArMdh8roWVFkFmdjNjGG/FL7ktRVuyC9m42IMb
sHMJF8aHbyN5tTk6OiB/pC97omGScEeuYetqWxkfBRhmiAfOyWU8TTC0anNvsR5u
C39P48Lz33ZECyk5mght6M7ILX1H7+Mij4ZFQ9KJgUThiP7h4dWVO3fspG7NxV7/
v83UoK+7RGR7fBqhB/n12076k9bgW6bGKhzEj8vL42fnD9d/bBz0XGrYokFgCmeQ
m+ACEuD62mGRrA4gCuoRgOXpPezIlqqDLyH7NFNeVSyr8wdPDw+UoPcyYxFDNJWL
gqz5E6h+iSS1vqrap4KG8cqGSEejpHRYRgv0Aai++2o2RqkOc61hjM3Kfv68gNr+
NYHgGjSRaLzIosNgIw6wh4a/HMDYdxmXnaszyUJZDxUMMohDqV6rqkgG0zbxGSRF
5u1rKF83I5/zlZwX9M58khCAtpghrPc0CobgxY0QbzroFd/bJeqhTardzB2gJebe
JzIKUbLaf++BkeYrp0JOsTEcIUxg64doFYMUCsVXBEIdlGQZw2salrWCJm/DbpyN
uJr+LzETzo9QZ9Pajm9V8OdBWZaGR35Tsb3OYi8qqiF9ZK0oJ9Kz5LInOSrsOyOQ
fZjwZgbIhOQZ3/GcDi8wZpYdU9lgGumwGNFw+zgI5m21hkJX95J2ZyycE+0nNsrQ
E7tGe0DJod0dDeTRypxNEKO3RhhxXBOWK2GujfaY5u7p0O026Oezp/MoXgggS+No
0KhIzHfVm5/wZ4HwfrA3TEa2//hYr8CAG4eyxqHXDwT33P5RS6pjd2gCeFdYJuBv
Pmj86dWHfigOdKDNWbIB4w5u2uRCTGZqKms9tq0T4s175gDe0YhTn96JWV4R16vS
zBzsWWK2P2Hv+lDWy5ck1BHRfSd50iEKtWzSE8f46ztVcQ6CjW0Iglw9MypVG2PH
wgCKXHzNdmuqY6C1SRoCVj2QiAyXwpbtONlG2oCppmSUEfsAKUha0tdOapWa8ljG
05Iz9oTTZJ4fJ/V7xaK3DFjKxTkcvTv9bXC2BrWmMAQVR73gmvpv+j7rWyYpnqLu
pTblytKIVpI+nX3x2A5gdawV4GB7IOVCqwvktjTmh7wVWKsrpjPKyGomQmGnmErS
umDdu3qZhFalKquIk5LcXlNCwrkXnLO4U/24CUCe8HKpDDkqOup74EA17gz1V71y
VFhen/TbT26MapeXwxe7lkPESu0rxyLB8K0LNOPhJjSSlbmxDVz9YoM4ZhVDV1JS
tNuC2QK4sTnVtzFnb0EtlrUp68LIV86uPqAwwK33vomM+XVFdOSVlHsou5I4e6mD
zEVedvFf7QhfOq+oXbY7iQkfSPs/A6tiNvaiSL6tMr1QhysHA6xVFAhjL24WuAgb
ZZ+azVMvrnUvYkiBeamZpOzAw5EokDE1sV9Va5apjK3kzT0EtJq/mqT1Zb3COXfw
r0Na8V1X4/95J2OA9g5zK0z+GejBDtPsmQ6HVpzqhybdEikBX76UjlPEyhuPRw9C
iLF1KImiVBjGPPyDiyTBOjlzJ1ZhG2dQjC2+OUIPRKvR7x8qCsBVSilW8PbCRl4L
w25BZr6s04SS8RVg1nL33bROY9OQj35pYALtC1Srzw7R8ucNrH3X75X/KA5qJbkS
DLxypWP7E1mqXnZUpSF3auN3fhqpZpvMjN1aTHxZqZ5O/dMSpJzCUN2GJLuzUjQY
oRs2IocOJe87tvjWAoCh/+MlCVbox7Ufw8d4rpCqpq3Uzf0F4Yq997taS4y6NSxI
3WR1q8RmiSzVOS1qwKCNb0BqZHgcCYskVLtc9Cmc1oe84QngfpSUvzcnxLxXInqn
xBXhXTQCsI8yFjOsbtCkPynoDRM9JNw0bfbflcnl65Bb4oc7DkQzRiRm1JQ9Y7yR
w5CWgIDJro/BTE8VomN0ukI5gbxGJwO6UZVOupNq7ztapbvv/NzkQCDlmDXfrInq
JaWWdjsJpLJ4sPe+S87XE28zD+fSxOkN2Bd1ya03eIpp/3HPSN5xH5t/NLWMXe4L
cZz7qK4FkqVw16HP+XGd3W/pYoBS1aLIu0gHg9uuPNSxmJol/rTGMuorIdJePEHT
+qWvI8koy7sa2DV532lA7DX9Ncawje+J3u8Fc+gZV8ncr10SfwIfRhxAAlc24lmg
sEwbVrtd0eLoVQmXTxZ1wSpbuFoM3IItvW4gpdq5p4WN5LNRIiD2mM9cxMIojuYq
sSwFEKRi1Yi17Cqez87uqp7DcpzS4YoLx04Z2/lngYwYXHlhjVZW6k/GMvfanckH
LsZdz3O22a4nvWUGhEQ4maui9h9JBKukSjDuivvtEKolnslXzVMK5IRA0GFsJ0M2
vq7Yzq6q9Jy92KDt5nLpzYekwjErkwE8vs03JUCvGqsSM7rsPOB5J/e5Kdpi/Hu0
G7OUUG5oomReyiXojR4yDG0e/j2RaAb/aL9oydGETGGGunDzyrZf1/83gEshayYx
kTI0PBfnDb2jLB6pjHkbRXnbs4lxqcZz5lLlw4/rM2x//06OyyWCzl1KejvGeSVe
yLm/b6Ep3xJKPo+tX2wyP5fNWCuJuaAVAxN/j7pElr/IeGIyuMn4ljYqvJdsGhAj
x38G7U1KcGAy7NPTTje+t4O0cM4HeaZRg3ZsUSgD3dPCmSVLkzNbM3ffyE7I1BEL
WeU/7I/SxDHhMeXIeec7FUwWFnP4PXdbUlYJoxljH6sn9F+jlNu0nxnLCnwtqQkM
AzNjtlijg2IU0LuOrxFWvOfR1hHGEQKWMt2qZ+VurRsDZo15BmY9wJo+jmNjmQLQ
gdqEpTfHXexOt1v05p/i/9rKt/I+61btrG8YlWssw7BawgLwUB3uZv9bpe2m4u05
aEtrg1V+jQLuPRoC8m16ZUCbQXEdB53xIGgepx7aargS3ntHZuZCs29al7Cc9c1+
E8uaiMBYzyk1V3RcOzV853JbNL53mEwl8dilLdaM0llH+sRd1zp3Gm+JT9TjwkMa
akCHWYiNQD9Yl7ej08SYnruN0PMWWnwC/motCpY7/cj/WMG/BtHNGDpmgYn+qOq/
aMKKZWSVXCVraZb19bqCJSFHC8U++3S3V3aEGWNLNxeRjF5GthpjrPoCXDSykOLS
cUIfjKajDxLxQpNNvhMg3+LlzRZtXh4bcgLQ+/Dir7eS5E3tJE24FVt9wj3Eko/z
0EmS0oHqE81LabO5xyI5bPD96RXhtGBIkaBEixKYy4Qa1jsiKLpHlk1EdSqkQCuH
Pi5V6VTOSWHumS2v8RWFUKTxdtX32gJhGvTGM4NFsTlZL+sVqIx+cge36zGjBYLO
b3B5BATQ2a47jRLMHH7OZYb1RCuflejj/q5ciTv9gv8PTn7NL4skeEUkl0ALatdv
GLoAzxD3MrI8ARAUTSliIhCIR4xx8pqwrRnh5+xT1yRofmMmoTEQaN5MqQXv9P/I
gaiFploruAIbab7wy0zgy4NOtLQpe1YfkBfyMAih/To7ILIQUMOle5cU/dDTucpQ
OZO67wKgU1oI+kOrIWIyIc0IO2S4wnXoKxN2Iugw0Z7GwCJRAlHlA/MA6NrsfdgN
mUIekFesfRCODic4NV3oB2ccWhKFrWsZYv+O2kptzGIdNQhy8LLb9jHuleED0En3
FjiQyV4QKFk1p+oRuC0iMPDe36FBFIGcZIvd4g/PobCIO2Rpkea3sVor5ynlwXFy
pLzGC0vXYFB5ehnmoyadEQ8I2nc3Hq1fW8TYXlkt5uaVsFNCsoB9XxAy6UTdmiB/
HSgzo4isvwqiPOvEEG33UU6quW00dae+PFQ+d8cWhxFxaGUKIRU6jSIGK+gRLigS
y28610x9FO1Zozf+H5KzmYJ0gIOcwTpJaIEI2nh+KemeeNlWH+IWfJ8Ug/lo18C/
3B9kY1uj3zNeoDNqnJC6Te+oCs6QNhm7h+MZ+0Iv0hzw4Rm6gWmCNynjw60ymsGR
R8B4oeZ+A+2LDRtTvnUIvROIldqJPSFwcSaRwtPd/3Xs3KFQNZ8zgr7RH7Q0B9eM
8YTm0wZB8qWLbUUAQpnfNcRB9oqWkLGbHCfeDY/qUoOZgSm/MHU5iuebxNS1UJlm
IytrPM2Ev0BT+Z8VnTLY171aitbD0WnYLKgd/DfB/cRKYNBKG7oP4QsuBDrPovOO
uL9SyfM7O2neWhdgdy0hUTo2vaPrf1ZhVWh/h983ucvroMXXxYL1MeyabwgS8OUU
U41IlccO87q+c0Q8SMOzIcWZ8TxmhjoyYgjYEjhG+/bwt4T/aNLpNZce81vDZrXn
zbdJRq8cIWNW0tJt7MU77FAwRZf+4VeOAW304ju888oqX8DZN8t4G0jGwb7gi13F
LKinTszNUJTjT7qqLxv4jdcQm1hYL58FEIDhKzdLknD2fEJTZI7Hm7eC6KDOX7iT
qQo4fP5lVdEA6JmEGBSdc1kmrygZxEYAx+HYNJt/vK7vrbko+omgkUCim13tgeRT
HL4T+P9PEoiaVyAHVu/uGZ0ZdthZpt+a6dt6S+m5lPYLjChtakPykjKVDAQn5F/q
MOAag4QvXGIbW07AI8HyvZ0K0hgUKRlHO7/4Sqt3mQ+Iiv3OAMS9pg1Yxk8sdOOU
AiuWk8jpAw120hq8aohwYap6IT2Xc/cxOGC1yhbjOlS6DHHk7yG15NZHyv/Gg659
jwxviqecTgskuciQa9f1ZMGS3xOnpAYxAY8T0oBVRpKO0M4ir/oKjdnImeTHJsVE
v1akXurAUULeU1ojOLAccTlpmIQMUc33dTHBgCNwUgxjDlnkXv3lxFTPHkwBnZVB
G6YPPfQZqARgRsxavUdFrdlLPpEgoWT1lqF7+KbzwY5IjOwA0jstHVf1SkRO1Tcw
X0ilJDH+3t1O8CZzw/Un2T8Z94thniipwaKtEaRNb167JNfZSUOpX3k9wMRQBtGC
HAwDrnlp9v3QksI1A701jj9/VUVPAw1onf3nEJ64rht4vrTSUp/wnZotNw4CK30U
4vPbtRZ82scInxFRfat3PdEtVFplp27EJUAxBwtnTv/4Wki3g4O8+Uk9pm+uIEJx
rqguqEkuHU85zx/oQvU31GB0Fd5w1E2P/SDdU/uegdMSjEus8H7itXGVUZuRZxGh
UaUZlIhtCB4Ow03Nbo2IcRI19zhEgEqgf2RyBIYOy2tQFiljigUzB4rqNohF9DPl
mxP8meZ7VzDdiTwhk92Chza5L81DmKTGmv75FFHZuTTLjUQJWolIL7YdwXJmhLTO
iMuH7Rotv1V9iQ89V+b7QkI5UESLLCTfm/xMX28veA/HxWFGsXqL52c7ipd9XpEJ
BTV7qOSXyBjZS6t23FhEiI1JkRVFV2M5mdZfImBIL8nMmTZKIFmf49+gvrABTCw0
epfl64mt6r6fhKozr3FoXopnjkPyqZXNPpxvR6yNSz6WrXGVUmJyjHb7vQDo+In8
6RK2KQQ8s71n2OdfFugVCkv0gzwa44j+Qe69JdwnkL+/dJu2eSqyUtCVa1pSBTpb
q6fQq+bHISxOlSRyLGOqcguiX9FMjKhbN08fgjZ4M1AMirjcgsVXiGauPMWGGp9G
vCvFNDix3I7PvUYJHS8L/YuZnx/QP2+jxrN6n+kZgXR8F96NnKtaYPIETGkRWj7j
09FmVIOMOi20rTCsdmXgEOFG2XIm+Epf/dPOJZ6fqiCbs5Qkfa7O77A8esIXbdcD
zXJ80T/1oMY5j6nqOSQnPVcEXxzmBLVMuKJX34fs3z14qeBJ66wejvcbTTh9UIB2
OBpFAyMD6tOLt9v7b4fZ6op7pMm6xCDeqhskuBQIjpCl5K+d934zIkQ7yLr7fH/h
pskvQUlB1OeJKY3Wo6WXgP4Lb5L2LqY377CYCPH38QW0FKIxfLMbD+E5bnZlpOhG
TRJfZ+n0kZYKwUHXc4m4BqdKw3kV3/A+2tOTwo3FuGF6g8hmg+fwF1p/zxJ0/AMW
ggJ8lTHJRYnpdk8ctgK4H2PEOkJH9iKGc1TbhxkbQLn6xEwKpjbbuBiQQ9A4e0+K
fhirIfuSsmgdBJBL0fDknu3FVU6El9jJhtcQeUB6mmC1PWthelmWv74sQEleLfoF
POp7ZihUrzdbK0bUm0E0M1nYpRd4E/pMnUo7dyxmpKH9rbYeRfolhiAU5CTHkSCu
Ehj5qAGOKXf6rLdE/mgEqjH6AR9QicXJLcsri/N22Q9wvKqFSieeUt5broF+ezvw
gm0t3RTkjaD5FF3Oh1+n56C47lpoW5NGgp6ARb486whkzEg0j6rxN8QNB+CwzPYK
8VeHhjWhCPFm4Pzy/Kwe6Ub+PQWkmcN+upBJDdVtyo0bvmr8GXA2x/8bL32a9z/9
PCTVM5FRSx+Ypnz+ssq2qCvJVP4C4RCqi6vC7XYQ+JSm+r7tr8Rcb2LlhZ+Qoljk
Ot/4g2LHg14wKkaJ6cP9VWmIKgAUrcSxUP9qVhYzPSTlON4Np8SbwzisLYEkkODU
PJYNGc4fKYf2deOFnAQru9ro1rGAICviFtWlnKvh77jwOb6A3iY9rRK0QZZwGDSL
yM9EwTSBzkAG16q4JQHlSdUps0NYJwsvE8vx9eywx1HY3RQDR4iDV9nE32gmeC/X
0chFBg4R06Fwten7nS10odGxPPuRRakADqcZX3gd0kgXr2gT23/jnmSRlM5bWtRG
y2UcUiaD9DsMmf1XvMpYr3ZKkMEoBUmeR1oSnKq0sHgQcI0miPpzZpeK9CEFSVm2
DgCrUTktqwsefE89UDjmA3gX/99b5Oz8d6CjkfbfbjZx9oyVNzOPR+p8PfjN39Wu
zHJAPcfg0fOP4XOb8FM6jeVKn26HXa14o1hUr3bB2MNTsfXnjuPfD1juJA5vf/gX
ucJOjSmAkc4cknozWuBUlZDNJOoxhB6/xp37a+JJ/YDHr/uAP+LNS0lsd8xyaXfN
qXKKR7TfQ7GsJtUd3BhHbnV3ahL1hDw9orTvhxjnb+8B6yBtx8BsmbUoWPqh7Ja5
y6GInShhEAEFNXJNZZRgegU0P/UIQbfPJwdnahJ8CdgWzEAhmYwPt2URU+ciXTU3
IWVUN08nM/HQetAyizYcX389Wysk96dgMB7t0TGhFQgRKICZ2v/LW8+nUSmYnQJt
XsrvVqOn4G2yVtcc0KXh8tX7TeX2wsOEpW9CvNmNHbmKbisfRaQKrc+UX9RzHYlM
O90LUUn+LDHu+4bV1o9Xt0JBy3yZp6PrC1EQln9uXWOWJA8wzbuQGoinuEidLgrD
CY8yNtN2DP1dJ7VB4FJ0sNEx8rEdjUs9MjZOF4PTcXYOEwPOT0K6ORbfy+u3TFE2
xZZHqIq+6wNC0MtDQ23JcxuHC/GbUYtFGBfcnPsxsqb53ct6MDVpbyGQ5eSP2FIu
wnNeTQrqtzFagsX4GWUy2UfVJyBKDsJzQLsoOiGrOtwriM+ikqFjWZLEO/VNCI1d
EjWazWno+HWp3/qH4nkijhXKI06weVtssgNXedP5L1GslwzqL/sB594xTvGo94sT
5813jfTqBK/S+t+GMEI5s31KJ81gQX+kkIFryy4NEBVbvqWWDPumP7zWs+pb9fLr
bUzufqlcCk57f/QgGqspKA0zJ4RnDywThL/pCY7TvC1cCZgRS4T5qJ32fPrZydjr
2LHmFSA4bXKduG6Fxn02bBAfL2OezY8Zzj2AUWYZcb0GLZbQewAI1IZDtwR+s9f+
j7msJ+tOIwjMgEo0NnUaczSO8XAKMbZmL7HeYPlETgs/+uEdKjwnh/SRSXm2FtyB
XkMPEbeW4ASptTiGyqxNJXt2DrlBHL9E+mRsl9P4TdTQVg2CoJPRPZjtAclMWKnC
Ln7Qh4kI65GS4MhXG8IYivcdwzeZpGU3XtZsT+SGZa+XJFjdj2ZFuOliTKeeOZVd
p/nHuPRRhm83AHFFTIXlB4YSCXXVcjs49gyymF51hRTmsQpoAh0znQOJwUxIzmk+
4feptn0+141Ky0ncUpJLQj+/vECXS85UXB/pLYXtOvhdW6JP7sjKXRK8yJq+X18W
b7vyUDXg+6+T4Utv0OmweJl2JLdIlDbU2aCVPAwRie2x5BL84kt+plMq4cfOJvEV
1a+4HWpDFlII+QYlF0JuDO5BA/1Y/QAWjRMdgCwp1TeJ5yIOyCWwclFFMCsL4sR0
EfRaAZmaWvpHn8Anqg5a350+aIeaqZBlfEtOquBevPpk+Q19YhDi3EDjWZVmOEuS
n7+hHa44mGkaFvY/xoKm9d1sQMR3fYzpC+eP8Dd8UNHT+ltNqf7s6+junMejt0W1
ekeueY18QA8pFp0lzztlvLZ7VxIjRerOb4g3TfQWe51EBt3+wJJa1CNidbl3rOa2
CTlfdqL0iPt9tLUSQjxI81ooKoqpgWfaRg9xBADNTu/YnuTbKQGD+s1qVWGYqowF
I+6qPFiXoShosxc4fpwgpSa+uHdIlYKn8PcQMhljSyR9KqJLCktydrOPx708nWhz
2Hesw0yq1Clr5peT13KxEFy+K4xXlBQmLkstjTq8swIMReDFZOifLclKdY6iJ8m4
XskoNnZQBAxqnbFHTINtR/bgLGtYn782+uuKrAJhnB5aeDBd6LTIu9P5D6ozqjkM
2y+y8Dpm6jjvCTz+Y+aTJBRNjlG8TKcEistKR5os0qqCLkqQ3g5eB0NNOFL1gDfx
ZisHdXXT5zbZPzyzDnhLwfuiQiu8NVBi7VtsVzdxtjwo52vEyhheBZXp8AmW4lUj
vemnbTORcOiqmpCHMXLX1DsUqoxFIzbsqW9Qlq2HWlDL+yr3T91qGqbSYV+0VCal
yAbaJ1io4TdBVhP2RB89q83CemLqVC6RwGYdDeGoJW4ltL9Yn+/4zHhoC8CUPtnS
RywwZBONp2MReRasQVT9hqtdCcMXSFBnh6ZN8+gNWbChy+8/bC3QK8NX749b2bWb
a6T7kVgLa4PEqq76jq7+82wHaOHWppYKtiJ8WwrystOIv9mgODpC8K7W5qgI3ftb
6TViopMp5UUJSqYjgbH86Co3fKetpNr+xN9024KDgWKmgvG+0pR+xmWcll20wUAn
997b8O5CvpycuWra2yP957bDErkpQ3aKMccfH4jY8Kqd0nFUNQHhI6pkIDT/DloU
CT5TCIDryU5QmY/XLl7VJ81rRpz+RVHde1kvIM4k8y8cGV1jhDHoX1e5f3pmZBEN
dZfc1VLvdv3DyEI4UZYMHoZp9uSc/QK3tWlO2Yu59u1Hx6sVQSZo8YPci/Ag717T
00iEAs9X163kwJe3Zl917LhZk1TX6t7VGn2WTOIFSvD6RFiCQW4CnjBHwVLdU8V5
GPTWF1ya2rvw4NYczi1JqwBGobBax+JrCsQzG6U46Q6GDAqHcteuBqHmaJgGjcwH
kL04cWKEvDqHqg5W72tprwVTgntcZkOMPSrxWclBaM1lse2raOBYw6J2Iudp2aIe
nLmvDrbUoVOY3HeaUJicRbLMzk8kSyIR3ZE5ewI/XXs0DP+je8d9M6uEjlPTfXXS
x8+4N5+MSxDOyFXtB+N7fkIlUPAKyi+ZEpKJOxOic+G5aA8hrn7cxXWH3V0aCirC
4WLxHU5CT1c2TsG9Mk7EMW3g/4xnUxk+aQ8ZECGo3ajAZbRTaP7NF4qjlBXYggdI
lJsu3tAZCy7B4UA7ZVMXeI8iGe+jMgUBZ2YASfPqEADYHYGyirTlc4jBqWY/ZYoa
a34K0PBzJt1CkJ+QI54qH+GTRBO5RJsiK6vl+w6kOmYRXTX8F7EFSXUDc7j8s5gV
n6SPHHqXMhxp0Asr61LUhOK0NK0SP9nO9p+/o/5tE3ZSWKQOOI6RhI1z0n4pWUR8
5IqqaLzmmEe7FUdBrrNmLlEksmol1kUKgF8G2MhBiOf6wkqTed1LVHewaaPydEm5
coMlQOs7QdiuvVmL/v5hRbPFv2yp+BUcXPObrVxTYHb88PY7dcb8sQF/F7Hc/SNO
nT3TNUfHrbWuCJNZUW0En+inKYYPKLKfjxzyQNNsa3i14tmfOzCKX6vxLHp+D/+k
ionI0n70hIr6zYR2M/gWaeUrBJGgpp1PqyB2aFMwxELUNgqy8NjY9zHkp770kIRV
FUby9826BiYj9FBJwaSeClHx3IFtcs2D+bKDnguruG3p9Xbt01uWmUNtuGl/TYQa
yYFDbXvL4Eog+1+64/7UNkzeMjoXgdCvP+zcVNHFZyEFb8eDzWNnc7Uanumq3NjS
hf0xXb+QYV66gM+b934T3S4XpoGFEJIOYwPewwpn9sKkyk8QmYU5Fen0W9FimHQz
6ZwKyIZwHnRdCgSN3cPrVfCfpfx3Xkfav4dCyL0YoLMwYPbK/zzrXUY2T2RPHog9
IAyTC4fa3ttqDY3ANhfsloRvH6MfKw2yPlGpiCEFn1NFUSTabEL3AvmDv8cyCbvy
wVL7u6Ar49E9EiFt/ZoqYRcELbBQh49sUsb0W2QhCW1LuZzV8W2IlKCHlknREO7h
d1RnB8Cfhl4UVpM2uPEB+CJibxmNaj/S8tSybrLOaXYKORwtVRztRMg877SrrjyV
uC4Hqcm++FEeWFjg0cgpb8GpJiGfnpX/ubi9U76CcYufl9qa2+OOnBT8r30wb5E6
WG0AlfPhTAjOOUmUZe6QFhNImTkMtL8D3sU1sREsmrqmfLOaJ9lDNlegtsNkjtup
PvJu8LIcxHTd3ECXEs/Pl2sgwszHvM2Ch91w0Ni3oGkQCUm8+sLhfC1XIAbuY/lO
hhmB8n6u2+XSc2pdgcBrgmZgS8ZIyx4wz0JtwtbCTZy7uTt9I8wvjh7i6dCVQA3U
IbuOUOoriAqjmrcCkeTLrHYhOPPetgSVRhIYgjd8px+tQUCIgfK4FYU2/+spn+cU
RpHoREO3xyZFQ0+Tvka+dXqzQYLCTMfX91VqBKdA0SEo9KpG7qHVKVq5aTU3nEsy
ol1PqB06BfFuiR3dusrsb4fuXQ3/3UyskEh6rI0dTbqjatirhhlBoCFu6oNWYvx7
qE60dhlmsf0bkt//6TbwQNC24D1IP92xpaleiArzV5PTCYjjh3WQ6SvnxzQZSnoZ
AtWQtOoHXvgrfdsbfU5WrfI1UlQiQ4ZWqCcRTzk9cQ0dVVNQpvPp6CMaF2ycpIPr
N1e9ADf4RE3uB1X0Q/kUrh6yKq06mN4d7caqupedjUj9DWoBn/fZc1gop2lTjxzv
yKFMSwUB9+m3TZL/+AB5scAuhYsabXlpI3fC/Qu7aVWGPkh5oZtjuqnBLEkLCI0D
STijqG0azbmZoJMnekbh4huIyauRdLLfoEkKfpBG8ipm/JIaWzEo1B3/ogWKiI3a
KEf69Hc9RV+sl58FuCVWPE5Gal6vXQPRHB4+gi4H7hy91XLiBMuadJq59Q2F3uvP
3Z+2GDql4vhLPQAKxZkQxEKL5LxEnLWRkqk57u2V/1jdH25R9jTUbIfQsiXlS9fo
WnIPczjp1BgIbv4qrMVIiZjQDHVBVAMOhNSHGUqeFIT9JVuROWgSAbaJFAaWddAx
KJ+w1IFbbwiM0UvTIoYiqTX1CxmP2VOqN2CDAaWhCY43i7WfAfp9JOvjp0d0y0cE
l0YDgoT1hX9tov/ICxjHpLyq1xNBFeR0/nw4NTL7LF2/80Bit3m1ZRu7wvX8ihB1
ZQzDbpFFqZ4/7eX0BEeg3ulHIXt8Jnh1TFIajaGdJNhp6U7A8e8v+fo8QltQK/IJ
eY+CywkByH8GfCpr8spigGf2Q7toKbfUyA2NtzKW8OcuZ1mP56iC6IozUdQVRAtK
YvbuChCK8NPKIVtx1lt5iTfdD+lmgzNil+rv9ytm9MDn3on6HZ5/1BAS9pcSx6ms
A1MDW9bsPL4ZHC+GEma4gcCD8Qt4JU2Y8elhmcQWR6O4JMKeaWYO40bZFq1s6/4s
wKZ7TqTW8gssDQ7akuO225vHB7esAbl0kObNa00Rfseaz/zWcddY5h6lnC6Ilkdj
OjIdbxYO1PqYgnYobfj42luVRse7DzXX1WyCZ39xprwcTr//GxabeNyzGK84OL+4
Qp2rvWmd1fu8QBwcCc2gOc6HJh7rHXf4i2nLtMCETa4KZtryK7s4ZN3BvsM+44TD
4EiBRuV2744n9XbV98frRAeaWZt/RbDJspp5pNrOqJlloidrH9FHVWTzdQO99Etp
G+2rt+1UZkDqm45A2qQgr3HOAFmSHh5ps3OlmdtrLlV3hBTMqHcnKctxZ0o1b1AH
+kFEm8wVobE6/NKKzydH9i8OXxWbc+icVK3EowuRAj61sJPnBM4GSnehFosO18YP
j+TBuSimjtuEbHSElRGs18lO1l3AF0m7SlHqPHlCYQDoKcWzoCgpUQTJFmLkER/Q
HkSHSTVQD3WOE5/WcAAenzNxiE8s6kwi49faGSeJaFpLJLElkU0Ygd2lVL2H/Cb+
Dj4cXOi59c6x3Op3KaP5w7M4Gw5X4Q1mNfxD3z5GgDD9YJC/HQH/sk1PNoOATLyF
qQOV5A8TMdXp0tRmc5cW4jamnMgpg5kmcW/uY45vinwYCCZwEU+PLZ/kNeGzdG0r
JiNPiqW/X7LeqTbNrr+c4dpdyCCLrPOUGcNjkWsJLV4EefXZ3sdrQfvEGzt7XrPU
Cu7UuuaslhgbL7U2C8Sguxqy7DkPCsLvykeJJVsmsFvf3C7Obm0B3FDf6ecY+bjc
ZvHWMJZbmKN4uTBHAr5c5uqj6P6cvJObmTYvRDfvzqwY0TNMXNjIUwq9eaJAo2ky
/jqgkwTbzKjLms3oeV0A1xCAbxYobqsdGkT0xh50aZZQEvye5Ok0w1t9ACWFs05R
PIgSNxF33HMRq48oJeiil/AKrYgA+bdExhRwm5BkAluJPXDQ4kr56S8cQ4FioqW1
7uda9t5zRpMnYzUcnJclrZUjwmfwlpJMXpYqVprd+oji6/KFdYi3pX0PGKcARgT3
TVBEyV7uj0RPV1iPhHuWWHriOv/xEI6rhlQe+FBV6SlCEbKjbae0LVuaffP9F260
ZPCEcBOG14iu35rwoRCHTxvS0tNedjBvjx4ac3GXjpokTYKu9wm+QxPWmZQoeOFd
RllpxyqvXxRKF6K7SM4XhIXT2OPGJb0xsGl7vJSsuxTJ+DsDGtcj5aeZRtik4WpI
krYBFn2BYoVckLEYUhAHi+me5U/BgGglR41D6CeqlM9I1lEpjHm+SszIb00oqGLe
WuN/+8zun67DY5ElSKtbu9bIEoyh1drgj8fj3nVqVSZ8zhbNaNawrSQ0nK8HImqc
izW8CccY1kLIP9B0/RRxCr9d8RyHbe4cA3gMyA0eM5JBwpXFHJjKt2zfhbUAV8Y+
3tA4H0q7yvXcdq/f+Ai8f75VS9P0KMPX4aSSm9M/9LTTjsJuqZfDIp2vwTtfapP1
8ApbyMViHI9T7gLVfIR+nwzvgX1VbqzS0DFY87y1NiiMuDYDWhc35Gy8hd/XpTDi
scpppNbQba8EHNCZ1zg3NKigB72t4D0SzsYmfC6wxCnsXSlmAVJS8qdCprbDYZn5
rwVvbehAACyGhU5+cMkZUbe8MruKlwoQaqwbIQJBRWzL5ALLkSz4pWOEsI89o1S6
hasp7s85+nxm1zjHGADx1udVjmHljgVy5ml7rpn3O4Rk+Atkjnde7CAyMIhoRW+S
iMiE1KH2WxJcgqAATAMRT1cA5EP0/1hRRMMnBQ8JU6RL/YTGq8sU0EImhwhDzshd
lQh9bjqYux+4IdSoncNQr0e4n/ST5sSR3bw0ZlQbNqCiPtIxtju9aqSAxKO1GV79
w5KFTdN3+kcfPRjz+RvLfj36WNIlxiUSGf+U3QelOkNKeqsiIaO8Jz9rxZpBjZHY
zQIKuGZSHxuNnc2AJGsPIjGUaVryw/U1wFcENmDibQCBKlz0X+QhrfDzvTIveBf6
CiuzEAh/5Ocfa+h/nwH9F+jFHCchIZikLs5U5wKZ8TRo3i5KfvWamrK92n+htwUe
9sJV0WT38RQFL2QOvgP/wyAoq+n7TrPiY0cztdME3EzW0df1lEPB9AXql5vS1O0v
/G5KXgwLRA+2n6c2vKEdUbipx5bBbQ2CsqDOM8aIQnDJ40wPDPqdB4a1MEN90mgr
hKRGNjV//p0WW4uLRcc/mlDXimZyyAPLhDCk1vI5LxooAwUAaE38mW8caQjvehIk
JAPNG6fQy2dhK8cyNdyErAn9JoJwSq4sfBs3Qxqr7IoLDj2t8aIRwi1ObUY5TJjE
RNejgHqVPh/uTd7n1XGlag9SXUTjVlOVFZSXsqYrcnQ/3Hr4dO33+A4K9w+beTvD
URA5XYTHU/ofXRCb+uqHaiBIYO0ERPB+hPMSLh5D4kQOxRQETv3O5nr5l98IYBEs
ngRI/bdoswzJo/R0noOr2pEewawCCMzVDw+eYavQ7rQN/NF0/xi1Dyz39ycH+lNi
oPfEPZ49R7FR6yYs3HS1GJIQO4yMFCV0CfaRjLleQvf7q+wlItJzIXyQC0dIir01
RXNB0Llmc9s00NZlkXS9lbNISWXv2tAEOr6ePhVNZFQP526HKA5YPyUDKIwzVOeN
njof/jr4gTvfuJcw0ZBxq3+ynrXFDLaZZF+PW9MPcf0aB6jw1wrskdm8pb0YF6r0
aAspIL8FF+9nAMHe4uX9B0CaHBm9Y+x41o2MAyZabN/2G8LMPPPWqx1Vxu4zMcab
3AKQ/A3HUNi7fVsuainieqoEmxIP6I3eGJ+R+iRqxL3sOkLw/pev6ZBjB31AK98M
yuZ4JXsUxsVTZ6LvrRZplSeZA1FXjgmjy8CZjVGsjbCarYVp4M3reuKjKx+B56TW
Eg9h8yn9XeCFkWrTuZnG/dcvG6bL27tbI19oaIq27PGLV1nj60B4v6ZP4pAcagA5
rjoh4epevEMtI83UxlOY4cP+wwZ3BFwLo0TV2NLvuWANpxqC3qfvT3X+wzVaQEfT
CpPG7xTJ31ptm1vW1A6U37ZRaz2mrTUlG2K3qC7u+JFkgrG8G9YAwj1R4dL32vfK
tT4dDV31D5Pm5CX2yTdVr0lKZs0n2GPdV6R5kDQXhaKHwmSyycrrnqbY5iM/YGRD
TfQNV3HMi/tv49gkIrDV+ImzGeJ/I9QCVn32WYBhk63Qjkg1Pfm+IxNtSIpyXAWh
4OOK6k4uwKG/ThlRdGRC8LcWq10zJvPep7vXcjVp2dbGx6je4Mbk/XmVTEzV5TDS
LN7HbWzPRbGOyknh6GIq/yNuOwzBb/7/M4r2dSTqup5y+Y5nUfxFuM75OoCSaDgk
4wftzSGXcTnsdXGls6EnHg7EDhXooROiKzJHTbynH//uZKs/XcMvrD3LoQSHbXJF
svaWuaMoh2Jvzacn3IlSkBZCMOHoWJdlROQgdGSiCZXvjJVog9mXBMq7AaUCMQtx
rxv3WLk21a+wR0fPCV9ACkey8UVt8tnn/7IHJFmQXcoHF/E5Nk0xHTBJilAsQYoe
bFiQlEARXPsqAKL+GdFtfk7xn7k8v1AuiLu7SUbiLWtUrNNq1fx/yiw210QtE7hH
kkjARtYTNOjRlIEpF8KBK1GJToIfovLqXlTQCAVdF2HqZR0gUblqpW6AWIAMVhde
G3YdhFjq9zM0jPC0zPHcGmo6W4DJl5xqtYxttv/6N0/Q1aiVvBZvfWT/C/fGWvag
nR9Kid1dlREmmDVr41wDT02NUUjJtNTGVS8yLQxHPvvqDto/Mom9vC/g8LqPQ25l
YlPfEmOFUjkh/N2PJHEJFNUpCHBaJ2EJphEsHLmsYrkPKF7AJ2qzOqOdft5iwPqD
YCG5HONapbUfRsOkdHP2mFH/snv/q4lXgEq+XRB9xkjcaeCKUfgGr6nuagHDkpO5
lNJEpfvuMc7QTfzvDQM/3asEurTDeEbACy0ckMj4pNJYtZYyIBL7cDOuwfU3Fuv/
z/JDPuRF2+m9UTPCX+kJkN78tPSUTCVYJL2eujloR1x3ee+Hk3rtchP8tvT7j1YN
/K0aWS/Rip/YMS5an0ejXAtjNZW/sXhKYusZXv8QPy5mnEtoYnHrNLMQuD8VxxNR
FsKIonmtphXPsEVdvKMAoTC1q1e8rLZ5I55rDmPXkP+l1H3aS30FD54c1nRM69nC
PcqvwLzxoWrRGeY9QztLGBPBHjTSIlnmoQZj68Br2B8XkMkK2dACMB1FQR/XyywZ
Fh9YK44lIIAv7kYnTAS5hmNya6vBO9QzTyw8MwNDXP0J+TFHm4+frjhxYsh95q/w
q0sh2l6lw/uakYqkPz88+kyHZHQtCCPDh0T0zJ0WzhCKRALKv7E0tiYugIy56P1O
/GlmMeepUrvStMsX3wvMZmJrXSNt3G7MEMVe+VW3aTd/6S6prjTVm6Z+ND4HhS6T
bVHCPlMFnGy99//Ni9dWfHuYdyXAkv8IVmw1t9LKrzlh6z4jo4GX/KT64y5Arau+
ZaPBRwalKL5XssI1OYF2jpA2y/mHug954G5zc3o4CU6ttD7JKWmJldBPxGkVp0mh
Hq6yZBmuQwhoCQrMnLOkpKtgSCWAUiDUJbaMQ/gHfkXzHugof0jubn3q50pumJ73
nH1hUNs9fNWK04Hfd8I1YwGVpn9gaBp4YsXw482IWg0J/NILLOvBGbNgSz/3fM5h
6OLIBwYd3d1Zn/NiOe3C5Rh7IBNLacAk42teGcvVV1LK3u0fZjh90g49Hc/YB6Lg
sGVvGXaOoRm/nMOZM2ORN/jNsfjErC9v8IsV96pY1bDscSx2cHnbcznJUFsfJDLE
Cl085TXMRhJOugXlqHO/g2RCYTYpLxgXyRUlJwz4QeOFN1DEXrPRGvUD8SWamwOo
iDr3J7/cC03W7Tb4EHF4jI+59ofmUZWeGbginLS8JxRHcuPFn92W7fts7qdCG7n0
GgNTMLQskoPmXDDXgicXdxFtkLnt3FB5GYAx11SL0Mfv+dMNqBEiUjZxCbM+T0c/
bFD/mNFlgCB3JHBffSFzj7Ivz+PW3DIQE7xPUJY+jS1cDjBaSd5fK1MMCq22tKKn
w7UaeMlPAcVd2GnKW5YPlFCNqmQs0k4nwKhrd6ybIWEwg19/ZVXfiAIkRYegsjwv
hRM1yq7oFrnp+mc2uIh6UDcwApZ0MBUP5s9427A8VrYgjoaMSxbPA454sxins4lz
WcG641vyMSlOCnkJOinzZWRFUAB/0uXXrEpLX5+abipMIVDYRdeITKG/vfAF/S88
kkJR2dJKghJ/ktFdT4x0xR+xaLsn0TJ6oGCPPNErMUCIB75ghMoI8kl+QllWjcac
fJCJXuA05+AODHydURZm1JXuDEnh/toUM+ehlIvL3q3JxwUm+g2thyp0xWpF6IMx
FQydKBe0McQmnG2D56GsHg+kgAK7c1ehm3EFvjAlebshuXlIPcp9xSrRLOd+62lq
ndbocBNNf9o8YCk30BRNK7NcRd1D16jIfqKyZ3Mqjd8HxjE0Y7xhckcNEKUnGAsN
+0B65gXIoPmrCHCkPot8KmOuLMnh+jc5NgxmELODpf9TjJ+lbUBGcc6dyfHUF8Iz
fyvAR3rpgdubgnJqRgTioUobt/Ci3xCDNRA/T1dFLq6SzcS6G0fRX8+eNgXXpj2v
ENyudKQdjul6og923cwhlnN8yW05u5s2ebQP12p5L5cp+EedAkj+MHDLy1Ezyx3U
Olv7nXsK0wk9rmrhkvfgoLK0uhBwoOaV7ZygM8P6tkvcJk3uJRnqAsKZkSUb63Hu
ilN0Fh+Gl2KwLYiNngUlxP4sIilm9I6bchWYDZqBdQt3m74F90mYZq87VOhzLDBS
n2aSmgYkSXDQuGgizvgHDOvAV9DBmA+1lTsVAkgmcbLzITmetAI/zxA32fcVivpq
uX34XFfLAMXLPAexr16E9mu/1uaa+aBQ6wuXNDvBNm6i96vEaz32JALErKqxY696
Spl7SzSZth55WQwi/19mlxgChRP0pWL9rqtwVslXlN3+0WKQkZ0zFDyr2EgHrJGd
Q7SDSVLYbxD5V1RlY0LJv0A4fBE5WOBIg6gjZ7DeLTL1y5fo0m9SGboDBIgQBlAv
6Dw4wEbt0NawGVGKdVF/dHiq0hck0pHR0jAwqPGnT0pbZvldYvK90FN4IgE1Jl6c
pwCCyiER2PLB+nfSqRhcXTUV1KyeGdXfSfWkrm4Cc5rEXP2d95qisFMs0ubK3yW+
c5/PG97ewBvWZzNPn4vLmyQFuyfaP/0gjqrT7lU/H8bgmBWnQJ4V/USmGfs+ETgk
a9soEUgrhQjML/YKZ1Ge835VnYiBu1Gg1aCyPj+Uy6JyurcYYqhyedqXqOIT+auG
PpkZa1qTEabefXKR9nAuVTckOs74c3EmNwnrnZB0bdL6jQh3KhqJaKPkUpG+LSYh
xMcK3x6/YaQX8fh1U2nGdhLPIk+My0pWC1xhQMGoo8+XOROlqh4WQdACiBPx0AWH
fbxnrq/ZzGIwlK+yBFenuYVrPFceHi3tmNrB9CpIUmgNx5xo/JOvNHDY/2KO/we3
P0KGGTibYP2aVuw+VzoXeMK4RfHdRNDjaDR+elHw+0Aw3p9yYCIKeRGNy/O9c2mP
/67yVarKuBob18Y9U7cheqmNUpSxgE54PxTmO1AJ/hqVk7ZYxiEPa3wWj3V/fbYB
91P8uQIoF93Ag/x5A6PCM/hv9IWT6T0yBNEXCgrlnmT4OTDrVK0zAfR7Uq7jUtf+
XN+RBGYDXqJL067e0HJecOyjHg1CKBy6bsrTqalBxSL/ohFe99XaNV19TkIQFOiU
OZ8AmUfkjov5UMXIFRYTstj7JQfnniT4w3dI+dWC2wZgGcawtOttp9wtV7fJNrc5
lXStNI2RPJBaIgxt7sTq0HEouACaE8lJXUSLsC/3oOBVsPlkSwg/cBe39ESNbO15
wysk3re/2WoKr30XIFfoa2MDZqk0G3hhcSCqzbXMvBmrvLOL/VFjJigeNwoKkP8g
5QFp4ko7LODSjIn+MxcwWBApWle4yU0LcLYLD6AC2anP9OnxEoVYXWhbGISWzUEX
DHNLWNQrUdDZnjBNB8o8kDbNxiiYeq5rpyxJDs44YyI3lQki+mIuslA3H1SfPT3k
nsn0y9SODpGuvaUoEUIuIV1ekgcK1JZiaMc2AzauUdRqR7nnw2LznxIe9cwAjiFX
6Mmx2QjzHx/ONGdeZz2FKuEq/AvnrAMGo+vFkaCmF8DMb+UNAlW8ZuKy+Q4AjhOW
zvs070YP3WDJmuIiCKArPQtbvtGOT805jlW/OTbDLfsnUnsaRb0/gy4JdfijUZrw
6zHU+GJ8kNp30crrY4zHb0OngtNXdYLQFJav53fSZlkLzJO4Gi9s05Yl4N3GUJQu
KUcg/ne2tJM6G1hiDdQ3e8J5FcvXah+w8NGjJBwB79SwnfX3nlyUXUnSnv6a2uvf
Spqub4VPiz8oz9kvYp9jspOOQtE5ucIZzF3SEWYE/JCyFKvSnWfaA8oSWtKVPKog
yjKb3hygNauaFDEThUsMNRmf+fQ7+MPNkiKDVHgx8T6BVVEzSijjVU6gg1aay9Dj
j4qJb0WZGQIehdv8m/KEVlI/BdcAi1AishZ0HA87RPk7mTtuuAsfsatlX1odEJJ7
rU023D17jyNezh6tH3XwFsR9NEnfzNnWQPqyYquIbDEVmcoFqrJA4zo7npngej5+
HsNcYLX6Il8RtH6Vjuf/JH43fXQsUagBEPObuHRLBQIYwwu6sDjPbpBSzuZIDGvW
w9hkWD9VWzg1xSF0nPJnE/6iYrp+yhHLEQ4fR5ywimKY1MHSueaMluOhRnWVREli
XRKZvx7TgmkJRRLVxC8bY3rwrRnV6BVD1CUaeeKyb4LFRXsbTl37XZfs+WcU2hrA
Ja9Q97tqJ0sFHTFo3Xago49DsBBQZvmiYsusZZgD1wiidvaM0/zMHQ5M8TqHJgT+
WLiNVcxnymD9njmZe67LIiO3zmGT/g0a0OhNc+yum+4+p6a27YoD64dInEWJnOpy
qqQrgVT4lwUVocM9g9pHDpCVSjxKwTos26+lkcc4an8z7FdOLCpF67wpJpzpefOz
3S0v3lce1kpstYup35o3V1pMXKPLnrCJAoS0EIN5sLs2348eToye5oeFG8naU3gf
asSo77ZZF23Qj2kjPT+5lb7CsI73lhz2MvkgMU0n1b0iogAzn1dqxjcQBXNeF8JK
4ROtkg4egSItPzPu77mmwoJNByi9OcyG6CRtm77hyKXrRtAVoW6ZbPfX5TlrRMaJ
qJfhpF1edlU4uBQTNXJCNlLlT2wgGISafXvv8o/e2hChXM0+oU+WfOqEJRtC/RqJ
bQ5Ul9TSBVe5EIu6+33ndWdltC0jI0/++LcIZU2agp5yhzBxnURcXUv3WGOY4dg5
q3NpIjqRBXUxndtFZcS9oOSDQgUrLao/U1VTJKnpHkOkr+mHq0jU3C+GA2TxtTLd
9viBtPcGb64eSy+Z6rTGq4RdVmqb8soPD9austOaQh1s8arqS+A/2AVSHmFW+VOY
65eBlOhKXwKjUQ5V59C5ZkPHERQA/lvSXykgpeMcdLWv/ej+D5MoP5D18s+IwM8u
rURYNKPaxctEPNO33JnnfyXw9gbsDBS26M7J7vJUNSwPt2FbiVDyWkGhBB8BQn2C
MObbyaXcwz/cG25QGoMBSVVwcUHX3obbOe7HbImYUIPDeXFBRCD2D3YxG6KeLvmB
Vmae3qX+W2yLdG7zpAi1KEmcNEgrC69mDQTq+2QBLa+Nu2abuumZ4pfdls8Pof9B
ad20V/OeqFQYP8G9fCskdMu3WuD85bba5dpUBQVt0BMxA+Ns2TKb+3nS0KXwgmSI
wICd3bN6q4g61HifkSPbayy+KaOS6MfR/qJoaL35Crp6pRWnJY1RgbGPpduQPJXD
I2hFBMq84WKHJDLt+EJiuTj+cErK3brJF/xmvpEmfOf5Uz7POSAr1jwoicNsvP4M
YCtk1a/GXvjKlSyZ/SQN4YsRrA8R/oF35Th+ZOBb71INx9A6LCmhpuMVtAmCRvTY
Hg2XLM2I5fkNLhi8OKpoK1fjtHNEefmob5zVo2GP8caDTBJZZaLzhj9fA9W7y/f1
1aBlv+yqvNjKpTS8j2A6QARFVfJLNO4eq4qtfskMQzYZxDzc1AMiD716wiVecb0L
X/1gUB4qIG/wpCTJaOIx4tDl8vhu4gjESibHC/q5lz0CEllemR4XlB3knSpiMWEE
j/ph61DhGYNjRh/+uSCVHJ6v6vv8H9Pg8nt9gVn3zbTG0a7/4bF0F38mQSLnCZAe
IVmbsltMr1Q4Liggmnbhf6OSJBijkbZ02mncvRl9KArmExrUDdq66gKFY240ciwL
fWelDuH45gyUtGv4/psKaF4Z+c0dGAuL8TbYKVvJvKkdwHotAV4biuTQxOKHF0vh
SmiT9UZeZIG4dbe0z/B5Iulcs2DxsC1z6X3Et3NFzttosdfxywRo2+oLO4DhUZE/
v7HcsCsppQoamYmF7EjP1E4mHuDT5y+jCoKj2z1F0iAFjtqOmF2qZ5d6WT2iE5iY
X76zaRRPpcAS/xqRfyii1t1aZ1kSvQTCzLrttkue3icTwQnBo6DEaj+G+WJiQCgo
PTMh9wADXVeUQbO1bXnCpZacYAwfPQRpRopmVK+jpwfvnZ4MEQ2EWf+f9rtmjiU8
BJQxEEQsZgx+nV/QNGzFIoQ3pBvC/gvHIwIejNHPbb7IWIMj0LNJ0xo3cdzTnMpV
1UXBc5dikYQtpHrJ8l1Ug+y5mU2T9dd2BLwlksa5+kLLPqyof7jz95QmQeyyE6Gc
nrLwDxfAzp7zx5D9RqEmKlRAabH2WdcKyk3lM/dq2hqTl/9Oi4a6aQ2Z2Y5M4FU6
fZB9b3YQNPBRr4+G0nOkkrWRKiVF01SXEuzZGgM9vZhY9CTbBtuD4XScORAWztNy
s5OAXMR46SwWSDGxs0WM8iexHkeWifwOLWV2dkLFZTmVhuUe9fpHJ0hp+ZxPM6mQ
eAgeZ5pOts/xyEfo3dTjRw6Fa38l5WcmnxMNYOBNJGzZCnQu6CiMx/GMC+WDyOV5
0lTCVPPRKzDmFlhJ60JIK6mftdUhqX3ZuEaIC4+N3OP4K02Vt9+U2f68ikMkgEQb
WWzcob7PN1ueawca5OlVqPZjDmmjHGtNf8mkIcQwe2lqE3otGe54UXvWL8lUu9W9
ksPrkX63q9BqqwhK2NIv6xuva5lRnGdcsCRk79a9ixbXqZEWQm9zSSucl12rhL06
LsLiqCqt2Ij+TbdI7PO2sF1uze0f1p9QGJp0lTNBcWhhtBOvygX8lbTfHyHgsk/q
x5dVvfTdWdCzeKtPSENN11K2PeQ23L79xFo0qRm644bFjJ4ohPDdTIe5KJHKAPJw
txws5sYifiRRhVdPdLLxGPognk8bfZmP3MLSlaWIa1ahlwa401XLvCuXCieiNeC5
zYxr6bqGqdc2ieBrqZHQrynIRr++0wBCxvH52SjACsiVQaHTnLyV40TgBtuKVdST
uN3kcsW7PH81a7Cygw5AhdeX1rq3vwK+IgIwOFrzjvbtcY/VUwuaaU3D76AP4sJp
hfH+1gOMzf36xhMXEkTOYL2LsLEblDqvvtpGKSUuzXK5C5Ke9S5T76rHFW2Xj9dk
8Puele+gdtOxQXEEgMOWX0+TqBRE6hruFQ35dIq7tKXYasCxCpCqwuAH97n/X11T
zXtG5BF33DUubtjCs1MXIEmAGfcA5/CIJPnG/YiwqdOck4gdDeww1Dp1tWwuwgXH
/Gkh+dtIQFWpNJq4//JdnX/cX12wvvHykPAimqmnHnuL27iYdhqieJFx3KTBavb1
Zdmlzobv3eQlIbJgA2P6R/L5+2MREWe7zfv4q+WnD8cmq6Oh4i9QPSGRU0kNNqBN
QcMiyZdZARcHRCKIwaT3K+JQ0ngcB1eHNcKAEjiAJhft9T5kVPPq5KvA1UCwYV+x
BVLu/qybzAtV3WbEPcZcmazr/B8TUoe9O5thUBDnCsW5M7lzFXTmuMlfu7ji+SfA
1x+xoIPXiCTAD01snMWLSAHcIUY/filpXHuKMegcqzkZWVUgjtnY/ZJxVUsJ2YIK
gUqulfoBe29nAaRclYBafMw7RET5OUAIFI8pNW5dlRKZb3YFx/5SzUCpgQDNXfdv
wWY2BOFSAxJyNjLhg5Dqvw6JRXZQyY1I/FmaHuM/HWlFereHmqNHPxRCRi9857q8
hcK+oexSKYS69BjD5MfB/sbWJC59kdhHik15v2vf6687M7onB4noREr3i3866oQf
UCS3gGuMkchnGAt4pbO1kA8/Ns4Iza4c8UOXW4AE33Ijw1qAL25J4NT4VGyECRZ8
FpL2L4Bdw/7timkAUGfzf879xUvL1IYauy5uu9UDE1YjvCrQHErND/Q3AE4lSJhV
vB4vJhaYx8HnYxhh6a9NphjiID7gC2J0KJ1MJ2MKSD58R3UQvyPuwRtDf+53G6SN
ydMpRBrGVr7hI1TzSADnQR71hZ8JNS+alX5L/FTjVqpuclmzCUtPEXmeWidVBnXx
7yYCj8t5jvYUXYY5LQTOOnFM2t0e9NUscTO9tK0jEScNwGYQ73cAm2hNLRkviK9E
fifFUVhMC3tKtfs1/idfBHpvB772JBNfEwH9mdvYWqSEEQ9YNZ8aLhYWu401CV/3
/LXj6HMQknGrDG8Gm7C0uP6J8XLFmsV9Itwum+tjxWjl4ubwzBR4HB1uCehOPfZE
vpxprAtOYwcr3ORk5H7jxfw/Sqy3a6d2ctaCVQym8A00MfOJ8gKjJ5llSfZowb/E
bH7wqzH3aU7Lm1KQXDB9LEqFomKvbilfHqz/FLZdPwK8U59RKF+kMRk3Ddo+ePhB
d8wHGm7YjGxRZgmfMiuNXqMHvZw+kW6T751ms1U6oT7isP4PDDFbP8ybzQcQ5uEr
+oksYyDH6DY1vSwC4uAi5MlTVENV44koadT87MAzJaVC97nMIGawku5idnwK1tkO
J2jX8T9ocrLO26r0Q+PA7BGgx7Mol5XfH+OzWGRU+6UHG71QvsBmv0ORHUZ01Daa
fVyEaeov1q4bCqz8M27AUXG9i4/YtQw7fghy/1BpJKsLLRjlqS/1QHP9WgA8jPdF
XvR9HHQIbQUXdD40h3Bptpo6i17P9Agx7eaSqEqVRUDnhxwUeQ8FTgoYHo/Qy5PL
iD/N6RY8PMFh1IopcKH0XcEQwrllVstX/QmuSoPpmecaw6LA8pULvPsUF5DC7vNs
mROjRK4p68Ii8o3jboSsXndeq68GmfWcQiOQAv0cbiN32XiwWmSjLzZ5aVgeA3Ie
A+w6w6xUQS5kgQV6GfOjSmL9XO8oSMZnmL17Eu0z7p12LyGryI7KN6/uacaMtZMG
Xm9hIt7t+IWdmHQQvFeG7sR4YOloEyKdMR1V/Bka2t6r0b+tHR9roSIbU+eMvGLX
eap0tJj7q68siScIhynSAqN8Ly1DuvKQMVciA3RaPb074MRnaXvgH2Mz5+v0gfG9
qq8g1L+IcYdM9o2sfyEq1Wslj2JovQ9rEHsp0JqqjMSg77K6SgLHTpHmkRPB3ZZt
zixGZqohVrN/D5oAF8C02YUz7FbINyZiofhRNp5XIHVOOXqBwZlg5a2jAR9nyKJM
KekU3xYvdMQQCBHrQMRHiZ/3BHqRLZok3SXVnS9NEMqmGR011BlvQN1mPgymVu0e
UyuLxtDGYWqnBSRQJIYXvdR89zfVTk+dlKmBCOD7uVAJ+RW2oGLtrMG+jV4hPKNH
6nSMpQom9SdRRyFgd2YPMBB1kSUDcA1jpjYQvw+UEIDUpW621KQMg7iKqt0X7n4B
DCWjIae4RHS3UROW7lurMY8fSz3Wogm6NtNoE8jr5KRUR82yC+37ZrX7M95WSove
1Rgaf55zVkNUSngCa6mZZUc8NvnyD00SD2eTAVFn9W2BVg3+aBz3AEky0MrLDv+F
fgn5TN/SQSWBpFVrq1ek+R7hHpyHoII20cgev9mCI5zVVkV2Lpll77HC1Zzjh9ee
+Sf3MjFLvmMGE3uRtLedukZP4WjVgFxdxSml6N+VkFYTuSBfRsm87vSVLra8IXxq
c4TTnGARvyNhi9t+eIT9Z0dycOHTyIqg9mNpQwd++PS4vrAWu0NRHAyqCUn0s6wZ
nsbDieG/BscKwpKOyulAB3cxSbnZXf6O65GOWbW+ftd3+rb336XUtBiP+o14WsUI
jwwo5ups3SGEYrp49tHLMyfRnXDTx+bhNrtAiy5zWL5vUnYZD6EMdpdzM7O8rtbt
xmBANlKhls26yF6kD9y5bD3zx4S6MPXbNWDffu76GfbyeltTQYgDvEejHbbCWDKO
19aHlNtcVscx2zWKOEkYNTeRautAqONhD3noFpMQNVgZjK0I1CsFTtpQMor7rvQv
xquOxC82/MhSS1Cxrw+5fEcdVst3QBEMgg9+5s2l3AqE4K0h+P5ea+NHoXAxDZ7x
TUOVllqkAGnO1k4HwU6S4l54hOEITziKBcn6e84VBScEWmituNRWGgwR5s+dvGH2
8+zPopli+q7cgseHnLVOeJMs8KfUOKN7zcy1ru495OujjkMBCwN6atzD9qIC2YCF
PgGcQvBPlNMo9saun0Aq+BhVbepscjqOuVXrFzp0pz0Pr4c1VdKVSHBLRWzM4A9U
HYkS2fGVlYJQj2O+1m0yI3ho/F+4V4cDpgfNLZfRvT2oKkDkGgrRyZDDd1ZnC8Ug
cSCZbZz+PsG48vOJIGBU4fr3OamOcrLSVzE3CGzjsxgLYy5Qb6N5Z4K/HaEJS97d
cfTJHi+VNLGsVbzCFsG9oYgn08zLIvEc5BsYL3xChkiS+iKQsa541e88XOzVke1k
2LUKQormCfMujoNzbOdJ+STQ2MmB1q9K1cS15+9O0w/sk8oMig/KTsC7si6OiSld
jw6EwhmxtMhRmTSe56Ys4ssuTWkOCqbiYqqD58tp356Olz1j6DQvPTf6o0KFvZwS
WXKUxwHUVYUQi9eRZLCNE9bui3rjPEn/stTumNXSMyQuCmUX125J1+VG3NWPZ30h
UzOxqYOIqwjNBX5Qd62Nu2w8oT1lJF+FrCYMlc+uczkUDv81CNXUpaRj20o+T5/X
nPCq2UHrj5xzdMBl9AowHpkb86lOVCwzrsbA2cnWRBXznvTT8Q+W/Eq32p16KHHv
TYI/bE3VJqUeDGi35GWoug5NJbKKGGAc69JfakGJSuUmERzp5HpyBqU9Gf1JOPml
NGgMdb2ijcf+xvC0l/wJ55tXS4e7/H+GiG/XE+BFbxvsHyWvfvoB4SwLLgJzUve+
QLcMGE1bCn0Sn4aB5eZcdHOaIkvDoouRO5IOLEOzHiDFv9Morry7xMLRh3UO0AVS
+DhrwkD0ykEyAkAxdmOSh9raR9PqscooCwRwCa2N2aeXjQQ8rMZVXKXNBNQs9Du1
XTvnWCiCeWpUMUecVmkNEsgHQ39xBCKHWB0NtsNXcPtdhFM5H9HPLdcPIY2BdB2+
V225GAqZlmyRtHGC7jieEZYdb0l0vDIGgjbGAVKPxB2o605PueKYQ/N2J9oNvjJt
Ef1UH6iiEmAMXgkEg70/7VcTHyPway0ty8rDXsehkAKfUelCpz/Giuzg7c/BeuDg
8IZoaru9D+nZ5CTwYtCgNXcDO38IVsL13/NE/4+SNAR17WSQJ3PbLVgIXy0kKi8T
YSAApuW4wFUgf0PzlO/brGalge4cbqDufqlTyII6tUQt9dw52FDJP5E0xnzvWa+z
ldGXwLpCJCRy8jx6gTAYl6H8pfYrLh/PLB33AgwvNAjzlorqm31nbZTc7a6hpYTr
J4zSsoiaennBdMO7p9rEEv/Oi2kYR9ft87d/d0X9A5HrZjQqEvQakYxUplLDsmxo
pGlJszOdkAlo9yjcJtGXes2SEccGravxh55HPZzbJv/YRRjGKvBPVm9I9E03/yHr
/zL43u+GNqGIK7wvbmSo+PPsUR/aI+p5wso+kysSj5TnT4pJNmMw2gtN8vhYVvQr
LFlFR48BR230Z+rG3d/MwzLkeA0HOesrcINWqE/pmZcFFImdsihNRP12OJfpa0c9
RzombkQE0p7W+JC2+J1sFvl3hU2F7PH2OQydyX0ybz/U1L+0T990xy1LjFlWFeOn
9Be1dldI7qkkp50bXi2Vtw7lZPZOKXNoK2pTMAMoZws5nS+VN4SsIALMw41gpa3n
po2UhzhpMehqWTSglJgoQTXYFl3oi1CnkWBbdjJgyH6oood1lZay7uBC1N0WeRBV
tOUi2WF2RhYiHwA+d+1YHbdznrb7XRFRI3h230LLafeWmRTBrqTeS4cr1hNNcZ9q
fhIZid3oO1rLVipqLw/H5eHiw+xcWizmNgvPaXbaZEQkaw05b2SwUpCR1Fh95/3I
373ofDDU4QK/DVCP+50ZUpBNwnBTi7nj+62v71j/G9mULvDHMKKAcfU7QIjrX2ar
vhbtc+dp170hnJE2OTXEQ9UiPkj6M8md8oRojiTdbEpBT1w523ToTv8T2ynVJKVi
6Km87JsuoXGAOAb8ojlPPVJYGWYLOhF6N2xPOBcIP33OmjxY4qC8piBBPzDh71Ic
bplzqHjd+0whgN2R2s1jbg5kcXonMmKGJdYAdkOWeoM+1JkrcEZL2iXcRv9X17fP
/R59AmryxNT/PQmrUt2MZT+09jX2TskuJ5j4Myl4vjcSsBag8XuM59VZtdyIbIL3
ZipoWoHz5KWitphXI+165Z6+nglKiaJYo5y12q9+VeD3wt6PbjN3y8ZXl1IxjdMs
IK+e2NUhnT5rIiZLwBqUcJhMJeTIx3pvdfc2OtksEqZmCJeuXH2qxFREFZezssZe
84InVMKqJc3N7pBiBQIX9H6jsnzNxS8XdDvmqswd1xlLkfoUnHS7P4l/dTxHO0LJ
cg4xxXPEDrpf1+CGsvCC8Bgwi0AC+gRdTHfU5B56AmUJctHAyenYS9Osf2tUgafi
qsUQjk0W0n0eVfIgb0HNoBmcU43LLxu7pKvDj/UPbiXoljSImNUMXTzoJktSKIom
Uvc8geckvVTMEvOgf8OOrXCOQjOS88CjVzqG27+F8jrJZ7lYTIc3ybMTOGDJyctR
N06lAfov5q0TSNRm2YKffPDk9Or/tLAOKe/GRAkv553SdpkPXkCW4LZ/gOq4HkNt
b3ZcG0+BmrR2YCSm0IdVOclgpvv9Ctb9ukhV4445sT1pu5pns3yJ4uVTlnvhPFGo
ojcyxfoHAzOa886wUdO7MtUs7PLg26iOYMx/cpmutoBPboiW8ArE8fOFF35m+0WB
2qlJD25udhrzeViM+c1eypTK2S3vh9mbIf1s8oNs6nt+Bx4rEmFKPSzp0y2a2N3v
nyQrNRywEH0XoiDbI0V8P/rXPlb5GHAfmDpZ/vg2tHFyOhMv5gMMhXAsZTeH+nCm
uZa3kPR9o7hZXxR3kH/h4piUR1BBhEUypkYAbV534o2eyUTK1sM9iJPdEpve8Bzs
DMaLk+cfVwXLKH2DeB1PtjqtO6WTW/42H8Bf2bTfySC2c6N41rJ2Pcp63zmkYCoo
Inm3QiSFb7qAdd4vkCapnuOgEZiShSWVTYAPVEi/yo8pE0Xcau6QKBZCIMrICEcy
wZcbZcsrqNQrPHbnkMUaQvIt7zw8459Y3iKKqZ/BeKpn3heOvjnkMQRhxF/RalTM
K5cLxdPElNr4yFGECBUzMQ4CKBgTo4C0LD4O8E7o5aMFp5huk0JTMwLzkUhd+hjX
VlfpTUA9TAq4PHoMNT2oWof3v2ULD7sZBrCzAA5LLjKKZ9+etALHwWM8Szv1r6xl
hubFBXMl+UJhbJWt83DvopjRCKMLDLQq7I+jx4eIMr6rUqoFWi/k1K9ApL3qFqK+
jIYlkaGf5oQId65XF+HWj15DlZvzqEdSqOAKgj+srGoXJZZNNvgokbeGsFRqBCtK
k2jxH09EN3Ex0oj+GmeISu7bIPeJfolN97A4I440DjWG9Hk0dcoJbCNWq81Za5eh
TQ++PmifvI/p9EXHNEwlqNgWHivmVccuEOR6ILAGOUijb8EpXUUHfyeJ+5Gej+nb
3Eey9Zxi7yT2ODJ1MXfybW+Uquha1LfpX7VohknEzPSozaG/U4TN00FHsvMOc1P+
tEpJ2e4dfWY7SY+KbLFZbGyPeFZZqFQROsJU2BEk8MrdUiVc4f5WrlMibyEWlauQ
ewYt72NqTdfDnBpjPbtjVnN8zvG2asLZ9KNnAYJ7FOuhpGlK2/7BIakfA1635HbW
P9zfrlgfzCH9/yWBI7iipB9k2Z+3WF3rUaf5akNw8NlAq90K54/D5F6Xq0/uvSQ9
jeburPzQXnsAQMw/UFFJv066GfIyfsoXR31NWxCUjQOs9E3+FoTzOSyKDhdt9Q4Q
zOUM27dkhKwOZxcw/myjDfICihUZ5VAEk6pyrL3VATAvPJMHmEkjWxC1GMCtiNhu
6VQizjvZmpf2qgQois65P9U/UL3N2Dkl/cvMQmoTSfq1Qz1IsWOTqPYZGkPuG0c3
kRa5fAsUNi4PSzzpA3N1ANMldhYYQh2XMZa3u8nZEjYGcmwEEFtdM4hho+1GiyG2
9h5XOCpZ4v3pZQaAnRGF6A0/QL1eKScK/iMQHpcCdB9+xunwPZVvJfqpiYRtHX3M
mwzJJGBwVHWacpNg4pFM0JbF5Zjm3nOA1J0TVhpWFEsF5o1EMyinqIGPdNSO2eJX
Bl1BO5PtxMtZwhuMn4V2zYnrDE9rM8k0TMwucPlaO0+Y1dbUCuaeW72Jda2vlzBt
xJqbUagxJCSH5vL+qCZUOkpc4bwwJB9yDtf7XYeXsQ+EF5oUsJ8zKo7z6Dt+SdK/
JnIYrwJoHUuhsZwOMg3w0zZIykVyQEPl2ryyI+NtuLxAz1dWBwsUtC/PcP1Eycpe
RPDPOfNMJonwKV9Ya14gIMSHTTlznMaQZf/xCf9tRP2t4IbEjKfiVQzsdhsu6hZr
ZX45nktf36GevjKl8/A+L5LgSPEkvnfLkr8oas4UP2T01xoU2OzOG/6soNQkV6/s
rERjtqSpGR/YziXsZy8MFRAdjHJhS0B94zqD0bt8TBnLNgn9PQlz2eNPX4hLeaGg
wPFqXS3w01jOLoDhSGj70v1Syhik+TSLnCYw07siMCL55ffYHaZNi2sUZUL1NnmK
4LU3oZyWII+1yJttXecyaSQLU+KCuSt/UilPaTY5Df9hyPdRQjkKVWE+RzRMuadu
RsKqYJuV32z5vN5Dhyhg5mSL3e/VELCBjqauyBzIdD3ugobeL+H1yue//xKayT51
c2SiuRwiVDaj4FQynd910QRLztki3xN6ssaitNTrGVnd6HNOo4ZAlVl5HrGQjeCE
DNPbTKKrtCWLHjCMPWLmQ61TDUAvG3NsxZNMcVrq/YMx4Yjg1WP53hAWYPy55nOg
D8R/c50EWxkVl3dIZnJBh8h197zmllg0WeBgl+16UtXOiLJXlxYER+YEWwUjpOv8
cZfwmHT1nbNEcDXh7TTU5KWkmean3hUCu8T+GY0b3FC6AZTPkFpibc0dzKtSlmtm
4IrL5zfRR7dSQiuo2yhft5qUxyuiiOg9inA9hHBpSSkLgCaGsCYrsrJs9lVrs5nK
sQgOrtZrszwSA5WUj11VG8PjPo1u0Y3JfC6G52Kd+czw3hXRN4lpSh+aLTmimKcX
/BSG/rgbL+4NcBkpNRpQljPOV4OsWNMwIxQ/E87pvCbon0UKZn61zHHhMlwGPd9d
pCcVO6w7rbER+ejofcAaCBKhq+NBl+aCrshNOp5gv4S9Xuf/XTXNPEnGQMr9NbJR
dfx62WouyO5o+L7Hkq0YZ1v5gMU3SmRKfGR9x03A0ZcQrz2pdfUB0f0xqrkxp9R6
tlCGIcv9DIlvUO3jJvmgfrXDtKdtzJCshur5PEW0HizKlVpB39ecEKmC1IyzFzYc
kpms3z7kN65XmKaILOuHmT5HuyTv0clswi884CwjrA7usohv0Juyx4TL3qqsUyS9
DivvDNyhsNRy3udYigAP25EpQF88rMbBwe52YqbbFOw9NnX7VDU/i3BBWRl7a7ce
0QzIaWX4NdgMHFZPNoJHwWcsV8NwLV8F9cYFfN8LeZpiXyGCP+ay4Z24CdkuXa+r
uGed0EoEwnkKFKzQU4j+Jv0ag/ZpLOheG1j2vVsj9Zf6sySA943Qg1w4VAZTqYKb
2F4egBE6MdD3WdsuKOgcepPhua/aVFeNLYA8svLEr/nmzycwY7WXdAxeOAv5NnpW
DiAB3p0e4YR6zHzsKRBRRk+lvlSUTKF996HZQy3Lgc5mDx4mt5st6HP8ZpKPfcRo
zdoSZuGFIdWth/0NTmoLBaWogn1FrHjlbDlp6E1y9NPdLbULKmo8Bo+/M6f7IVOz
MfisxVgHaF4qM8j+JtMbHlkDq9YYYtKaMsF71Nk897MlBArfaPuqP7t40vxl86bR
9BfHedHX2faZRJ5u22MLjqShxqKTXaPkehPxVIVFa80e5CAm+kzGLc/Gp7yM1JHI
7NMDBsAkVvIHTyGGeoZzpiHK2bJiynHQMmXzLnVI+Fv9DSpqjvdAgoEQAroCq663
D92ZD/iu/PkKfONC/JSW4MhjBcUYUpBBtnJGgODUxAUfflNWxwK8XYlJ8s8QLpOT
U/YDpnntsdd4DpP/uLLVcqXSDixAau3GY36QEOA5Tp4MkboicW7Uva2ZfUWKhepl
AvbiZdb5VAtgSQvy78xiWsngiwiFrWg8Ynag1MjIKf8zu9x4w3HTucsW3QJuLtIw
BPh+8gb3X1G6SmW7D0edhT6oOsoIxlLnpOuW37lP+fI+5J38TVGIie6l3YH4d5th
LJUy5Bdtr9rSAyyMpR/5VLW/+2V0D1ZguwILT18AIuTMB/46+G4av7d+uJysGYBb
KDQLSNsu404BpQ3Q/z7ppe4v2kJlDNB9YGLktq1zejSBKGQiPLE0JkMWGONcB2MS
jeJFV2QvemVmNYyonPFiRyKnnbzdEXWPGMemVJL4Ql952ZSRc23tdv6XqxkCLbti
uAs4KzhpapsHFRb95oatOli9Fg+Pu+z2LoYxggijgZsyHvDPZ15DIpVqlZlyrScs
nEKabNJsBsR6BBzlM4AW9yvIiqzvifB1EeOC8sj/iCvC2Blkdn6tda7gOogoFRIE
CUg7gW+Xi02HqLrd74hZMm3s3nAHwXPb9FPz+2yh3469PF519nZcr7jQ0kB/GawG
zWPoSNKUUYwMaMw9r41lgco96W/NfBfjIjHRi9HaeEo8NcDA1yPA0Xa1BNfpH5XT
86oYzbqjrGtWJfjRlSTLgL0xtsVgndPcbKeSA4KQ/vLDdqwTXV8nj/HY4rc/4PLJ
iwW1bwIoEqEAiou4lqpoMsFRRvyQEU39X0IVs8DLPse4SxE5MgrZ7YH8O74snoZl
yirTnPqnMebhHEhB87j8Qb4FZMPYT25wpf5JIgXBLU0WsoAV/zcP7Cn9o2ex2dHo
sKaSdxFokAkvGX25vkuTg11MqFbjiziLFD5YjYUh8duVvCYVCt1urd+jJSM/caZq
C9K35u7ErkPu7rH2Fe2oJt2tB39eK3EWG5cd3x9zgAlgh40bA76IPlqh/R8pK2S9
Kf5LathgH2fG605450LpLDZfCzs7eVcn9vLqNqpBZTOXDFydZT+XlAQbRCMC/hU/
Psrsjy7vho3TvMJV2oF6y7UJL7XjqOmNBqhB5E3cD/KD2SgccoFVTAyeF/IaN299
em62RtZ49SnoqEACeisq1rsia0TRNQ1V9TN94RhrQSTcAw5hKKXIS78hIm/mBqxp
bg+DcPFoB0KOtv7B/M9ly5oCpRO48gfcDxhF2LvWI33FBc4LVLPf2JxVlzLHD6xV
WnEaWTJDTBU/G6D4VMivplIMtRMQk5y/AdA794cEyecTbBLEt30M1DIFgXl4yT/q
nT0uGKIyitif4T5USJLQMSq1tot9PNm/5tRp27qzJKUl/t75jMixgktGByDb8EB/
JIDcGYX84/VWbFOVa1fNqdmLocuL9Kk3FiC3dn0mERuZs1+4uuWfBzTh65+69+Ki
53biH9RKQ5i3Vfc+gf8Tm4oHizoqIfD5n/XFyXnvvy9ZaYet3NvjDriWfuZ61KjO
dwNlvFH3Olc5b3mwrpvIAiUTb62127dJ2k8qcIypxrYG3aQEn/ZY/YnzOPAC1Cs3
EMy1usqcRc1+YCcpOtgPiVvyQxvk0Cz5H+lwcPkSm5m1Rk9kMYz0CjKsEThctjEr
ZhYkoUzSD2Hv/WC++NslYbDvXVfkh0EE76IytVNn50RIV7g87XX1xIdoTiCZ9pHN
CpLiT/NTGueSJmEQUAeuS+59efJXci/7/ec0WQ+rl3q7w5zlyiQD09t7SJSsqz5I
leMivGCF5XxFIEjBVoZ8jrQbGrgepCRn5y/jCqgIXrqzzNvlmJmmikj3A+jj71ch
6ASuakwYYXjg3GrxKpKpujkN4QkVruQt0ieUrib4O6A0ZNiOvFjLlTnpJIsOOpTt
JkzbgLkDlh/AQAlv25vbXuMWEvZnBRbyIJIetNM25uii5t+MS8Cy8bFzWqAxOyQ4
3gDmN5wqKeGmBtCQ2ogQzgR+GEtNsAKZNHwYeAjJ8FLFLDBV9U6Yw/4MVegs9CXG
0vXUu/Fatv68TihOi4h1Hzsc3sVRfcJHY7Du9OAJwRBq+6T2qg2piUI3m5BD8it4
TOQdFCFxjPTDMra0VuNUqmDJ9MzACccJL02HrzeHuX0H3B2gK0PX+XHPbjtVNbUV
rNdnbEPD47iwkdeGXQldozq+mQM3DUFE511m72YEaPz59y+ya7dMf/vg+D4uGWyt
5/pVrCdn+5UBSLd/66sAcRoFPNUWfSJCkOsiC0MXacsSN4ln0zrL+WiPzeSd1WeG
uu8Yi9qpbA+pYKWpcwZkzBGY2S0SPP6WqDWrT+zX1kBLc9bwjCpyEtBWBbgF2f1u
DH5OraWC9Q08s4AX388BFPEn1A/uDV/2S8A6kk8D8hUmuBvlZEVUZbuYCthYk/IV
KSTVIyMSq8xybCUlqr1Q4GzpiWpiVRXawkezJ0IfTRGTIlwpqE01bgyXxIfGkQyZ
bJ1uOpxpyW4CBDQ34v+8+I5ofJ6l9PSrHUPdND8H3L4TfAWglYeWYxDhj8HyXi+Z
hiszCTE3xPOQmSfgO3F7/tPq+Ty38KyIZTvIaoDq/t8YjBzNb1+mOZWCwgeukjx/
q+8hA5id8zkd1nmbVmrnrevOagBjBLlncTh951vhRZ3/Bv/qFKVrosZ16crIxXCD
+WZ5LyUfr3yoJ2hYjDLjcoJu3bg162tdUeHpyKpLhPMZYy2YAzdZx4p8Rrv0S28B
T0hMLPAlFPFYLZRHhO9aYDgfJvHMm6TTH9WrhvuBsMaZUWvbbxvFv1bTQbN9i2s9
Hf98JKF8sK5gugfuZnzD7s9mKuhTanh88pxgteBUxZQMORSuSpqmqb53P/h8M0RF
9kxhopUE/GUQk6AZ2/Ars557e/sfs+drimXkhYMSn6nxaoO4/3YigPWOQPmykq83
g8s/cefUESC+Bztxi16znE/+HSmw2GmnTwmq0Hwr+CreCVfkJII9wemU2JjnfwEc
9KOnYmXsCIQpKmUSSUgRsYmT5Tx9pS0k+xQoYEg2s8qZSrqSUtYkzibObgOoLRv2
oTXjVRVu6GpoxqrAmRTLjB2wJo+juitUXECuEFCKR2lCizXS9ZFq6aySU+R2o7ED
Y6lHfmynlcz5GkRp5W28RF22fs0X/flKug+/d4Se71Dey7X7F5Df3hAVLFSWHCbv
0Lzpgs4RrBV+oXMF36YEAkvzmDrwOVCWfiLpXXK40owhekwsTo2HGbjX5yqXt1D6
Ac/HbcvmiJi45ZVcmIe2A4zYCvz3KQ4luoxQ1h9txM9l8jDick2GkQWf/iudL2S3
XrpCukn9gyKYG631v5mxIXdHdwe3PHKXPuH/8WDPJAeGwAPLi6x2KRaXqxnz/h3G
KSUSV9nAejpnz9ipEEiM3IEK74Wk+jt5MHMEgD2jZUzZ6+4CBA0mWy3vSOLAGj6E
A4xzn4yoF6m+OdnxBnwft/9t4zbsm+rXFrlRcqVC24nq21S3EbxraxDYV/+AidPF
3sLzCKLQ71F3G8ZuaOm5tsUm6Tu3IzmqHNqtORu1A8GLKXlsoKaN7nfBT5HGVFQB
26d440FsONyngiZV/JQ6T20LPtRDU3ld/kmN2Rjtx1wnnhIO+8HV3lxYZwkDzymU
JgeE6Y721sWjyI84cSSEkhwWeEPLQSMKO2d5lmum6yvcGRFcUxPQObcKL4aoPt2C
NZRoDqVsZEiEbBySqIRrerVQnaQ1qy9xR79rvT3fSfWFwA7krC2NXZs3Gv/3x5yd
yslsQTOW/xZpuari1fmNpebxloofQqMT25PXXwvO0NCS2CTIgV1JnffGXSDFgW34
uGnv39LG48Ffi9Id2VZT/Rtyd75goqPhG4BYgNII3E9qFhR+SsOrKdJBhPIdXH6e
83EBjlO+z82/qD3jVMjboHEBIaffAKErtts11HW6s5ia/Dex/Vtn7UEdVpZPEw+t
1UFcoNJVbsjdz8+RGx6ryfnJC8y3LeQoYrqt5r4KlUSTOJ3ZU8TCPzedb3ap8XSw
xV67n1F2dd6cmVqKEVurx8AtO/g0TpSbgBhaRSXWBMK98aSuA2GxMuTqrClj9Mx/
OMzHZ+s82Y0yfEOWhI2OPePyCtDYzMT/rZjlsCyB+9pnqL9l1TV64+q9lvGfatmR
uSdJOjXJ5enahcRIZIzUBGAhl7uV22r3cOHtq2BhZyoi4k9YAQQCk62MNp+XqURl
HnTGmSZFgXoBVwMXTZIdk2DOnp5MVyWrzHAZeUm72W8kkj2zF+EwlTgbceF/9YjR
MrdrrLiVLq6N2ZYBMO/y1zEzZibMVHe/kHT73saRBBXrHdoc0SSXyyiD/G7LKrEP
N8L5keB43KteQSzAX/2lNMZLlqmlieT04iyk+wOwhEtz6veXw2OIgGmk5FvTVdhy
mKqppjDj8611kLWZzB0HKE7xSTHGRQVbW9AtV8/gF9QJUSmNf8a1NAtnT7yd9kzp
ozQVwWKlkY20V42wKgG5p8jtNpfUbSX3Ud9cwVa5peEcl/72rso5bbJB1PQv6y/6
P8peIhnBaUiTF3jEy9AR8qAoRur8UQ8TVMLqanATIOyHZFFy32L26gYS94nFCfCN
kUzcR/2XnEkczAWmmS2Zfh5sLWVYGDRRk2xILMpL2ddVewYyAjC6eM8Y+fGd6Qd/
o3JRCV71Opa5s7wrhb+rwlLmeRw80TOlmReNLtbKv92jLizP9f+eJnPNMyl8rqfS
rCnoQoRgbdlfDdVpYpoNDdNGn9rI4Ur+QIlJ+GctnaXIjAsbvV2VjlGP7GsIou5H
dekCbKUOn40bou6Fv3oDNMcRgkK1L9pcj5El/cvb0J+iTsiuvyqtwn3j+olvvyMn
47vyUANJQo7Mx8Icrk0RRbQG15d2M6Jmx8RCfCfMP38LJ/7b9rvpjCqeiijURuCX
MVoT7g3lFcnuHF0y+5JaK9Xetmp4fHK8IlZ5s9oQwxE3KmvxsQh3gpEYLth1noWL
AaMgyj5NCCz4tU4NfgD7YxPejPM29lV/vMrZeBayvCLsU2QYtktgNINVtKkIliAm
aZMrvjUz7KlA1N2eTm0SwA0V5rrM8NOui7BPn0gIhHa7dspiLSZ4Re9WtKnkMmUN
uxqWktFM6ix2KCLAYayPY1aZJqcX8cw9irjfRJlwZ1JoorPoCaACFg5B6im0wPFC
dVGbtwgX8wphuLdgKKJxJjbfDMjff+pVKazmrHPIBz58o3bYoo6mz/cM0hd3Ade2
fgs9uqXwlwzoZ2X9LyB2QzH/SqrJ+n8IISLCfHnOX80sFXbQElrEXWXPBZ55+mvP
ctAoXVINvPZE91gL7ypKrPxXfC9kXCkIR4VJVsSZJO+xTY9FBwoQ91D4iA5fse1r
1qla4oHFXA/6p4+VuwfMpS55F19nTi3EjYUqHd55TWfrA2yQs0+1zpOQBVBVfasp
EvLa3sWnRKXOMZSOteyqEy7CvEOJSp5dlePYaxaL/gPKjLHohdkdP7/j7O35qvQt
NqjFmWA2FdeAu03d0rVvNYtDyC8Y8XKYXX5dYB2l9leHy4woxRmtH+yHv8SF5To9
lPcrb2tS51/lyyYClAK7ipEOpzNxZqNO86z+Ij7mjTEPMhg6cppZx/iny+PYbg8z
3LjSq5l6MdDyg60VV8OZ7jvRFkSQ12J2ARIbXa/xHQy/5Bi9fClBMdcCdTp7mm4v
+FJAP/T+CxMQq8OVR6k4sY762OWj/66mE+IbR9JWg3S/MSHWFCzXQ/wJag/SuMPp
8Wj6H/NKbHlmBaf5MnQHBC2zlEzHFyO1rnMNjbCKbe7C0A0h2FAUCKFS5Wa7OIxN
Tg4ZF9fUq/6uq7+Q+BtFcwoKuLZeDyHM1FfOD3GAcp6BmsN/yHMzP2Js6KOaLcUo
H+jMvp2MlS1aL7ASGFzU8zoc1TIjlU5aORoJ5xr8s5+wdACpr2kLfWrxCUc18Gx/
T+ojJxSjxytWrXR97sAFHth29Lq6AQXgW18ZFnSuEmhs/IUEuZ86jgGjzYoBAC/4
IGO94GPFRT1XdC/caqJuD+wAA1UJoTK8W0BpofVe6VdlU3nTmEBTU5yN51Ss8Wo2
XRyZnK/Zi75FAkatO0qbOjaxU8f7jPQwWm8O2pfRVeWSztKa+x1EwQphaWEgmnCD
7TqovCaQWLerwCG7ZCSGsnwti1DZah2Ps9HkHwqq2Hgj6na98na6F0vO/7gXb32D
CKTAYRo1yZ/iy0NPMoTZLyXNIIUjQWKrJnh1nsST4jUum8Zlv93P0VdRHk7gOXVX
IUJe22I5ZsL20Cqu5iNQr46i9fmCyDSRmi6NjPcO7xliy1FlPN6pdIj+N3wBcBD8
qUtyF7xWtKSYfdzVsJ4YbiIF3C+V+pfB7yn+HMB1mB7P3aV18WJzoIg2Vkt1FxH8
YpZuYFAnvkDSzL4dCJUrbq0IJx5MLzfoF+v1IaT2u4GjyvhYcfKX1LgdyW6VPFQG
Fiu83oL9KPrmTR7LD9oy3WeroQQogCuyT0zmVTeiFyDdSMP9W3FQAavqEjuLfgXr
FFaMOp0KFQjABYw0TOY9k7Kd0JZgJhm2J6OfNSlHpWoGVwwAR/yV/ZS46FCovHG3
bobTZCgyn3Zb4AZ7XzmapiVPBiYT7DRnRpi3Z31bhitTREjQsy5Pm29rhWDUHOaj
RkRVoQUk1NodDNj4qY1cxtERPyn/4YMxytUzLI9GtQfuq2MXe4wFclF/Rh3bxPxd
z0Udr6yRJa0Sp6CW1tzv6AEaJbWdCnX8Rd1kMWEKuFJQ3K7WSREW81VW9HcQwj1u
pI13+LjibyhCsC3Gc4zk+hXP8ZIz9y08GeK6VTzhcO9aAB5cMUWn8DdZmDbRu36v
bekh6LdAHcn+zqWgQhMysZrE12PY2gpoIlmP0nJMHHl0lxN1UOpi+mZzHvDt5HU/
1FPIdFqTPUJ7m0iumiz+9oq+U1x0CNyvYIzFnY+sJplgdRl5qak12GmUZlenomlF
ztmhZIYEkXRaI+rWa0dzHWgGfiDPK8k4dgAabLc2Kg0CiHfIps5yeX8Jk0rOifTo
q/63eDYYiGd6mxuSMwxwzb+47LBldhOtcjvetCcHEdAjUo7nDxwDVitaf7M5RCvx
wYVJGnljnC7EOBp0Uc2hOvWX9/K6f5FPzZjzQVoQdiQgB9QfeD8uPJTAhFmWeKoZ
6kRT6EwKy56TkcM/Nck6yDToduS6uwRTgpwoYfz/Klvdd1ZNHUZ6LaSaW9+fKsRw
O2LOBi8Ol0AFa/+xx4ufYE0NSUYnSs6K0wyhTkfQrXBmqkVJqJrCO+35cVd4yTDS
sKLMxcOeiNXhknz1ujoJzQbvDVzrq5dS6ICKmg5zJ8h4tIItYftFDRnV0Fr0G34y
/cTdiQH1n0J0S1/dd/awz0A4heZa1x4/glTd3QfdwT4yqkLC1UolAGjFbUhQ25eD
Z1I1UIJMzcSbWk3j+S3iS2ae+VXQrx5tHPA15y8rAIV1gSUtVUoVB8VVK5ZyCQlo
8e8an4w31RZbyHwEl0jBJ669gJNAdvWJDV+qLtzZdB0zIicb2hO8nBJGl11kbax6
OGmTWXnrXcVIgXzJfI6iq8NYdN3/4spd3nFN1IFtysESPQKWQ+5fNmIcmW7os4nh
h8WEiAkF7MF7U4gU1aaAjP9m+T+hnK7Q7UE6SJsGFtoJY0amRHlTw19ISdPC1f2U
D7TUYRtNZVU2JJNtarA4zr9O9ga6y19k1yFG/uMllZpLz8R+yJEz92JvaSu/+gx6
ZFVDi5bywMq0DS4YBKm2P33hefXPHV2ZNYU5+iEFzhJrg7vVB4XKsojcIMY/I/Dr
whcikedSOO1Mjln3vql0oF8cu2nzi+Quve429weZkaFRD+nfh1iqmijIuvAZ1Pib
Cnp2lkheMhVgJ9E6GZlPO3V9aFd1efD2qk5rcdgtGowi2JofBcf9/S86Z4WgQbAS
vw2+WJP8IFzUIb8+hQjfEFq4tM9Spb3DkapJjuWNOf8MQaN63uwk5pveB88nyKw2
nhxeLDOISJrupxYfhyaaX8rsxqMnuqlOTiT+8dZTvbU09zYgiaiRsomffejC0pEH
VLxbft6VCcOaQJDliDPviBxMXtHKmAlFPoyXSaxponalqBfCGWdaUnmFEqAtFN3O
8gtb/LDAsv1+hNuIxB66HE0cfm4jJA+CNCQfmLu2PfYOIXe8/hUQ31Fq1cfRoqYq
xG0KYjW5NEXWc2Xj/utN5s3aq2s32FppF74qQQkxREHranJoJQnfgNViwwG8dMlQ
TN5i3m2jbIduuVl2zoUhsfY94gYIbuCBBUsPjXl8I3ahBc0QIh48dst62OmEFLLJ
zspkGGE5qHExEpjCgFyDvr3m29boPmga93kh8CZUbxdvm/elplb23U0EzYqJCahi
OXYC8HOJM3AvAZL2R3Fn5KXzsq6GQDYWm7XQ43RXI4ZK70Mzqe29j1kVda3aCFgI
mOCBiWbMxDuQkDE0mCZRZVGwm7epaumijnQwUjIMeU9rfJHIgadOPo1Sb2hGwXkk
i/O4QNu1B5K+k/aUB8BHcLhuRadaI6dw/axAwCVAUU/NlFsoPbcvBvZOOlcnUvHb
cIEpMKTQDYWa3pJzOL6wRXWmO6k1CBIxqpZqd0SLOsf5KRgh+Xx2Kz7aMBOWhav3
P8YUGdZY+id3iSToPOmb3UOK6HwyYzqK+9UsmsbFxa+nfTUS4CDaS0mcTHLktEpX
bMGeXd7Y93qGYqGkw9DZXoTCc3nL9jcCmqynYQ28LSkt3XSY38fPtdctRLY+Yp5A
KiDyIgaVFo4t3mUIW13S8Mdq498Rh8UXlUy47apexZJ8YvLeMPWC7CadhVEPMEFl
A/KIBbHqkdLWCU2Ic/xRr0D6Mpv6s9FX81KOaDUy5FahgpBpy6kqUwWeYyLTklYf
c8SSXeeSMm/56hjjhptLMasLdAQBTeap28XvIHFljW9uDqDxepNV9ewMmEOk+d7g
q2lT0HGSNld5garIkrii6LuY+buMdTJ20pkJ1jQ9ZOKDBjqiwPDhyk76h9e2fUi0
SW/Ash9+cB3cbmvE9mNaviQdJeRdFOkAyErI8+j0fUyRP64gakaTmB2vHVDoFuu9
xZggul5QnDtP9RybXFPQO3pEJqiMgfoRtvwlI14AyDBJXTVbVavdGQ2NMbcbsZSJ
+JuTf2NpQmeVzlsP2sdYCFAlQ6dem22Qm9YRxN+3x2ip0y+d/xs9MdciwSRF5zmM
9e77j2lX3VyJF6Q7yDrtlwJDFCPLfjqtWPAV/Qn5yn4UaRBLThGcmbLyF06/9Bwj
rEHqtyCRvWcgSvnUIAQtXnb2+tj4SXbQAJUEOnILqaMC4jgtUhFMgX/ffYy1ffQc
75gEkjS5IySUUAZDj9yWxNWyFSj52Q0Mv4IL+nretoeFpaJY6/oO9UQv7+cPv3A6
mBZ0Vk1srhW6W9fCXprxEStzgSCpXsbQzYXIcWumxks5B3cz6x9mz5bFDMpwjZ1u
Q1UY+HzCx8BgB4S4ThM5uDIJ/+d5wp0AsmJ4wR7MQZs9pYuh5mHiPl4+grjpZwyE
auHz4YTLJ+Tyk+76mt4EeKm1k9OV/DVkvYQ2ZCUmXU52HCRlF4QZ/H12sXHa5TzZ
2Npa0u64ajGEu3G6brTIbIHy49lxKAEQqU4kDAU/T0xNCEvrU97hkD/3z9mbu+ul
ieYnbarpGM8fGb8NRTd35YYxcRZtyl4vcxKHp/ixUGz6BsF12xNB2kgPRXpgZZZG
v5SD2Bevp90+YBy6k8lSUGgrobiL0v4MlLJTzzQy7iHH/u1uY7CAw1Rw19rC6a6y
Gp4/n6B7/RG/pVg048tkRdLtVPchEWWF+Vpr+w+JtmHtSpwrxxx/BzKmaouOp5lY
fxW2HBcWDwq83bPIpCbbSN86S+HEH5DwYRzaVAk3YQWgM9r79xyOvHznJLMqevpi
0Tvqewccj6VB3QcPWyps6PX5lhTOnJloaGRPglHaFGB3GZKcPNYQSJveY8lrHhaM
9cF4rOI6DNRs5d0fOJ851hRGTk8HtVMiBJFr5Yzg+3w6khle2en4DUxbaYhQgR/o
BD2Flj0ITH6JzhUIty+wsZBpgBhkRIbTA8pCEjbrRXFhJIFRubgSstB27BjPWGse
lUION9fHm5qv7W2sCGs6xd6Vhb0j9eQ8gvPd2pJBx+2kfxkFHwoiym0DonKZxD2F
BPTho4TWotIlo/09UBlEMbBMYXlNXK31bP6Y7sHtFN241D1WOJ3NYhf1zqUAGQ4o
fbIbTn/IpgedO3METfxEIuDXzSWV5LYAw2I8xcL4UNkdIFYu/xtd+1v2+x+xmaxz
SqWISzj50Ua/wHL5coE6ArFZpWFOinoGFPkyztNGEb6klyIEAWqFwIiWM1d1G/ws
JbruKG6MgFBUrBzQBH31V9GvKw+irLbrsRL6ClLRsFkZ9W0F6Uea/PNyAc/twHql
uHzhIeGVG8/y7pQ1HBIyhuW/LTXkm406+xKlmy+MMePwjTPr/fAbPj9tZNYIC1cV
qV0mTCsYF3y7brXM5dReilYkZV9Ii8HpN2k7f51/0PXCkB5pTsAZFuuSTr1ODc2A
/OOatZGaZQ4uFg6UFqc5cDnxku+uAAKQaQp8NJDMBPVbwzO5fXaT1+95tadkkbRF
PD7Z+Zcmvv60d/rTbr4YV7TqbO/tah9QY4uWfkaRp4NBsrExSC22Ubzwxux7Gehb
PCvUIAvkhl4/o+d8ud+GKsjP3mNIhDvgCm98lXbrWWx0WWi4StEaMLG5q+b3t0Go
4IKpU6lwhC6CDtkINzJ3pnx8dggmzL04Uqb3B8jop/3mMYSSIP5qvEYCzEPYLkhd
B1ikcFk3Cg5mE9BfELuWTZ7Bis6K2+pX6R4mB8fFGEwcY2Ip/6UXL1SXtN8u3wF0
aLqOeSLEhUfBz6Gfnk7RcY67T7qeg1zlu2gyr3+/9KN+5Gt8syeieFPCgAQnSK2j
cyBD9r1NDToNJChhNazvAFXF/8jEnEiKd3LdMZJA9gEwWOb2g0yz8czK2+umYg8z
fdkFa1WAq/YOGgwpcHgGGYTnzmu4gr7ywDz8BNJLfiJpOFgcD4EJxeUk1SKou6GD
JNLtmSKGbYGtDXBzgFzbUH8NZuzH57rQCwqzCqUS6ZjMu4i+UiQ/HkgpRZdEErkN
ayIOR8bHJeLfU/w0SCyfsUqHQFbdkgPZDaBws9VVYOejSOLDQZOMkJhP5pLUkmuG
Mz8w7FQx8JG0EnRIrqXScvJ8fvH5i+CaQ/Sd8LQLMyCPSgwtRGcw3OatSg/0Q9k8
6mc32Pkidi16j/DAABGxMvuenckFwNcQRwbsxmv6TeL1yK/Q9Fm8nzRMKpauHmZR
l0CEKD2lkbwr+pU0cz4C7YKbnC+6f42FAY1RaJ7lUm5MH+oKbh2jJwq4iDt9SIZ2
zWkzLRxOAO7a9gy5qiPzqc8xV+yFVqXtzZ+PPAVVaReKe4qqrc3pDPGE5+g5ng4n
34GI+uwH5zOvsWBgZALsTTFL76lz9h944oNQeMlI/CyJyy7ryaqIUxelHqzoYKa+
As9nWxQkkmHM/29hM1qdqG9QQhv07JlcXt34Cz2ga8EnRCRQrU4+1mF+lMnUoGA3
+Oi4UAgNqEOEiPae3/RTlfxbt7HO1TNhxJDxtMZuG+qsnzGFSYsfbTMGB7/+M5V/
pGsCl7wdSQXkkK86sZn0Q36eEwPApg0bE+OMQJUPQJnv8ptAv6cZuC3zDkIdtWq6
VgyIcAnPA257VD/fx2ALIlb/GNP0tisPAwFehlhQnY+Bfsq6JimVc836rW8wlvId
76Ny1/gy1shmyZpso7uv+yZnPiHXIS888IEKdZJECZqISHRCcEV0RPUjhTRZqovw
svyvu2AQODDu+gnBn25TYxTyvn0KtxLOfUxH+YAzzvvaTtpVvoegMIHP3ZRaVwhB
m6SV8FkqzJ57XHGnh9o7llio3/G5rAOXMJdNk4HR9K2eeSkvgkfBERPemZJs+Mcz
+nf+nSdzkKrXRwSX6dvl+C8uUW4DVzgaufk3CHfuJeqCCG2436ECzVNHtHFmYLwx
uSdVPGox/eEubfOdjjnzmajuesCxVjksL8rsJTjgo8K7J9yVpf68bIBtBm6FRZuS
R1WkpqjJTKpT4jsHIbrcyP+nNynX3QNPQ5nHSyTbLggW2bFQkjR+Vu9H5zJYHQvj
oojRwXMrakXxvWk8WzW+5r4wtygzEhIlWTfXmi4iSMPVo1vS3QCK4q1naYz0B24n
mb7Ir36Y3G8ag4/N2iahp5Ny62QL2qsPZO1VmMCB8i58ePZ26SUDp5sM/J2w9qSI
eMz77U7KdurXmr+ExzVlbPtalGSdGR+1y03Ot1BcwhwoSzvqzYFUomYm/0JcYvVt
E9b6fEkiXOgbirk2rbCVfsj721O5r24+kSyyc2D29jp+KHGdWt5ppq1HEWAYdGsj
aoGryT2T27DIhE7YPAJh979i8yK5/5GvZMmVQXfawLf9hzLdxGnwd8CMPz/2Vu/L
TAF4m4vP4N+AkmhGud6nMLyiQYgzm2wPIJ17HQ4K5IvzRUFX2lAvmNxwIBarFsf8
yG9VlwV0v0ps/OugIJKGUzSoLfFsWrKE65b1suXbq6UgLMONcv0GBt6+FqZTsLl3
9ABjNJPWkpDEfHP+kzgvG7bdoFxQs78ZoZ87SKqTOlwmmxW1zAGV/pg0qhCbeRim
/pXyCYn+7sSx/sLbIn+nlKG72PGZpJLEL9aTe+g9lBz4QrSwrJeamarUIm6ipzzj
O63UQlvEYzpXbG04NQuCiJG+xNOamPNgINVe+xXxiVBFjpooQ0u1liv9Oc+PAIEv
W31iAXRfP6KyAnVbHCThbzOz4rlIvlCrXfNoO+ORCzOIdOskgbERah/c8Kw86P1f
ppwe+epNfJCunERneLykJMizkh/DVlgqRJol1/+TonZgDpUEdWbqekxw9qyeKRAf
tD4gg14MeN+Eghrr/sLJg8BxqfzngRjyzTfa9B6QZ3TJIFbjwSJsvyMfElsEi9zu
f7cr14Pb8aYcNAMSFOcQgSoz8qJ8cLckD5Nd5/jNqzHXv/nzpDopb+Xs2i2mPP4e
8vbBlNNI/EZTgavM2mulDo+0PKvDHUvgzeEOHnry5neUDPQtYWScQleWc1icpSOz
0iKxiQmjHWBGzEO+W3/HMYHdOFzQGjdIQr7v71bibl/iu9q0P3RjHsubflje+Hrq
oywRSAN2LF6OYx7/lX1IdHPmz1HPgioUMG1ltevanYyqIW4N/pjU+dFiuwqVzy6k
E0ULv3T7ZVNdwVUcg7yXKV8+vll/brVWI/BWvgZ2fLlbM5YIHGHLHkOqN7UeWY5G
2L9GqPHVlw4Au4XkVUn51DE4zfqgAGhGKj71voHx6HS/2MGZEGOpquU5sJ5mmXD0
ZrgqwattIyDXczJYZXhv/CaygE43lFOqAQnF3F4UbsjQ0nOc6KlFepVGID+tH/7F
iWadq5/1Y41HBD7/GgBmXlkZrlK5Sc2kc8zFPiNHbg/j4z7wbhAS5t5kkBokVNSU
2dRjkin02hRj45BFdgrx3XHjSABCWib2LxVeDvwWtF/d/KSQCahZChV8Q3HLTEhk
GKcas8fho4Od/Mgkgt8UV1fSlcATvndOLzl1jR1kQhGoL3rgHVVh84vTfP8mwNh9
LwowoS1W8NMxIi6pjfciaQTgp1zVEQjjGNJx2nYhvfVf4q/sHNe2iifuMV/JDu0u
uGSTJKOk4cjHmi17WFkfWcNQ8sPGUxdIct3KEjTHHt44QcOnvindQsxwCrMo0Apk
Xadlbku+AmPGbG1igiU35bs/LpVsfwpxwLQhB7pMrPgjhzKuhWmf+uAqC02p8nqu
7+ra4HWZluclHTHBbo0m1nZY7HUGh+RlvQJINcjv6NK8gFvlNbsi2YaJNV8UjNa7
br8qCg4ONgbC5SRX2czVN01z6uWH3RQutt9DXVcq2SsdDv8MeHNtOMk/SQVQCGtK
ALyfG8Mnwd/+1+S8O3wGWivQYA5BFCX4vYa7KiYaGYPMa+1nA5PYmgg3/bV+AH6j
2PF3XiSXKlt7nkId5ZGS5LRXu1fjlTMXISeaNuVpuLPxF36TS3Yy/GR26bjD3gqT
T3lbuJ9gPsqsXjvVPfqwKyQZi9OnleVoy2Nko2VDwwQKAdqtNm0qPlz1VZxvCIrS
xoMcDi58w86puMmVW1vIowwmO2jyoMck5d2VJ4s4nejv0G8NcZtA9lFIiKMtLX2R
W4J16Po18dK/P88v2dl0nrZMGEITJJMyGV/kYsxcS9GpqOhXK35vsXw9SXlaEbym
AjtOGPZfdkmaF0TGTfZD0vZ82CJmkGasNHOe84/XGD7GKN+LiOIUB6OVGAEvzZhY
PnGueCUy8SXR/fFW6PR3upai2uwMT7VeyVS1RcQyyS2IBw44PU3LPxTGX4nj+J4m
8PkquF561diVwOhE1oWnlcVnSBJKF3M8jHreDLUjcHpFiKVqCxWJ5ck7ikh1hC64
rzyHw+9ucB6QhxhG8WJxFmUWnWlnbSApswApHXLZ987qi48r1kt6zd6xSIG7lzb0
TNWwXwZByA32pnO2VYUJ4ZmDf6tgFEjqBRBC4s88RgJRhjC8dbjx3BjFAD6ZMQbB
au1tIPjFmWOWIayNKICKwde2RSqpGjQZ6STWaGeUlQ3kaSAt1LxC++k00vtLid2z
6ePjMLZIJoqaVbrpd42Dwm8hFh9IN8mQVAaWbM7qjzc6jh2HMuY9GqoZqqL2ApbM
MPOfXeZHgjzcU8oQS2Bj5yHNPquK4TJBkqbVeU3OluGKzX/09VP2gRT1N6uT5FiP
Hwyrt+VIM5mfuMs/a82Ru1Qt3eUEn7S66x3BmgrbysomkSel58vK2LoKaGK3owKA
RZCmk0893G5eCCjDa3Dr0WewSACpudrBvS+d+jEefbchu+f6jN0MdKr5E9l8fmvm
tcCBGFTlwi4tIrKJhzXvTLd3A0u2cXabWSVFH+Vvw7+7sQ5w6r3Jh/JvpyLZtpao
rhjQIVS2xzxD5L5OuWvRvkanE54piomQ5vnv5cWcvQDq+oBlkj5qw+q5l+rgvbEe
zVJiKvYQFSNKTHOpCmc229Oi52C1BXahYiyDYXLWEskQaZkuAOVE4I2yo3Crv2P0
dVNkImiQlinS3XIleuK8RbcaPO59geeb3hIsoXOGZyAGpWvlQpONcVYV+eH/Wk4/
dIiMvCyZJM9YVdM94Iq8rBsDZgdeb4Y+beN+qj9SLy4RHITvmpOvPfO2pjNgWUoN
zWKqucFTKoBvHrwIVPbpT7AHBGbjZ8QO9uujvaK1O73ntOj16B2XmoHDMjmQOcv+
Lrhgh1prr1TB9L3eRNhksvCjL/vvOp+ciWJtqvjQoSNaz6CSMY1ozLtDZGRPdlmD
p3GO5RCSA3dG7IhPvIp3h/Li7UXNPG4vEAQFzPfGeeSm9QOOiI6PcwDloSFsfQi2
syasxupMWH4AmNOQEncR3m7gG199IxjYfVy6AeGYbOY4LfCHXh2RIioQG51VwOur
VgNJEPCH4SazcdDcuaSdoTzKfPEaZZsauCFAV7QawmnkiNcrdrnEEVch97ypkb+s
CGeMyPutzb0aX/8ILEUxNCXTow847oXnHHvxQ4SzEIcIV9aW/Km0SHNHmZLN8/jQ
o+wvJn4y4TlRdCndT86NHU4JpVcCToYVxYdpp9Hj5GrevTl2ystIqM4qNPGkjngx
1L9IkRXmEU5zU+Da7WRWJtImhST38ECDb4HPyHYFFf6t61WgU0LJBvsD0z4gBFTb
NgADJJwQKHeUxLeu4UzXqoJ1fROgzVuYAbNCqXFOXKcwfEDS0j8VKURIDkDx/tlM
WV2kksNIiZ95viAQGmTt9Ge9NHmANQIwi5LHoPZZGArP8d1dOsL/muGE6r6dmErF
TmqdeqFSG9960kCtbBowGnbKPVi9FYaTHPcsI3pYU2DSh88JVn2YsP/uOWNrQC5i
5adVggg/Sn6kVRP9DyVzd+rk3b/aj0kFI5gL7pkpjghR+guy7uTRaz5ECt4NaasI
W7fYHV44cR+OPyJbmenJQPopq+5C3/d+ALXACubkwo+INmQNrW0pzsj2+CafMwA7
um1N+olcy6R+vyk2ynlpswJl53dctd3UsFYfQp/UrlmwTDp1pA4p2Cdw/SA5Nzk7
MYvFdVahUhfZnk8ZiCTaK5v4tX+5X2wX5KCm7+oqtBa9G+wE7fPrdA9zHQXo2XA1
Zymqkncu6nsp2WDQS7G3eMDBedKTet89bc8LLuaWZ+xRspkqNOSx6BsKBiA+lsv9
6snsje0jbCO2HtpEfmS62sIEccASjdp9A8vlvl1Po2Sz5YMdgeJiJbIb6zvrtJnM
fsLHL/uLxOonTepeD/G7wHrjwvKaxtwCq2gRqoFT5lzyAHY+lBWp/MnSaVHmRVlS
ewMxwGvDbA+OvcjAalZOyv8qTQ337NgrxkXxvtDLwGOS8HwyTNGSyI73iujLX6ir
OHPBXNw8pUhtlZh7sphxumouVYAVlYGuiwvFgdhD4Ucg2p28biv6poPAvBBUGfVo
sdtglCP+yNaR73bP289pKgSoqTD+avh+JGGwyGpbN/oPrrPlybjGVn1rGh7QQlEs
2P1uaRnyyJRywCbeaG3/aunsLNFm6+zVnO6zhX/FjanK8PYDqqp1qjIu8lVKKPd6
64kgcChIifcJz94lXWagEmpW0qN2EWSf4Ug+OEy32sHUS96jnAaOo2ZU+OO+nZ/S
k8X4ZxgL8suusXaJ8Mytwocb2z46kyHWlyW3T7Roq052+aDXVrUf5yRcjri0Fjg0
CY2NGTwz3PjVEjJjVWZrr2d8WRvGX9bC/XVLpLc2iAyruwy2oO+P+vlG9AlXrHQF
cyAyd0KoHN7Hz2hLCoEY8qDgjihOo+1mbSMqhq9t2zJ7HwLNOfDG5Q5Xgu4WOY+m
2Jortywln+/y1SgfItQFQRiYvoMQcov5j0CfVkHNEcdCUAQZuvJk+WPtiAb5jeSY
6G/FBddk3+ttnSEZwE4ZOT/2b77E+pKsRzm7QG0ccNIH63A/jKKuKwc4RdaOdyzm
QZgFIA9CQ0r4qXr8h1O0fW1e0cXYwGxSDTz7SZbDIt1GhOyyQoIFSj5FT5kOaub0
przEl/eUZXpk4185mCuAFyyiZkAPb7PdKcVUDihGVh8y+VPNu8hUgUY98KJYFeXB
1NfoA5PM9aDZBl60nH5ygb9sblkltQjf20gXTFUSkIDSaN5rw9uF/YcAKm4Y9kvl
A5Q5Jw8nbWBBl8NrELgAx11jzHi3iYO7JjjBIm/7mCH7+SrECarcUoKGGq/YiCjA
z5E5vxX64YLQM+bjz2ca4cvp0KZJwBTMQwlzJw0Ofd5/+8QLmw0YVOEQrJ2ojmbs
JOx51E3np0DpoxROlLWc/fCUUWTHcommUbo6tjLFD1Ay6vYSXGnwrQluJg8YSQKS
tV4q5ai02daCPXqkEV8N8TG40h1tabJcHuR3YqS5ULygYQbGseIRn3XMnLP2yDJ3
5c8J/PI1/vGOmJknN6Cd5zcjOqvTLQpp3kyQptB40Bnh+VU6vaAoFntiPSveezPe
5So73plhMxB64BpwmGQIc4iWsWrn90HfLrUn+GkvzSltqXok26bvnjOd5YHcmova
EA39wbxJePIZnhlO6+MN5FnLKtAHyH3+XUuy0u8D6VG2Ef3ENkIogMRW/awOG470
GPyB2PlPWQgAy2CVVHJtL9lj29spXbdgEtK6lpm9zP4gDy0YriwxMxMWu4rGv81R
7ofpaqooAwjeXsOVRIElRVrPy2Tc+vhBMQod0yEeKVUa1Fur+7fi6khm32h27MQM
xZHoJclT3FxplqHIoVBy2WhoUEh1e0uBLfOLNCrKNwAPBtST/U5NTobp13Gtmmxs
oUN5WQUtnsStDwZw94v7KsrqHjPinx/dA1h30rRaH00WW8GAuiTdFg3AeL8CVKlC
q0u+S9DWNM6F9Z2fhz/IRSHS413GfOWIgIy6K5cPTmiCB1W0cn/Ke4YEzg7NaLx8
aoYe7XnPR2An1uJLfCzdxvv+F9rEjt0MTc+Q957hy1nu19vTHTki54SWQRes2yE2
Qfj8JpGVmcB7fVIUL7wcfaVSemFsuIrwq7xGOsW2/95t5jjjIeiMf5I44C3uE+pj
U5Tbeq4xLgY4y1Cqu4x8JOTDvyJB9Nr0+K+8boiZ9I/ynVPKTCsq2c5HmPOvGB2o
LOXjVgi2TqdxReSaE4+Ud/vMmezp/bgxAF35igprl6iEmj3TqATC6AL3MfnuH71c
i3YnjmZAUzWiamf3TBWOnvRd1Bee0HdKImMETZxlJ0nEvj3d3V93lUFKxhGJcTU8
qQXkTNgUVg0A6zU1minwn3sz9JZDph0ggcIly0MxyHuXUSIPSBzMlWJBZoWj8HYR
sJ3wUrVQITagtaFv1whyDymrRQdhDeDwGkEWXNJ1dC+cgl0he1KavJBKaN9YTnzj
+d3avXtkZaK0UKh4MCzFOpnseg7zzNGz5uhVKsZushzgHqeBC0DWmhNpkB4yfN9B
zMvWMuAZMgqKqEcGW+/HDV0vA/Uh8CNvb3oXneQNkZgcztMpeePm1GsIuh5abuPK
j0qu0UFCfTqjHYe603UvgG1r4uiGMjaE1QFrui8DB07bmWRtcZl7l7HEQtkmsTM8
N07SSxgYXEsoKmXrAA0nsIiFppG8fd6ZV26oj6i+f1Y3uVhilhPOBBdXXzyrbc5w
FcMERBUsOdXXseg1k+0nqexxyFs+zx9EasFpZgjBxJbOduCHDqcaFyukospgUNw5
QnhhIXaCmiDnDZrS4EcCLJTSFho93VzuUyKTsRtznAX4Hcel8sfMm+9m2C5QOGiY
017QIEHwpZysTKSfZ6dGcCKLmG9w4m5L43IWMGF76fzVCXSpYbHn1xn+sUh3oD8z
+VJTbEI75nCuc6VKi3g4ForDAyvSD87d910OkOMG/yVBV2IPkpd/w73ZT7ps0KL9
3cB9NzZvG8DgVqBBo2pR9no+Nzk8Vw2M0IlXciPbMrfmSKCkeLYJD+xJowxgnp32
mlvLqKHtovkv7hnW3p7WmYMEAdkEzkXX/zzRypx3Z+uFIe1ct/UwKX1sIy3kHrWe
bOAeaWuMkXX1MB99lgVqqHHpvatqlGGt36VaF9KyNMVMQRjX1cVwGLhNOIP+UNjC
ynYncQSNX+Fv2WWKGwgss6WxoQ3bruYCEa9n7mSH9MYBA8C1xvgtleqb3QOL1092
mL3YTnbB6jgq8AjZFyLdbWuVpxsuLD6OC3pZaRYQQVvgtG6jg6HwMEt9RkPoU5YX
G579KGwnvQh6ipP/rd3F6g0Ki0+HtwI/8x5BpopIZXb8T70+8Mxb6dHZWfDDghMu
FK1n3nLU1uZScmiuSJBIZgxg6xTESo5YIeIgWcYlcMcQ9N6vQRxx7ALOP6bCpSj9
l5+tFTMQOGNhYEig7Ga42p6P7niNnFMg7PtPpHTFCEh1/XzChIbLBDj1Gd424LHB
M1MfHi37mj0UJjNar2+uTbtJWRZWUNsN+wIKExzcPjlFNYDIVB/4WO5Q3yHmgLKu
CmpsVNW8QWN/ZaYAH9+hJyyYzuZoqmLkux/DCIF5TzvrZwUBeh9j7whJBpOscmll
yxHLJJQxqsiIRMdD0V2gd+M4hIGz3xFj92DKHCMsX3R8JutHVwi+Qbi6ITkNqnn/
Nbyp0wXGaEoS3hyvzKJqpwmzl1wwsnwaTcqs46CrMzqPsuv7k0k6aJzNaP5R6kyZ
X2GlW7HGuAy63SWLGfHI0MqPB/VX1qzZMw0LIqKKuQSGASfseSM5RW7+Wkp+cQc9
kloZs/pGMjJSXkVZBfsxreUkYlFnUDcU2jJEny2QxfuCI9RzXwkeBXWVvUJzx4Ep
z7wleU4V8hsCmnmffc4CAINCfA8bcNKsuUwghCGt1x20+DjQH970Dg1Q0gi1RFgJ
9N/GXfWWHEdtslw6bK3u+NlFQ3EUi/M++dbngY6Pt1lVVJwZuuH2xjylHSvzzoha
mOfjge5kfOyZxmVckTP6ZUUwi/MsuwqeH9i+K9oHT1oLNCCs8dtOg9cBWVknAar8
EPR7nI2ZAPl6rm+VUIFcD1kC81f5OXUkeGxd1asCLpqCA+y7hCksmLCk8zZkNsYz
dFGlRVnQcNysPydinwCLLY3OOmO+vOnxuB7Xw7HWLt6c35LA2b3CE2qHTHAgwXqv
vfuXntfoTFZttP0Qax90XWVmGmdWkVagkX5s25aeqXotwgagmylS/kG1sq+FdrwG
90ieIoTMYVf3VYwo70G3QK/704Ik7jDNCXpR6etPkaxWOsuYvH4Vlu5Ien7A0hal
fd3bCeZvlDKGHOggR2hny7hdDUfYjcNgEkJ7NFG/V1zlNVm9iOactRndS8QO2iG+
LT1HGn5dv2OcOzYynzhmaJlFz9iP9VPAqsfnPiu0HJ59xi9n7e2G/W6roTBoI3bX
nilh68dsmZ5VJxBK5zGnkeOuMhfbNrPAa43+91gxIZalbp1JHuyusHeHwfTSjBYC
4vtvh9fx4mlTjaB8URtrTrFkX51+AVIXqYq+2Dt5Z+DNrkco53hzD2RuOUGkRdvu
/j81UCtKNUQuYxx94q8odZomlGshaGcGCYlVl/JA5tkevPmo6pleRP6qenbzOU4g
yGCUk7Q2cwab6bMfXgWPMWC6BNBJcVkFJD5utyVbKGVop6DxvIAlORW8d+1Pa9Ob
3xT2YPA8Q1dc5WXg6mJdNE/3Htwizf064fzCsv/SWrxWKIqSEeqfYs/XKuzs5z82
oML5TmLbVH8hM1SfiWnFxlAvaZJ67rABkTpu9CmwhO3L6eNxxgFUXXWIr47/hDYt
rCnvK0yud6BwttyCKNQ4Oz3rzfA6uxjxWiONIWQw1hRT/L7MWBM12T47ZeyseyFJ
gSyfrkurTkyR+5P3nrovOOujwbGtDk69KSYA/rBJt5LiBOggdx+no9HkwcjQSQjl
PEItir4/6V0zL7pfcnkMSoDWsrBMV8Sw3HP0pDy5S5aO2RikwtcOKGPEB7s5HHro
vP00OCs21CYFQoImz80t7iZ4Ao21NFohQIjnFYcogHUADSaBWEEK0EBOoGf8sPnA
GOfw3RTjOTKVTbq84+h7+tAlUyHT1tdwL6JNtv04okRPSUxme5EaCATPAhJZBhUU
hYsNmzYVsX96xCjijDPmD+Hrkk3POFrlPP8s/EmhhF37DwAjg1i9oObdtXRfHKEi
hFDsLCZ/XHombuJ1+GsQgSN2SngCQ7Mbp8Nlda9EUllr8VYmIjvKsB680IB7JVCc
LKUBeX88ZBbul+46JKag/r3BP1tKuJsU5dMvQ4HAkb2e6SSbu/m7QY3MRkL0gavN
S1JrkMgKrCqvYabLAnG3efBzPvLnGlNRzTPkClJ45y+PmORtxSEp1DK+164+Q+G7
kcRo9/dqF+N7Ofd5PBPDhz2qQbS3sOipDpF1ksIKMNBUamI18OU4Oxc4jAObDLch
1YqYJCdvL0KbUn7azyYqX84E2nf31Wx/ePtlL/Lc1XTT/rKxresiww4Fax2plYX3
wdyCLgjIdlkKTvEI6y/WMdxhidhRvzXBgOJzDgDnqGQYWEWRqsIKLab68qOz+bpm
+B4naSAB6Qc4CcXTVMU38l/rCtBNF7Q3pfpIJ8KmMEziCJES5hu1qKAh5HMFFhhA
7S3l/QKeFdGf/ADBvU1AWVkMfvoOvcr73X1TkflDA8Sz7RnC5Rdyo6uahM4w1Exd
1AH0jmBlUy/fcFvNq2HiEnYrA+ttgKj0DdYd7cO/GFXG4SA8jjIdc4KJdjxQek5u
r0Zenmhql1Kqplhb3w/wBpytwt40kSMkN1ZNbnWmOJeOC1i/fRmX3Ju7ZEQSY7+B
OZiadN/p+/TpyHKzVcvPShWE1qTPO+qgumH3BTs51N184kqJVfGVH7irqoqlfY0h
NlKpycj4wJDwflH9yNoWOtFeCfMc1ujR0V6yc3WwSAWuPGvsYjFZrpTXFXxy+0Td
3+d2TXNiLFrh164olBL9cheTUJ5COY+2WVfyw8snN7pxBLgfplmvojRk/KGs2Fcx
HQUkgAqxR9Y7ST1YFnMpDa2VbKn4Fgb389NNcu+mYCZgl95ePz8LGlOul9hOkmb6
mc3wFESYA+K6XFhQPTAOvdlH4gQC8964IgUDGf9BFZrf/JJqlpAqAnaviDiU9773
mJVxEYHwxE20VruSddPODmG4evokKu8zC/f3gydXpU0frL5Kl0YRb5X/ECkLV44g
nFUOSq8iNVhfzhkeslqZ9E5smdU1cgM3DPPLzNSAq3NY379PaEsnfY/UhGKOLhMo
1Jew9sfTthJInnNMBmT05GbDxgrXUoGZtfqBZZnTAQkkAGokufyOfqRwFxA3LTXu
ZTdVNKtjobk1s3C9YD6U35KfgnMSDeSA8aFoMSz9qv8Rl3KSzPC5xh+RO/Q//YMV
a3Q5JGfSkz20IH2suN9EOkYoZyWkl9ivZ/OnZcveG6zcliwC+nNQI4VxLevGjyes
nxsKYiFthG0f8xnM8gMLfqAor9ZuqoQ+SHRgU+Zq0Pm9OTGYkYbhgHikTbubGLNk
UV1ZcQtHbt8pOTlBfOwiBGhCDDfIbCZ2RyPZiM0jI2dsVvH1tyLmDDeNmk7hlXoA
ZMM4olf/tLO0mV600WgJLqYHWqwAR528R3GXL5Uv1R/hPjlrlXkXe+Bm0ZponJMT
LTyLsLdd7/PAL1aL2GKEx2EZ+kWoNdRaff1vvMQRVgGKe8dzPd8WPp8980g/QT00
v19w9wLHFK1FXkBLQUZWPIie+aRiXQWiKWZvtP44PSpQvYFAn4DzsApQbsA6JI0K
OwhLZ9T0oix/NRRwChlXyCc/F+QHlH3hZpXsoagJdoR6vS1ohn7mKtejomngXxIZ
uKcOAcfVoQAl5sMX9liMWHPp15wf70Z/ABHN+Y09QCKGEU0Nk0RK0SkIkkKNveuK
MiHPLTM7/DQtUddYmLfzLiZ2L/E74XLJwOlI0C8vzcQzeOTXHX6L1dXO4Vn+Jykw
pd0JpHIk9pJP8FSE9eVgXNvvAZ5Td2mY5PLyPxPOuVlqsGtQOVWUzKO8v14roIWE
2E6A2nkFU5DC4NgyjiZxYDwiSTVUPMIXQo542GS6T8LHRgKWYzG/NL9hlJ08YPG4
vaduLqtkZLiWJF6FccyKr2ALZjIHLCEseSjrhtyVO0vnt2cBQLqgA/ZsX9VV9jK8
xqeMTWbRGAZytoMrU6KVGIGCeHJY6tgOF3hPI+xj+8GDbDtV9n+01fSFjPGPVbcI
idvdxjAk7K2Qd25FANLp4CSmEHOIVQJrar5jHLH/cnUsog1bR3fcpamd5srbZjUt
TzzLXILO9iFo61hEzneJZvCKOrWHIetftEcca+0p88TrcW7lKWTVctjEKnkfI8N4
ULFaDc2RMsywIcDStTcgCFrxYumrNxCiqU/G7+djx+zvb/1uoryvx/g9kmOPRG37
XtZaxV4qDZP/768j7Yw9/RLWO0VcB7qEBBFnvdZfNPVXCbrHyhunb6Oa3wa6b+bw
ELeQ5xIXJJswoVgHjXOC/K6tFalkz1s7VijIIPNQnYqBLoZICVIyz8QyvkaHFr2b
5sWs5dUs1fZyeEzEMjrkUVqEswa1bmoG7uZmXf9Oec/3jDA6Ana6Cvr/rj8BrhI+
60KVhJMduEO+F0AvJgWT7ZG/uD/e6LjuAh2PO9dm3iVvXHUtj8m6gc4yNFm02QT5
/+nSTKYnClMif9OFxHl3Hq4eyrGtJox/e9VEyf+mZW5TU3gTgNDlpMZUdFAJ59fy
qI5NWbcEzk0qbAPWaY6mTqJTNMERslUhrVtIY/0eL6qGi+dsuIhfwuJJ0WxtZNAP
m0nXrMwyFSVH7+S2H5FHT5J0+F/sHrROee3KI6/XfwdZNxHbaMu5iioBlOtafXsQ
ql/ySrk/Fdt+4/3jj9YujHqaSMq2yz9ntla8flsGKx8ynOuueNueGjSaSEDozZco
ifC9IMdjbsLKBwY9nAqIwB4F4IQaYBsbTF6V0PzsVzL4IcwhhtLRG4qiqpUM8E2s
eknuyRO78ZKCPlQDxgXHjwelaG0aDQ0nJXED/yP0T9+ypDTa65ZlW9EVryQ3hded
pJxFMaQrYqqMyZatZVnycU0+5RCBIHVUw6MEvRtgfiWENkgP+/2AJQY9F/EjdYhe
LLvMqpzI0YqtoUE26/D9xCzjAk01XMATetgxFq9Rsysp/5wJ6EzhVHSLMrgxw3dN
LoxNqQP9ENi/0vj1OsNn4D7yysQKoTqkCUFZZq4L8gob0rQmJ2IpFr3UEt3koJ2I
cuprrIUjyHzMrH+bzm9yupByy0LpqmoUUKK4RfJpj7gg1bZ8wQZMrhKlxJPNBYPp
6DhD3gaoO7L2rXafhsxXuP7mJPqm4QNZXpQaX4+FIl4awuuNAGpjzDGiBThd2E55
21wvDjVkf8CBVp2qlDFbTd2EWWqAYN9VSoLADpbD3hH7rht1mNsSeBdcEQVcTN36
ktImKbJx4LkM59hpvOUoX1QJjwZ241Xr7THDsPLldDUtS/tJ1om1YUUfwzFXEqGf
vmBoO1vjPW6Y7jero1c45irMbSOqTIU+MVsGGtcx8tiJcc9Zvmd4LeWFycrrcRcB
b+lppUuaZUFb69XkGNUX/97AslG78GzApU3k/HagRVpawFV4PsbOz+unGvVNXwQN
8bxwx73axTs0ZIj8C4L7lryv/Z525oUkGs5MWl86XsL6lYpWD6s2mtM2phZjmZQJ
HriRTv3qTylanGFSXNzNRQetmNaaqNQGCqoeZfP5st+878G7Ujvvn2ZlK9PaLyAe
F1JAHLegcGC2riwyAuCtIOGVO44tDIF8quGbkBvKANihPkHO9gpn7V07tJZyJHkt
v5JkCxf+JLcddNwCIhSAZVSNkaApgANYu+FjWGBf3L1w5cncc1HwrrbeY+Nwowox
HaWMTu/G0raIdR6EAY98iGdDVWYS2j5vgR70aXAWxZ211zhMwUDTGBfhy1GgHVq4
Fv9DgElSkA+WrjJ+UCmTjX0QZZpOG9HZrgijOIjEfC1a6UzNHiRuCFg8Yoxp5+vc
nZ7w5Bn7y5QQ0SuEe8W11rIQYE1JNxO4e+n2vBDZ07+qxnNXSVfq8uUVBFlkpBpY
C6YPImd7jL5r7XaEDbWZLQRfAUn8bll+2a+Z2CgNJiMYdURiEXpAo0wL9sImiFVq
mcI9EXtrfmJwHfOfmUOYWfIaWjwZbiF+kXI5xdPzzVMabuo8jwONcFSgxIFZ9qGG
xkRUi/td5MnTtRcsYMYNbYKssOoDm/5PfuL38UNudN0W+dxqck7UyUW74kjojTH5
ke9uRpXp6q0Eq0cY9likMZoNHS+V1tsahs/AsAMidEdBbxSae6bf6p+TsN25KFwG
yDm1Mhri4ZiAAZAzacrzrSRCZkfSrLz2E3FXRuNtx+KvZGymkdvvZSQES9VhPHQT
q1pJzyWdkDYULM8C8ymkTeKfqsKb3K4JBoNMwKI8U8PQM5iOXZ49EgOBVqm+BX3/
m01AfytAWo8U4rh8M3jKX/HNPBXmMFcMNHJdvBQ5jkPHIkR1GUdWxHWYeW+kREzm
Wa1IOglq58/kfSdeDqZFcN8j4da6/rqJ5GPNg6kMPAte1rLn90r0XIPo+PLEuTxN
jmeO8mjkr3mfkAO+q0HaG4n7K5u6X/kXbJtNEFFl1qTGTnOUVd57Kyu9RkKuyJMx
XYkLIIpPC5t9D42kaxJGpoyg86SiKUAIchONROvpRJU6numbl9sd4SAqeoDfA5v/
Kyc7nsB7KMNteEUgCAifPRtrxPqX2K2i9UK8KhElsCgv1TnuqaZBCX+JQVVNPj7V
lmrgsKWIQ3enZPp8PnESKsU8lvODLuHNcD6KoAnDqgznKH8TGiq9t+sVLycWjTyz
1jDvLQiOhf4cEiVeDo+QsoMqu/JwFJUllQ+fto5Hv3iK97JVEGSug3sMRfuHOZAQ
Z1eicoEsqVWgyOJP4up+g6bnzZsvNPphtBE/rHkfJqTnjHDmAji5NIgK+Z0btdHV
qkc8/92aDwiEwxodM0hbrI/2VVN263S5mts2jwDcTLAd9uDM78uXvJxT50WpdDv/
z95JeHW70Jd4FScuQ6YWMLm/ckeBg9hzfnGQ6NZ3iyOlMKA4/yhGDJMrXfhmnhy5
JoNu61d1cwbLPgZAUnHKp7aHzMeLRYYaWFHXpeO0tsyoZ+Wz2/zKIQPn3XgnX7gp
f7UPpFZKpK3qtFq2R8IAQBeZNNmEV3VD+ZRJjoPazt0Ss7c8QuqgFJmH6fZCMkIk
MdML9hxpMV7++Wi7HOZ+qTrPWLHw5iB7gVuybDmFlL0lqUcQcS2mpoh4fDgYvLLR
+KRVLX0GoTaC3URF6Nj1DS38SZI+UnMDNHDXPF4w5Ibmvu4jJ+nYdXLaX0LuDBU5
5CIAycegF+dZV+yz0J/HnBxXNuzG6sCXoclA1iwZGA/5qLAOHmWSIun4KZvPgNFp
PuFXfREDLwN0pW+vPueipWB1rvK/ChEwv//AJmANpglVAraGsFt9I/qaRC/p+tn6
ZdJrxp2c5Z2eZfFPL+2oB11uqYZ3ivmB4YUkX5LXcuXJzhukswrjsegmqfAP5WfW
e/4RoV9pYsjGdYd2yRMw9CRSkspD4XtQHPYtTWnmd6Jj5Tim2Peo0zbxfWZcHx72
VUpoM3BXHbuVHUDmfNs8PM4/+P/ho3fkQ+WhAWOkxgRndbidyInAvkbrtsTa0aRk
Fq9fuL+U396l8AGa9asMBdqY68yal/citrQ7ZvUoi9L/VYy7cX5uoOXWWRV6B743
CzsYof1fNxX0PRv1GEreCF6q5O7RXlIE2lKp/dMYDnb58SxjM31N4Wt5O/AJjBAi
53p5AND7tKD8XC6UheqebCnZQwJ5l53wjSTtN0cDo36Vw7HXoGqTQA/51rFdKKSo
oC5Es4iUpLvMWc1PelB2+CgQ1uLardh48nkevzDTaOT6ae05dosr6neJ5oS6PAS+
2HPQ3L88Ikl09haKWwHgd2TkRLDvJ8PB2L+HZQ6sd3WKLUKuCV6rM3W4OCK6t4A0
V3m7JA1naC2d+tRt40kQIjz38wcfXswhJg+ZBzQSsDjm7eeTacvtR43Yxv3LG4Pw
vHktn5KbHpq3m9c1fudrz7NLDDht8X8g/aX8uJT5k9qmAsSU+ICwP27q6hBQi4hr
vTU6G7eMUxq+46AUkIOcXQNWNrYKh4cyP2FW8Z12kOSnkqkfCMOcN9ctg7OGK68t
lz4kyqyUkLI78mYyCc6g3NykmlPxNVVcVd713llplAlFLFUZ5D8GS530D0HQqBiR
ioN9oTSR/6n8OgOaaJ4htSHfOQaKXl0ayctKZORhMKlcGPdiIrwxI07LJIgyt9OG
5dRuAbjoRQPy2/FwGQzgWGIMK/zfA/8Yyio2cC61NOdTu72+0OGjkQLbkaC4lGAq
50cBjviRUBwJALbdXYrk5tGLZvfor5o92Tsld1enYOzRkKTLP2cNMnqKdkKkANAR
dSoRnO0kc8adYHEckW8OiKjTIG6KT/WqCTYxHXCd4VSrWpZOAvFzFg7/N1UHtgI7
rwfCN/GMcC3UNpSWQzc4FvZ8d1lqjLo5nrNVSWOPpqLU3XXhjAS8U9qxhc09j7Pa
v7jGqdfpSUPNIqnrX5mp9kt1rMvMzLJHiRniNdSEofqKZtzEBmLzLrDtkKLhEd7y
q1IouyJNF0Qnr3iZShRW72DuLHWUi4rlwolMyMMSn7+FWklft+fjldw5a7TkCdYR
J1uenvJoeqlDlLN8jieGlmTd/jQ21Hb6MHkq2QOtMLtJj+/dG/1ueW/Sh2THpnI/
2IbmnjHAzVTBRJAOj75cTMXWdb/vlazF3dlU65MV9juGC8o+06KGtxn9qkhl0jqI
kOAOEu9gfkajRI08ryKXSmTVYs318ilysf8tlLInmSGERxmqJ8YWz1vxyT+SEeps
g1zyiPMKnVEx4RAeCWK+4NCrMF3xlE0CkpOJ7AK3uJ5JcTDnk/retYV/zok1Qfjj
CmWowHpmS0Kd9brmiJKmEfJ5IwFpQ+r14Qiw5XtV+UUhrnbLp9WqbuxN9fl39yl7
JwVTeah5d8HPk0w6B8ZQQfQUmzb0sn8co7dmGsCyDBVS4m38lxpe/aArPIYpL4S9
P66Y1h1A5Ctq8v30sClutvotnIVTb5DEhJc7NV/msXwHJEe5Mrz1VqA2MzKSpybi
zPiyPboenOLfZ4WvsfvBz2iO1gYbva6LA2AzpUoJ1KNGYaywC59Pe1002/8hLTSu
IIieCru2j6R8ek8rsUNW+8S6kT5JsNU/3qvHi8DnVXsgPrnfB1QEb7jImepWe+dj
nBOTYqoQavl9xBjMS9+vbcdRsoT/SvQr6ZPvXHq25vGiDyoEd/rZxNSs6u1ESoVE
iE/JOyMwnXNdx9xdodxCD1VNQwHnaHkL/YmNeDNNySPuoGVLwP025HTb/SmGhjhN
Nvof+GepeisjOvCvMwIIjxICfmzxkWT4LgHstyCQj1MqQyFOvj6XjpQ87KApsVEf
OK2q1qg0+mXAfQ3Qn5VEcrSdC7eEk0pJcPxqtCwARlFZI60z9rVbyokrUM7Kb2oA
buPfv/54yViMTKYVJlYYqnSndCxxmmXpxIFvwQi+8cHeVJ3+a+Cs2BByE7j/5Lvc
/ezjXmXcPGXWO0/sogZxubIMJK7gFKFQjEj1TrNr/2Bb2pzw4/nOnOiDR5T7YPDj
oBQ/3wv5CxoZKHnKC48gIZwtoAOZahn02D0RZ/hh7ljjoosnSXSFGrN8PIGF6jyo
GsWvgO83elIsgnGobuG6md7LywSmm+fpBm7A7ULU1JEHfLoxyZ7o2VDZsLnAuq7D
WU12kRPZrJj0LuV5tEL/0S1zsqEpDsc5pECtGL/dQHP+drOhc1s78nIfo2lhkz6m
6cjisNoKbJAakNWtRcI42DkhwSs3lXSBByLbfFMjH/JXgyLiK62kDTbcJ6YlMeXq
BeN35HbP3JShDZMhyBTOD+giKsfEzNY9P6etH2mv1BDlow+QMgY6W3D7vIY5aQSO
q/NJIlP0J32dBDHcv4y+8SdRi3INKHuhQY7C7fEpxvEXCzmh1j+Gxue+zBJ6gECE
+iwYmrzFapDKOYaFt+EW6bUug7OcQSxci+ArIeUGMahQK4KKDIbefjiOzVyu9roP
ydbdemgj0dmxcjncYxoD4KzrEQvsv+Ll/D0mybdrSlM2unA+gyWDJGYMM50+KC3h
wQeg9fJABZjAhZ3/p5dZSplbeN6x17AeIw0YBg2q8t14oRptqdI163Oql93gUkxD
wBBwsN3gY8PAbOsJsSJTZesBMDN/SRCK7ky7JvJcqq1aNhFoBwmsvuMxjOORN/gP
sosE2YocQlNBWi0JWymeZKjTQqMugpPTp5cDDIP1CVur0iqfyYGd25yu4kToz/iA
JmE2y/ZNPQRuMn/aE3uxGKv85Mbm4Nw7daYb0rMkq+Uc9n6npbEzITk8JaHGxL9f
hGBXFbeGYTeQyv6hz6PIS6buQ9rIsnfx0yPuLg6NAwXe2X74+mD3A8CqdGESuyfy
2dy6NIC2z23cmE+nDz1mkzmrkj++bqt2U3U52Hh4ClceflnqBmYqCe7bgDUFcC2M
XlkvHeu7Y8/gkPumKnRJSwUszZpxXiyORyV+vT/xwa78iLHPvxFcTEK8ejoGbEB1
9ISg5RSzflj1AZFYE4mDaR/6Aqu5mcOaL31W4KIdRTxhBzjRU6NkwlaY6rFp3NHK
Q9RFcmLpfJiX5bUD/B9sclLfgA2YuRn1Vd0rv1H3KxVqzuf51eNXBe2W1v6CZY+t
48C82SCG36hpln6wbSi5SXK4JzdB/uYMRFhRevElZyx+EfNTkb6/1RmvQZMY7Q2d
p5e1ov6EfH6I2wEjWbF7X2X2Bz1zmylr5nvMlnqZXaYkFJIaAiy3fAXamNCOq9hv
AJsabhLXaAt0O4wbMhDrcbFZMYaS/t6n9hRyMjhENorg+gEQ9AiPac0jvIF3w0FP
V5KKa6BETbPRHxiyM41Kf2p8aX+NFgZQnTFqwZBxGmcdMh0DFG6uctxjZs1XFk7N
MIk/5HTrM/UlUa3wLiCh/MRqJY+4+iZloKedeA8EXTA+U6dmUD1c7X+B9iMeHDOb
83Ddyhuo52iR0t6jrPZlSjuXGeLqWdix8uF+mSO0G79fODiz9UAig3RtWnhZp8W0
YKnMQgiF00gRQNSOnaJQJDJnFL0JwlY39ltuQxiLkGvQALFtqewuMNp5x8HEXN2T
MQqFJu25+fYdh+rgKDI2fKnzqTaiuTg/UI3VDa8j/SKzx88YFmCmLF8WA3InjY33
IGG2JykcydP7AOV7kzoggGHFBL39gQiHtJaGdAjbkkPKaaTz0mEGT0k5jiiEjbqZ
bpedMDxuQNoex+AuB6wnWoH+M+Wm2ZQCt+AkP0y5mk49GqsuO2V5zR1NvDU2tC9n
awvb2yrN+gGrHOZXhgKO0y8Eh+OQPKBuMbbUWtiREsJQBiD/Wafb5j6pjDChRjGQ
VZHNzKk3FGJfQMinNOGb27+ER12QM+u627XS8NHaEwwRMFYK0Vjent6whKA//FGW
C6WCF6kLZ0Kvao4lq/kwFclA7ES/5vQaAGC2zKE4cIwHAVJ3xI8kOb/5Z76ROHnN
wnb6BsMe/+fGWkrwmaYnS1D5WllvW7fy25HbZ174LHvZl/h4PhX95ccHBJcC5u+N
Y9Ui+5PAPVL9uqV6z5AlBbObcqikrViNa7POGfrCmq/VFjBJVjnOupdCnSLzp8vH
EQCpSjL31uemrzOeNrwN+x08M2Is0wjZ8HkMX3UJg8ACrvEgUw+4WklKDp7FyRmU
JYq026dl+dJaqHiU3rXm0sSODvgajVQumhQNN4aNqi4560BOfdTldZ7g7Z6+FPTm
VSCJ0ZtKPKQDe63nTWKiB3Ur0VThW1xl2pO7nn4DcJ4jPLvKEjFS7hqpAcj+Cj7e
n0A58AZPmZmPEaKOdEPKD4x5nmQX0uJpi51QmZ4aeMQEor2kDQWR02PJbRL+S/5i
9bCI5DJ+4DM68to89hcrS0mVAw7SDtY5213/JPD7jR4HF7zX2ntKaK9nOrRV03B8
ZLze1wk78Ro/gUecY3+XvKQYJuM8TrjFpwzBXY93sYc/MvSWRXMMxZ9UvwpIqyfe
3LrJSHyH0UnJofvhlJuI7OjITp1cHxjT/LSs9eVKndTXwE9fFzBD2jDl/mCx9xnm
Tf3deMbcpzamskizwq71Wt3zpiSlMwvAuBUFam/mQ7kcIkYt6/CVV+pWhgDHjz3A
eYbFKNqJd4QMGlGyssdZ1ekfyIkEcUWj4zyBxgEZy3TeYylFgWSToQB9fR6voInN
F2ASFbw3IV/XwFH8z/B4WpaX43FuCxTyE3+aVbi933cKyxl5FCHNSUpXu0CMf125
1Fu6zFgk4oSwRQUB+VMqh0QpIBhLQ+PUKrYZV2y1zOLIGtiWd7vscLol4ry1XzMR
obOyZiZ41fFPnqoU8ZyP3LXtYkKcyk35FsXpGDa2PufXbhKRZfciKKhphCptRKek
QS0BHD4NVu8p4WS3SI/x8PGA2g1M1KpwrdN9LRMVasPq3Nh6rrqmCs49eYHyUY9D
vOMcX0g5TajI3F4a397lhpcNKeQ1L/sGAGwt4JMs0HqdsAaZ9k4hGiyykgAWU9U2
yngvASZ7EWYUMIKDAOSz7WzgYgRdYnqH2RYvry8d8GeBm3bUduZ+6ilBmr+Ztcm6
dB1+4kZR3Skr4gkG83NXc6WNXJ/3Ec2n0uJoeT4ccV8zQN9b9GySzOnqs12iHkL7
3JzWCKQNtfKq6gPKDWKvmbAU2Z34y5ik7AgVksX6YjJwrkTsif7MJv0Szblu9qt+
gTYU3j682mPgqvX31e9Peu5BhSGgkBVa7/0xB91UfjnVtAHnYdOMS2NnMiofv1wP
k/voKLJfToEqdCAGoJLqv0K3/VTz1rmkoTFE+Rer/J91EiF12ulzjMwaidGVp1Hi
kEn1d7rm/6qXHWlEIWXSLc4NKxh9T+YIwkckfUnRPV4ToRWBAqSF3TBv1MRgcllu
lgcBkhTARk1BH4rKeulahZ6HcbmyMIc579QsSvs00H6ilSa8F3VylH+rLP9xBW6U
9y9MEpU5qrVHNT0jK52z1/igGsvJW4dHAQWg1/AJv19688c9tfr3clWLC9ndmUlB
KKYAmrWfQeHtYRxvdnr+AeZq0cgeq1WyRAdF6fIsJx25IEr+UOStl2rk6sDDI2xu
EHihXOCkoasIqKtU1U4RVm9jB5eakRyXB+0ytFHUOmQjDPYniJDu+IIEKcczKn16
qzPi/TrzY82zckhDBFm/AoGR+HUoDHTfAa+6jg9jdCVlK7/1YzRNDk5BiibUQ0bI
iBQjeymtHocSFg76OxZZN009yFTP1agF4rPSHKE0DWIkB3pa755jXBV8vuZes7hC
KhXboUN4xTZtoeMukEpWkhaov2UiH46NfUcKxhrVWkQlN65jsUVwmh1W+O+jrD/4
i19Ze8CDDyYAG1RiVhgZUF/LR3Sjdku67lojsBFiySBYbCAYZPQbLrb0Oj8o39EU
o7LjTYjOiZzoJVR8tMH2TKv3xoWMz/AG6sCrWBVV796R8q0Yei/L7TEnZVO/7f3A
jdlogz1Qx3JUw2vpogqv86h0tQJcr+5C0AF1ylaNZoyPvXGKi+32oS6Eq5s0SrB3
5mVBc3ZwMY+NMC/uPlVEurRBRFTpOo27HdcBpxDOMj92mwSvrDe+P6uydIVvBBya
sNalQidCNHvLzo3ZOHLWaBx92MdEs6XDSoBkB/ifpIg0TJAP+VttczkUX68V7P58
SH1aai1rY5Ejb6lRTL3QgZMMCs5xxV23VyqM8LdNicejqt2sk98QOr7qlALNZsmh
k1rr1wZACyWJmtDHUSrkprdVwZv46/bTt/zukXDtBEEbWC1jBMP7KiPmgKnKs5t+
WIwUXSP5CWVtAdulewbfIkUXSqGCn4lN5JS86+TtwrH4OCSbbR7y9RA3KaXTTAib
1swEjf53hfhFBpsErAnL3doKNHr60IKW14NjO8OVfpccLQBHK/+xpJDcLNlGAyix
p+H0b8xpEkeudu3cjoV7hqbwjPOl+oSHCNjjkgA80Usrh30m4azI516eZUYvrl7M
pGd3hMgiNSEc0ZtqUcUgRtGa6anohBEbxD9yu32pIuS9ptUeQl9PeVMWcGxxscaP
PAvy8lau8geqVarYV4RtCqaW28GnvSV/3sL6vQ0VRiy2CFlYYOn4AQ6xs2y8gAJl
xdLPscJWAmzawwiZW1zBaiLpxCBysvL5sG4hMqokYivDEXzqtG04UclUegxC0kpP
UaLysR64TDPjmR1ROAN0PDumj3RbP9GocCDP39dWhP/EFne6SSqydJ3kWIRchBAU
Q6rqt52Oke5D9AOPewr5sPq3xGbnBtgvuUJ5kG7U/6Nh3f7bGT31fp0TLuU8a3A+
VUq9v0njcBM85XdU1FOdS7Ae7vHu0ji7mZHzzzYW4K4yXduFZxkDeuzscc5JxrHW
M5WfrTSM3WheA/v7zFhcSumD/TfPJrDuPOuzjKldFRy1wEipVKY1cDv9Ilm55l/m
Vcqw3y9S3CPjBx5lzvBGLsTmyJnEjCigTOwPWHH2w0+PRm6ltNwVHhOe8ub6X0CP
WgbY6B454L9i+ZtOpPG5O7GdphJq41hHttZX/9qFQaftZtRytEk7RGd+JsU7IZ84
owJ2pCVMXzhTjx4wIp5xTKGuaAddrYYDYf8Mc8IpmCkRCL3KiGwDvSUxoa8VqXKE
yBiRgmB3KFqkfxU5/eI9Bn8Su6QzFAQA3M1iRUGtb1AbAN6vpDmXgQFH0125m6cc
nRF7+jw+8qsZgJwdwVQzGB26AFD2TRR9x2hdvD7NWLIqS3AVPK+6upKiyWedfjff
/eURqseLVDLaC/GBMYD75eIKgzonFYpyiyeiFGgPtXTPeriqhUYLiyJTE/UrVdPY
i+vwLs7noPOtMGzJixdticJetORy9j7acG1/HjIhhxXeKRJiNZ2B5fUkZOSUvyy4
KB4KkxYC8wZw63pBdZsaDlUq17QTreep0LJ8gwGFfAk0GrVOCcNh7AHuwPDPRwMd
XeAN93qE/Pdj5yycYjT/xDTHaRZrrxKPZhjYVshRPq4p0X8X226g+ojCwOr9BMt6
aFGRVANJAstxt7+A/bXE/LVQR3tNcW7/NrG/2mGSuUwa+SZoSLLhY/s4xEFkvPAC
csjCLiC5mW/5qpzMyfqWCQycKcjEgUg62hykWmPgBe1jHqlkBpU4bvYY7kTlYEQo
Qdsmsq1ITzv0MXyRE3QqU7RNoV5gKkS7DsfbKs4uHeX5KfJMJJhbOF1K69ksgoB5
kZIH3pQi0cyNaEiQC0JYC8A4fnsyCCi4bEfYKR4I28FX8i4afex1NjQ1BVZp+5Zq
J6lFx35P6AdG/F8F6EmOLa8W/uHGMCWzOrJzGFJCwnGM+kq08Fjj/O5KAOtZDus5
DpxSgg1fB4eXMwdIV8vBV/UAwpdKvV8qFAsm2gJ3NuOOLYfy2aCUZcZCO0/mMN0/
cUV07zWiHa839ZWanUyHoc/NdZ0lZtvP8w6rcizXWOQYiq7bHYnd2c3EO4l2RJYM
Bh1W82Ci6WiY3dSAnBxs5v5h1IpJ5N9P9zSYqBu2FNKGNOFkxswGf/8tHs/A/Y4B
rnFYBo9Qcfug620zFrthjHrqtNW7b9lXphYGP2fLm6+kBDVWkUUJUsffx+W1DETG
vydJGd8iZeNPpaXLvWs9aPz6Xls+tHPj17hO68NsQSluspdsJ8fabWynM/i3ImKu
po5DZDT0N0OjPU5+JgH/Xm6LSqQ8shQnsbZYCMCYO/foWDxBv2uBfdi5DuTioQwS
VcQQy2t7pxbDc1H+2MVt/cCdBeKcVRfIs67hbM2XaANVngKGJzb0yBB7abMF0gYz
0vjz2/Ck/jSUrZRotzIswN4WLGRSdTEFB+8+3kAqYixUpUndmpX1dpLHPp9lRzzm
BLUHuonofSVAu2v7v4TN3O9HVCxKWV+XGlkivM4ea2OBzUvu+fiQ+vlBq/Epd9AT
bHE3H3iDskaiJBtgfASQKYhacjn7gvQw6NByg10cBwB90fO6oTCuBSN3NSQPMm6l
aJJu7CK4KlqfWQHtr8vUoHm2UrIm5hp1C7RscYH9zgYhE56oZMsELpDDjoQBrKQO
+UrXS/rJ7kItqdXunIGrW0hXvUQT7uzgx+FuGX7ZXCba3l06hsERxfurfS6a96kA
QV6H1ajZMXwdczTddnMHLcUVL40IDgsnZWGiO2JFXrPPuzdZk0cZ+NKVGp7x792X
VzBEJyM4eBvWokklgINHai9tA/O/mc8ZEododw0xPQFFtYIvy8fGaT309K7LloUd
WIUVn3Fq4D9oqqrQ+u5jG9CVdF/HwZvgBp16Z5wnvmZKiNpt5lyMB1KQJi7qdjku
cztqQOVpt/Q7oMclGKrgUuAZ5ZW7DvtWWRa7hstGSmsmXZRa/CBC0OEglxv+22DP
W9ibCGe2u6ArveW3kEB7iR6CoglcmqlEqOZejUfbZ7FHt0xrh0fdl9dtSoVmwNIp
7MSdSG830Nwc2uPvQe+1ST7Bno+9SdtnG8hCA+FHUY2KNSW3r2HBApSRAMuKo9yZ
g52TgzkzLhcvhHB55hY84EficsA/dkyCC+KAUdXNZp9NcKSCsyimQxfxVh8pqxZM
3CmmHDudt42Wnq9hvo0R3cUvFi+rnK7J9D2LCa9k9kbwaNnlwJa9r6UQm/MRQRlm
25IzU8hMG5QqrMHU1mhFmkwSJgcrSXBfuYG2Dy0BLF7oRfXMeasEleInyc84ETk9
Kwd0FdvNxLl3Kxda0gEC3DZdy5XkvE/ZsSZV/GKorAqeYvasF0xKV4bn1f157FA/
j2ePmKZkJ1CqJowNI/OMp0PW75rrV5j96TQ8psxvapdcaypMpjCOAMM/tNGTMc1m
2T75pdfWV9/9gCA1Bh4baBgCXoM3fPhh+VQWqjeXVKEMCqrvx2P2eJXf1pP2LY/g
C+IE3f4nRFjlUdS84W7oxqS9UGDwjz+QRL58wEeBpt6gMDPEBBY1I9utJ/8tAeBY
O7g9CTGgT1pRva23W1jn5HsUooAH17oZistP+yimGE1R5hVGFCei73bbfrBJDql1
DxX388uqCb9lpCvuoiOtzuvmHMw0QNSf7FgUHPkcWdlqyf7IKK+z2r6zbI2pqdS9
1yOblRNXJEISkzqb3tpmUHUYrBx0j7UsvcQ0TBlX+1hHt4licC72EdrcCmqaUo6N
w1jjLAM3q62SsTiUA9qvkI3SbxL7czHkEQa1fs1yW8U/dyRuD7u8SmcV/5aCBN8h
yXMRZhoBK7gDFfQjxeQQUG+l0XQhjx9v+/e1bACJvoYd2NwdEba729OwjxTlTEEl
k8MfACfq7iPqLL2i2wPYFF+Q8cXNlAoT3N+9cQKDP+LZH6HUY4zt+pmOL3PZg3lk
4IlmxN7rCe4ylD7EN5XuawU8eXar24hQurw1XbI8L6m75xDS9d1tvJalXMiFX+Jt
bT/4Qj9DSChAPEBbb9qkWeamIutQGQJtINTmWTQ/L3spFg154uupEwN+pMuxLt7p
pcyx0UY3HMxRXBEXRic2iIfzquFZs3EAyaIXbSE0Z3ioR4NT0VfjeKBKlgRVfnh+
pJ8fC27q0J3cT8YFkXpA0Iv4mNRugRX6m1r3IKNxYOSc+m7be0PIYgW5EtgxkPUs
cPVrY0BH04sXwDJSHFngsSi3lVBrgm0pzSACuLlaXE+SKBZJPpbVBijCaVdJwUOT
kjdOVQP8E7t2FygGFxdGyis7jUA6VtP+sPscxPfPBJxhU++RpI6NUP+wkjwfzyvL
Zi9eRXsvc/Jo/NfFlZT2+esGHyfbvqSgcq9DiMh4ZJxJRXKG3DjMLCuUuGre8rxy
/pBkEsJL7kN4OcF11O3yckbi1sH9+ge7zKu6yAjBzPr0ABfj+0YOURqgWgeB2kmt
YAC2NKianZwL9eAXXgU5nTLFCHYu4fbAI8GY+vFjkmygwXSui359cwq1ShEysmyh
yC/Po1k3tCHuExXMYxkbXDLKmCMMyPWVQgwUjUCuXdyx5QOK+ZPbrgLWtYpkv0cn
b8EDG7qVHleBeH9wLk6pMMcWIf7QTZ6Iyh/BlWRjQGRml/QLJfYTJOIYh4FZFn3k
9WZLy3DCWiUxdsSVAH8NcxNGsHnhbWBdV5EIxYfVl/LYzP5uqGG70DJ9tTFOLi3j
QfNCVCRgWET4DAnA6FjKTSp/Kc7xp+sFpP7vdIHVX2NhkXXI3LFwE8W0RS4lJzxf
MAHnp0zMd+e4xoceZankZ/egjSxxvHcuGYpbPoZqYYLdBCc+zGxQX4gWibtbMvaQ
SdfKx+icXpkzQ0PiEZEskPh7Y9veiv/l0VUQul7fQqUmHFfR/GkLCoEfq59jzuMr
MTlJBDJ2Bg6NVvLQsZK+pNOm9ah4aVcdZZPN28adLtdTbATVBYOBauqbe3sEAn6o
qlaDZWbuHXRX9mpFNotja/t3eu8bfFvnIr3zzaEG4tUi1MC6HehzWsBBqWst/7NG
Fpu8JulHFrzCuWJkzkcJ96T6mwwHKRk/y+xmzlclUZRRA1VM1XDyLl2RWYA5q6/C
mr5nBa/sZu9m36ob66/Va8gawo/SdwZ9HBm2TNdoCQJDKDBuMIdMJWNNMtBTAONW
3N4OMn5+1kDZA6VfXheaGRfNvBTnzb4+jBQsYIPjF8Hu3/Tdbm54wq9WmAi1Lz3C
bdT1xX1l7GxCXxagFuQfEWyYytbyKjk/gNL+FgLMN5392LE7rtzddd6LlpWoz7nO
nAd+myXD/mgG7e5ZMtKiqkaCU4m2268HpszN4Acd2BZth7w15mjAX5GL+drRkMwV
mj7X5qss8E/e9pVb3AWjcJ8q5n+zO8rRue3ovcvF+/Of6D4Qe8aUn44LGkbA+xlp
uIlAqIC2m3rQvXbGd+lboC5C+f0gDxLd86wwSh5ODCnInkUXK2NvPXCagycZl6wy
hv4CK/eZYZapyxYAt1ZMD3tDF9KHBL8R9ClnnD9uBYaE2MXL5c+0na0j4BPwhvS5
2SEXBk00cTjGXwQxPo2PBkBkOSGDd/SCbgtOmuCxDqooT82vnx04s7w6b1y1rBFD
uFBkKjuEO7FEjOGb0ku5csgNQV2l21yE67mq/1XeM7+V05x4Uf+EPPb2+iAnw0te
poix2zxpMW6foBCC2G3TvrbzZbnviXZ2E1oZqwOL7DwLgj0HCn1HUZ1dQg9zqvJu
opPE4pGIe9wul2w7N5EvZQLml7OBSZPw3taDIMAwUZGnb4GtoXZRWG3Ai5ETpCml
r+78dH5fqkhKvv6tRL/n67XUa9gq++G45D+oPf7tUBJbKxRt4y6MIcW07lfqrcMe
xNzufmfWGqMMKQHFMPUSo+bLRRmNEpnw4kvhrxBZ+tsPLj4GUy9S+4ly1tyn0NKE
mWCr8jQBNv7QqCa8OmPHArDq4t/V4Guu6nnjxYUmlUPZC9PbGjCI4rke88kSp6gO
vqUMv6oB2vEIH70jzzv5FrGOOr32oYMGHWCn1ioFbO1Hrv7aMRr4t3XqUgK6MB99
K1tzsS0LNnjHqAeNPSsBZq9PzeoMf45VX1aDCdbQQcVD0OkTQY0pJB8ElQx6yKmR
4209tGWUqnAS3uA6gAd15f/6w+2UZtH3mLklabi+TmCT+zBoN3doCaUJQU7W2p/q
JJRikGAzDXyTnwtj1j7i/x5aszcsGVx0uougGu5LorMl/3l+QFfvE4BCHsu6a/40
T1S3//xYMfdUsjMvAXrdAAofUx8rLJfb5nwbE+JSIdC50dUvOkivpS6nKFwipTEx
F51MQ8dv6z02rLImiqm1GZfSB7J4OzWOm4lmZ1D4282ibxLPE2y7XDT0lNXVzDhv
sty0RFT9tQwub+NRsiZgke1cX7HDTiZV7m2uAy6vXKjU5CTneWaEM0uH6Po5sbxd
Dqv6IT8DjbEG+hiX+nBLuJMtddDz5LS5MTR3QtCy/dzAQwu7GjjhbTSwl79Afjsg
SppGLihTBDp+XUmpVMvjCQgAcXqgNqm2hTh3rJOSKzwMecOEUpcAspCOicZiDqeV
WkhfOfk1OS7/TVI3TJVUs+dP1lhvny2taPoEXYvkSlyClt+NlFhYlZhrAVKYYcOI
cCR4Mi0yU87o636Ba6sSRtx/aGEiwQlwshgW+4o6kl8FXB9ccK7u2+RkHfrGOqx2
mEgOzDjzriw8fhOcTw6XSQVx71LbzvSWa3nJBJUl6WYayzrAu0btzhFwJiJNs4fe
54DXFowugGaPZyLCLGME7CerG4woO1DtBNzdQGFwbRMP/Brff3lC+5Okd8GVjJ4N
u5bYg94IXYC9423YYcd7Ukz4QfDvBSfdCkavshhfKGzyPqglIowJ3MopSh5j1zdh
M51RKyi1N36zc3a91O0GxNZusrGwbXCd7t0j+ZHLFf8ALEiQbKavbZufC3lh/4QT
VQ3WKoUCnzoD6XgGdvrZXhr7VdhB+9WbrGJee3zn9WYP2QDyTOREfGIq9Y18eUVy
PGUxWskrC6LSecMegTuAV10vsu3yjjQmO8yw6Do8KUD7FR3WS+1DLuezJzT78bI7
ZO9fTvB1AKbtrTcvRtSRq0gIeevuMF0PZ1tLKzHTuusL6czyosDr8zQRWlHdsGBR
EiqCmCELeLM2GSdEHe0CnSGZmhLTPzI/bZIlhSZVD1XSbdTrjBf/fTDgxdgwdzJF
ewvkO6Po2Qm5vH3uvESyxGZPlp8wKcPXGRvxekNQRQ73RVxbb56KtMiEGFFu2+BP
TnMNDg49mDQzPBJctQ6YaYRv2hE+0bxcU0loj8JDgKAYBKpc/0wsSPlDaiak7M3R
iQ1r1TuRsNwv0gjlDy7xOVI52HDz8oGjffJosG3HfT6UTz+oQrWakwJPf4ur2wO7
cMTyxGfeNom9yYt4sx761WRlzkxnIwTcoleG3xuHo07suEtysQLgcRT6vuUUs6Gq
FJ2ApWCsy6yuwHSqbXhRVpzvLHuI2n03qmT9/jy0mARmA4cuAUJGkrneWIHRWr5q
N6Kb/i1IlOaYIznUpICjlkjkjWT9lxyaMKEdwHaHACzBOyOKIeCESAtqeEG11qcd
vgePlyX7iv7eqbL/ni4DqfKu2ArElY3jBzKwS7aQmbp5GXK7rDJ6FD3zVIniJwRJ
mll09+cf7CsEZZgPJ+leqqcLNNgs49KkAkcWsBkCopTd7/JuYP2h/MtB14i6ZrO0
9fRS+kNRahttX7nttzE34X0qdbrTv4P0eattb5qjDjh+WNsliZfkaFy4jelQXGsh
iBVqAc4E8e8JIR4iirC3DIFW8ZDUVgDGeYwx1viSvlagxxwvqsNk8oQmKOOpMxQ4
/pZmb/iEFzVT2HOyDMLaGAyaW897Bvi8amlKABj+Q6dXrJtFk3UH3in/DOgrTNC6
lncDDsurYhE2Fhkw+Fn3bPOpr7AuT1NMJBt5UK8a0feZ7fdEIhwG1ELjxv2nCK3b
rorbvLi0fbgh3ZQkv05er73DJhfrrlqPn4usQC2H0o40+L80W450WGdwLAMhy3VS
eW1xVYbCParYxKV4sxlggk6Co8v7vh7+RuInMyzlp6zje5hapWbKhKNO9+mNMHaR
T9a3jkihGCQRYM3xcIcQUoHl47v0B9mL57Kxju/N7zpmiRVik0mtowXQTwO1g0AT
tyzeuMM87TlIyt1Bx2oj1Cf5W3NwzLlqWompRZ6rs2F4wfsUI5gIidk2E2zeeKEe
iv6LXZ8QBBHRpLqtSipv3zZ9Kvp8GQ+qkANXr6GmfWy8igr3M+fOdZZg5SeUY+OO
bissgDj0dlSy9VGLFEzn2kC+Lu4tc0tL959mCs8daqpgbO9vdCdCD9YY4KF5Iaw8
6PWxIwe44i6MrSrI/0BDlUkQoLOf+6+Bf1jxCN9mWrRFHU+0R+hvQeQwLkD9H/NO
L3i3bsGO7pmGXAmy8g72HpPyY3iW7zZCzx3Or1cLzYp/QmMXvDC8dkEAmYJQZeB3
rI5qwr3o/rbgZqPGofZesCRYn+hewhFAJN02G9sxE64VBsLNLK0MSe/NhnZL3VPv
sEJ5YEnMxkWEJMdERMVi0KNDs61slh+cOHgXS1qm/sNw1sU74ohZzaopsKxuEZS2
HPS0nZLzNEh8Btk2Z81sPjZj+HtrBULgKn+m+9o7PuaFc89O19O8w342SK0yzBCm
diri4RhcfcGg7VIiraD7zk2l+2RqWfoAtTxwGO7TECO+IzyCGr97TxTTLlLjK2vr
RGGG+wFZkiK2ArjMzeAQRpW6DM1HTcmCw6tOhuDvVXG4b7EAcrngdDiKW7IkaeSG
xvQvyagRhVzxMQ2EaDDZRRWEOD1otbNjJQSQ9MRKrv3G/tFHH9hS00e/VeL6vTRN
f1hU9MM68odC2euwFudKSbUj2++Y858Pqals+6pTh7Hh9sag0/YvN+fzyYqnKV15
Vj7VBrbLonU4K7qlbgOQ4Tr78wnizIAQZYpdcyiwzXCQW6wULY8JBUjRFTON8xhZ
FmKjO0xfDozcer+JQceKkRFVF57RYmPwwl9kzDHoLpsqPFeCdE0tMW7fyvrRU/h4
IW/Jdw/X9142hBcioNyao/eriUSvAdrhyAgqoxBi1d89ExrUSYg3CgFltIrLPTNW
ZFs1UP6hZoBDIu5K+DBsPPBbgbgppfEUeKvUQiBm3fd3mYjpNqo2kl2xYNobwcyd
6emUhMv9+J7Jyrp+T3bomcajRflesQr0k1QZ3b4SFd9PjcTuBSGWmrbI9IE51dmw
tLUAK7vjWvl9gsfZkTvM36l4jSM37g/lPhgLVGnxNB8wf8SIZOq9L8xPIIqM2SCU
xpGtt4CapomSUneHtQA2tap2txHWrdw/FS1+trz2zRU5IDHLViM9CCtS/YcUKA0k
3rPx68H/vQtJ6K5ZiscgTGeteg3OaOIGqQXSw73e3I0gJDCHXc0JX2aKia43Ysl0
Xzb06UGCeWFNN3D4d0aE3Aw/P2xH1Cw3QHaI91Uyu8ZnUGfkmjIoBNi6g/WwPsd2
26JH2q/NI/5R4oeXkoKCeHY3ZEIheP2gmguRwfcbaMJgs0NeA+7kdd0COw0yxVja
kBce2AQdeu5YDQKOp1yLooKq4oSZGuMej8jzNXoI+facwtonbQD77oQwLFKHmX2B
cxWcqAP597+4khQ5AneNWsBGIR4D/EhqiVZ0G2bxpAWbSiSSSfgC9nElbrx6RHTj
w86yYlUXxLL59+LXK2uJzStBfy/mV3tO22s6BnBUvDHMUaupQ6cr9rSG01BG3Lms
/0bUrW3x339yF8e5oCLKBCvU2fBQx/XLrBV6tXy15Fubon1mb9sb4afonrzlLVq4
mop6+7DbHXAkT/7aXw0mH2tGw6Egutc0h14MSDZtmhNMh0iGnAMQ7jZIXQZMmflt
1Cm7S6X68ij35ezoubqXoUmP3Bt+ehtddv88UGG+dDFdW5yV4aoYL1+1UvM+s7OS
v/QUvllU3wEVC9txEce70g9isG5K+UxdwKt1XTFJiBRBRWlI4wyU9F/4KoQDyPmK
Eqt/g8Xd8xORSzjIwOzWvjAV++fRiRULEVcPhHmDpVAIk641sCqnfBiK2f2DFym2
3K3EUSJyxLwiD9kWBC1Kv3ZWsICa5F8HWgOqcI2VRtCb5+sSKpCWIOgLw7qCrk64
OHTA1d6Xlmo4JXT9sik+UaNLuBG3GkIb9cHIbtn3oO7xzTp/gVFAMhAZ71GXwbwL
qcAJxrkcxqPgZpK7Fi0phsSzY8gF87xvgxwi5al/K2jxab6YtztvIKjNcpYRNMPb
uSQnxw68firIWzxz7x/gx6LfS2QnI8IBnl8MWrlIXcM2AsvIiwaqvd5vGmNceoH7
aIn3NXGYHTPkpiM+Sp8J02xHYyLNz3AKQ39VEfxLV2648qwvegigKyjJLiILvTWe
sOZ6fRqNpjx0uU1E/pkSXSAdp7rjt0UBFheEiHlVwosxqwuUt0Ft/F97tehHJGPc
+HX6dYWiFc9I1TCkTt1EHAFEBZYB3tUB7CzAx77dCWo7bx8S7sOWzb9mQ9pE/pIv
4zOJTtKRqqidyKMpiJkGl4KlX3VNnnUpDl622Z5ZZjk/SXtmUDYHcOLe8FJleTYm
PMmF31UZSIh6+SZVxqPVfGSBQ2t7nO4HTvbfamobuQ0dn4ksDrZQRA6OC3Ve0bpL
dkVkd3/T2CUpDvkm/M3CfB/Ehri38vjPd/kNlmf78UeN5OluNEUQnM8WGqWTytlQ
XA/J4tt81n3zBXTO++QUeQksXplIQTHwq1kVeP5SidiKlVggb1K8kaLje3yZtPZP
qibl6HgCkk11i4oO/kDIajpJEHTbdSW8h5EI3Yo8mQWLnibrMS8yNNwhvegvEvpj
kDH9E4agLvAT0D4wxSK6U3YaHIsR3vJ5L/DDLJOQ7wHDWTlAIlgbKD47i2eA2CNj
InAcKwy8Munh0CuCagX1qD1ikSf3IML/RIek1oc2+OSISRW2soJ+EdzAwvOvcTzC
qw7KjrLU6RhMNFg2Qx94aF6p2BQoVNnnaqfo1n1y5zRGiMqknRDmkrtcO+0VOxN6
2cCxF05SlqFJHuqwG2jNCa+pvcGZug1mFRimUoAivM5/72GxfxnWWUfKj0ZhNKS7
jmKZm1bLOTeQ2IiiIRE3jZUMaHuVXsagGXLlSUdbQueS++onkLAfSwhRLjnHPQ9e
cNwgjG8+S1U4J85rP+tRU2zNtCaLyub31550JCpTyenyw2he47fUK0VxK1KSzWgq
1xL+AVAXYlUhNZI0HPtUjWiM46QuK7MT/qkW6nobK2Nb5awSHd7c1XlHGm2++7l3
hbHEJBhKiKm9KijOVlxDHf3JOcmoIY/h+NcENTytnUIeNq43hldkzS9jG05JkOIg
7+pCrA4Tub2Vz/gAatWCocmp9Ttinwvsqnqpcx9DJx/36u+HyGr5Bwl3iKLoGx56
hdVjqknCYSUpUlGbiWMo3KCbW9cIHsftuiC3vl2W8UDlKGJJ9Ai73mJJk3sxzNCV
Z+J5YW1nlO07vu4OCIJJ99hAvaQ8o6wcziea7iqIJ+xMhlIVzxnR+oL05zyV7cdK
hzB2MHfV5HNbBaowOfppRr65s55HVvO/LJw0XYY1A9r1qS3NaffK1xWO7K9VFTSC
VwjI9DUbTQQzU3ulb5XKKGcJCkMAXvyvPx1JF0T1vlsMGhpNAwpg4B1rW4mbDIxK
ngKJ4sUe/9kqDJaeLL5aZRWygVql82CF5TyeEmr23JnI2gXWE2tpR8dQSjjwQODy
jetVmCoS5OpH+xDKF5a/8jkQwKYR8t3mHAonI2D+cfXkrSYu5XKy/A98+760Eh2j
411ghUYpyDAm9Lso9Oe+/E/faSdhHLD455RC0/Cof0F7hUCD0H3XlDNKCdQfNHYt
qedYRksjHMAnhnzfh8cfgJ7CKpX0ZfP9Q9l7cpg6WWjsAgpmRyzsJsej5ZLYSQ+c
l3gymIy8CLlXRVEazCM38B11QuvFWAEaPXrjg6a/m5XukNFgeLN8OE+qiY6uMs+5
Lk3pelaU/tvR23K5HKe+SxbNaicT05UH80RUOCnlKZ80IwQh9oyqotmduRYAAnh9
y+YuxjsnfHm5vxRn5rDmxmnw0JHToDlSKUr7yZm+ZiqJtjpVxmt4+yBFu/bboOHA
hy+GAxickHUZog5WInSlkTrbWedI55cOSIzmGBMSbb8BA7dqbZrXRKcOt5E3lnNa
LMbSba7OqNJ/nHwqHFpu2SCt9bWLfYLFr2snHcTdKL3HgP0PNavdCL1OIaiCISjA
Ho+92h2+kBJKu4eFtZQEEE9tqJaR40jGkFtblu/5WOz6N0OPCycj8ENm6tQbOtZW
VVQd0gx2qryWkB7SGxdXUrwajPKPzRw6ADSOQlnX8EsMOQyiFNJeQpmZA87K6Vfg
8a2yi+iL7G67ou9AN9mmNSIx7W2iSDfOHV0PIL69lkRUDRGJxdFkrRTJUL3fOtW+
QdTBGN+4DPBYGehFJbmCphU044skhs0jP5o2SqyirzP9dPi7MyAMjuoSbVT7Ldsz
tTerBT9MrA+YKF+S8hGWQ/aPNN6RWO0cN3JUh9abrqnpmhIYwky/QnmdxGkj3EYJ
uH4UsctfyAuLfAqhIrU7Gn5c9bjQUG5S0/TaINLNRknsuAk6CusYzrhhkeOpi+WK
cav9fP9Nf+jsfHMZkykDrmKdpwAu8L1Ql3iiE9c5GjNX6+4Z8N3npB3peIoayCqt
u69soLfRFo3up23UH0N5ZicCS5qqYPspDpyoPNBCy9+YAVVbD8WzrivKdtxRbz7q
6vS4u5S46hI+URoQO0SA+tFrGeg+9DgEjnJ7Vv/iBhyZPlRCcovAa8ej+lU7UHQE
ZRzpTnaDs9aCjqTcjS9LEaHZ8cgQTgsMPuEeVvk1mjM18V05kAoXE8WNvhsakFFq
erZ8iyn657piBsVUPjHpL1ytPSCVgkjsqUWw9NbUenGTo4W+4NfJHfoy5Ff5dCni
grFUA3F4lIT/Fx2RDXatFjcb0OF/q+87MkuNRu4wLdBc4/g4V/UQ6fDPahejxoiS
7usrRp+u5orhnxyn4U1x0HKknOYFdlCupc3joVJwWasYa/eyKZofqFKGnC8OsN5H
e6Man0k8YF8fL9iCLB9Cx8vUJ+u/mAri9Uv0ciI1X/QswAaUQfcgkprfFrZMm0CE
OKHnqKD97mn+iCmoypU3ZMcvyYMt7kyK4YelvMO5DbDGvRLlzxAOt2xtO0KQK55R
DkAUx8/PL4XTh+2/bmOfm7vP981eUXZ0gHBg299s32dSZuLTAbPkk4poKlXwvvoA
aAu8aW045rAo7fUEfUrM+NaTzi/wypNK77I1U7a0XJQyb7UKKRJzSJsZq7BEzu89
HzrJ9ETsPl5mxLbwvHN6zrEsfmj0Gwereox1IlArFEYdi/TaROXPi59jwo72OwDf
yxf158OyO2tUCcX9TwApcb0pUXJ6vchDhcP4E9Vt7GKxBnhR6hlk9LdKjUqFmdiD
CjlIhYXdNv5k2emNtRXrU5uFmYl+KFijl/xrQ0QqZ+DuIQKbVDDNT2gc40H9MOd1
XbFEMmJ0mSAwmDHt9gADDybC61o7iGRsjcrMRhEIoF1JNg8iZid05ZBpBudMBnCt
8Rdd2w11FBC37H07UxDd4SbOlscWdzRVNa6cvHyQLcSGPzM4WHFmzavWAbxMAdJ5
9osbKTw1q0A/j6w10LkVpYZzX4Dj6aD9vdxRTS9bp+lKLZq4LuZviZw3Jiaz0t9+
Zui9DLJR252C5j2lpuWj+US6PVsroWx4gSwKKsldOnuPwT8DrVmFFgrzF86METi2
xQV2r41pfx0RMIJjBIDAFUjhWuBtuiyBTzIsZBxCE5O4gWGDtDgsOqeoqKpgFR0U
YL0JMJQpOn+629M0/w8dfXYxpxckqmdPn0e/UzDDaD8s7Z3PasgX8Do3YiAqrZFQ
Fxpy4cR3+qN3i6SiVuesjMGwf7xCXH8vzrFN/u2DIXjZTKEOsK1xT0Ha59y7iWtS
4PE/jLyS97jru35FaeFn9Mz/LCzX3XSmE3h/demt5yh7z04K3O8cnkJRQrid8uJx
Q1worXF5NgiY5Jo1pnidmV2KKTEGQ+JpPfxcz6rTp0PcgwHxaYMxFDg1eVAgLyK7
NDy4kqFBlUFYfx+9InOyjvsoKhJ/AiwHeM8YkWeb4eIVJgxtNP9HRTogV8MlHqZh
vfxJRi42vwG7a4LU9yYQXem9A5oBRt11MHpxVPwTRo5KF6TWxAJsbzEzvupWFlei
wAebO5lN7ER/eQBrJ6R5gKyL/E0gxTihJBni8hColVt+5axSRQnHZl/QfmcceQru
N8CRkVYkXMZPAKC+EpqD2hpbBQLPXzU3MOzDhGS2XgTqdxOl2JMpwBFfEqgh6Xb+
sC7pz/64GIPDVkYnzlhR4FPXFyGhtsWFttvBIznd4t/JgwVrCbjIW1y1bz9BfJkY
eHNGxSZKXIANqiGDxW5GCFp96veegxEW09cJg/eUwtktm53wxSVSRC6i5Ys6jCrR
h6Mbe/W0C+MYOxpOFIfdToowl3mK1OTmJGk9NkdQCCYnT7DGmnojjiK+nN8WvuYS
+ZTrycptx4907xRxsmehbNunrtmpA9A6wpHOZo4y1vSYvww5vrNkw2qTgY/kkDLm
fwfurf2mHavzIMIlhX/S1M+6ckCkT+y99W4Gm6AEq+WhUBXGxy92Ew/a2gJn3PDd
RnMFJwCTvxZW4d1ED2PyzXGX7/dugVvjAHs+fgXb47e0XwPAmHanQV1gR2QWp7BS
AGpKHTOheeZYtVMp8LoqndZdsmc9PmeWhM/117tUxQuujj3HRDXTD7PaW8zX7/2r
jWDZIfi1EG9HAafIIPLNV4wPuNGKF6A4uM9F6IzryBfZ5QiMjOIoqhAVCMc6mCIX
R8nEsV9nTFeMTkJwEGH87OHRV9GLxZBqmiOCL+iZFcV9oAUmjDcSjR/4cYqdviM4
1iUp+xT367MtG5ZrX8duB/zdWXAed/rCr54W7gbeVlSB3Vl9Do+XvFkWLknazjjH
Z98TWrqD0i2XB+ce+utdO0oC+ABSgRXvuFSF1Q3Er+E3RsAuq21V5eHAKYG2e9G6
B0bBPvG4LUIbM64l694p1HQYxjydUTYHDLM6jW1/dBX8m02x7HE3DqOCZDVe4mUM
SgFNOoRx4oLObaxest94oQVJ26s9usd3o90z8J0bA45EcCi33A0O51iZtAkKDYv6
RNXlA29j9WSW7OgsCqTpZrLEqX4+rCrPth+Y/BHZRWOCpMx7ni4YVFbvrEjWauUa
47h5uqs221tFKsJ0jRnc4zT+vTWmLDNWgeL0PHibauT4g8NQTEQGaT0akVS447Mt
BZQFrDav/OBbTnYyY+qdBuui2kYCdWI/8xFiJJ4DRvv5VSiIhR9dXn3pfqzDWkxK
QOOStPeFlcAEACORSNm/LRY3B7ZxaPYNtjHcfTGEB1ecdSrvp3bv/7Ii+4nBvrgU
wBTf6T9W6Vj+mzdasYqQ5myc0CRr2Zd5KmeXAkBBUPgpfUJiY4A2aDkj4wG0nnS6
2m/kQ0i7DDEBNaXgAZXOsrY6PfjxJu9bU9stwcdw7EW7f1eQ01Oxrc5H0H88tJ8i
dnKgLAKGScxNpX05ux5Tab1hhhsAlGJn9ISYuDdyv9QJM/p4TdjWp+z6b8yVtdgB
DH1IlyTZi2xkilwqi957Oox+wHdgfL2o83wlCHxzkiaKiwR2kkEHchnQHyFZVcg7
kQ6Yd/ho+NbgJ46F2j4AYulH1lPuRFvDobIdSL53Z5ChuCiPI4gt2IPx4n7qX8LM
+pVNM1dV/MH3quzDqTfajJIOTqRTF85TJxFbjNwjJwTui7vfoynxdF+lQfYtmpHS
VZFpV3qaQrWRAsUw/iPx6XGrbPMUv6zxZFajNSL5OPw8PKskV5ly3QUPPfwX4nPS
x8GgpkHMBR+jciWlVBriWxOcmx83YM7yEnYk9j7HGQT7dFTkYbt1NIzrpmJWEmuY
aTlEL2BEly5mJTIOS9LtqBTpGpfAWoiSjv1mPNFxjtwsrm59/xLY709MlFvPtj8n
KI8HxQH+ku2+uQomleI9BI8mHHQK1jEZXOl9vppv1FPx/UsoBMNaiHfagmuiJ8Kq
nT824HEh88j5+S2aBcryYeXm9KdMf0sXj8n3kr99QjW1BiZVw3dHFJ7sXZfVLcG+
VGd2JpdUKQu++9pKSNZ5oHnmDQSkJY+ny/hkJobpLXsAhr82IGRGyCulO0B3Sg5d
Wyb4gf7HEPN4wfGPsyGnTOIWLrfXyyp5kSObMNVu6iqFCDiQ6b2gOcN2FXsif+sx
u0ppvtT1IAuC+JcFCAOT3nGYdSZmZiB3gFP1NQ7+0mORndKtCpriKN2AE6PjU2JV
oMbWiUReUyhPS8Y+J2DkFRwtyUgZrIM2+8gmDdzywQBvrRBFsJFl7sk63cXWRCqy
ouInpZoN2YNcj1MFKcK3xKgj30EkE5Q1PHCgaGHmL99kEq+WfpLJJU4HjAlUlhEX
502PVjMVA94HgEAHJoh7t9LO65vqQWqXBVJBhvZph2BxpRykWEhuJmqdJuRw5/DI
bQdNwiedgeY4htaePaHwa65BDCas9vVpWqvl1acTSMmRdM7jD+wwUOo88Xye2Cbm
v8bwAGJwaELUVeYQ7eU0iPvMnXJ5MKCMOVFGS4uf7sm0PimjDIn/3mFYQcgRheYs
ZZhunmAiJFQUwSVz2KH5weDFjkHG8oCMLJ2DSQZXJ0lfbc4z+8K7k6DngLJbRSAq
wZErylOA+zR7Ojc3WUoCT+rV5XgNjI60G1Y+3QpX8B5JnrO+NYglAD2ZP6fErA3u
/t2U01du7p+2bRVT/lRE3pV7dCuMo68xNiM4Gp6MGjIffItNzP8Zm0NV5fJhmWgf
jnJLgE9pLuq+4ObGd3E1jg3avCOBtbJrpldBk4Bgef0wNRnDUGZ0nv4khrWXLWsY
oHPOYAtyF6RGBv4tJPuwbd9e9jwMgqR4YjGptMQqkNEQoaGlcPxFBpKOeIH+pJ4P
uIUpD6nftgHnljlf/2mp8bLkKcfVBNIRogt4PrR9Xp2XNRyMGJ3Ry2fjOlhGBp+Y
AesEkWTF9PaOsZTygSOyXyLD2r9rNABxpiOTS4GLPuMbOzqI2uNCN+VvD1Gaqq+B
DN6gONHRRO0iT7NBGmpFAaVbsoGgK18vozRG1Vv2/C2S+ZVWppJgqPYZHagqioaf
1DsPx0W68p/qpdep91j86NCTAy8bwhGkl/+yycNhyqufLbSAmYbo6p+bqvl2l2lw
FnyIkh2NnMfHuyrmPlBtOkfRk7Gr2LNykONINMJwdc6MmgadkPxqBRwp3p1e3sAv
RgT2VBTqXvZmLA7o1twQ68/HEfijIxxVFlnqv0qPa3xXaOW9AJh2bNXlgbBKrjgs
pJX9EcF47eDI8ZagOASltq+eu7ozSo8iM2sR6pFpboAhD2Jnx7QwVXe4qdgsDk7S
GosKj9qR8SlJ2ZXeZpvtMvF2ZSz/7/drru95tSgnBAfBdJC77T0Ir9gUzzR2pXoN
YtIuGzrpQ3zNT0jNSwc19dblFxuE1vJfaPl+MltjfhqmS3avk3PqWjNKOzefauRt
t2+P4sW4Sjd/GFbA/j+QxrCegHDM1V/hYKY4H+y6xtMVr8KlzOm5ZrGJUNdrDplU
c4l+LVjHrz4lTxcSt/oUB58mt3i91XtaqmQ8Hw10fNcwGsmHSRQX3ayxI1XzMp3C
o1P3lKVGEZsAzn5FRYBYEv3dYt1VhDxv4P8UMAiPlxke6Tb6mTo/8mUb4ZvuYgKe
Ue3ilDWlB1izz+8cRjf+S34gBPtHP+qih9SGViDbKTumLSCWvwpW8PUHM7PznB8d
8E8LjVPucO/Vd2pCjRcnUWw4G8hHBGfuv+o3/8OeAuir2s3XzFem/jTL7v58iKa7
V7cNS8bZK0SKeAmDygOQhcm0ovh/hxk6eJK5QTs7APiNI7ZEVQi845T/hWDLRhW+
sguXbmtn2JxKiyYPd0x21nRvWKyzXazNfUT+dt+3XxhAa9IwOXkI8V8uaxV3PRq6
ZfnaEtJsMXtzAFMkPD3gR6Mc5SN1ke5nIS9lQUtqIzhXJ4LZsgix/Rl/yAmZsxtp
lRYsJhoA0DiH3ZgNfonjutdEAG7npqnYusnnonx0bEbz/u1cWkpKDevtyqeuALI3
0sIXFPxOa1u8s4g4yrHncR20xh0AuQ6nIJDDABSuSv3iOm5PLxb3r78m7Qc8H61N
b+OvEZIioaF7qtCTdJ9L8o2CPezsEC6Q42GMuRJNtB/zYhiXcanbQZi4LbRSnQfq
3p+Oudd2p04nHykxEmfyHDk8owlXyBqSgANy3w6HUEPtfclkndHagLeqPLW3FVEH
rZVX+zxAiEUIFM2UMbpl1GEp9ixauZZmL/CtZjtVML1I900UstLqzRaRQi8Og3f+
0KNP0QZmCcoKJXwuI3UqEXPSj1VWxiTyfeeTTbGMmZQUk9Bde2gSA6z6vxVChRFj
usv6F87T6CC3yxLoDI9VBv8aaXRW7/Y02DJU3tANKx4dywhYy9ijxHUoXIccuWKh
rrqPE+dDAI0oGYYbf5gthLZNxM8oztdG8UcXRPj9ZOh7QQqSuuY0EzL6W8f3L0Au
spp1m6rhB6X7VuZuO1r4O3lvmg24rYfsCPtE9fDh2H2FPiBkeO1UY+B09gSdaHas
tXoC7H7XA+dfKwesclpoAZm3dDElCIGKbMse9CtOBUq03RpUyQ6CZ10VAHT7uen/
fXWAbtn9i9qQ8bfM+qrKH02aasb6OP88o+a2TeJjOj1jnxt2NvhNrEU/HepYpunB
CdfPTooTbMyW4j6FtrHCHqUQ3qQQz04mMAPrW7MZVY16v9AYXk9HYyXhmGSuDiGs
lK7zQBdnpMe0rDZJmsBgxhuoq8kEKu6fSWv0KccJXcABr4CQQxogqlnUyvokalzU
BKuSH/tY989MtSYuzOPUv2ezNZ4asytEiScyjlvPJzdL9PyhNJFm+P97ihDaf1Gs
nDr6Ltiyn4cbvF3ckZPjLVFxwA/OZAc93wE4qb4BwY81XLkGiJq+HWVofjpOg7nO
GHCpN898KLu/JfW8e3Ji+94HFvIIOF+kBBunLWPC1qIDq2gq/URcvIWOPhZRuAgV
UN4Ob27ONjXqivpNR5r3JVdf1NdmmHKynknu9GHhEKb7kqfFLyfFj/KUS7IqJfWf
lj4nnESCV0cAYHfD6QNMdueovJ0DyLG8o1i4+bEyYVgNJXWbaS4t9DeYdknpsC+Q
NSVWnOGVVr5TXuU6A0uPlQzGtDBV+LbaLgTi8qVPcoBS02FDAW19D9pV+cfp0mD2
t6Hg5COlJ7DtH+vV5Jid4OfIOzgxkJDZXFw+iF1arIbfJZb9bWgDNmGSbxrkLvFG
j5Kz1Ha9wFSz+OVcE4RwZUqKhtB+K06xnfXHStJSsTiVGS29i/J/JK9DyL704KSf
SBiern8onyulgoAveB4V3uNoIN5heMQyuhnzr4rhs7fH6Fb7feFnIVcN5ldXH8a7
GRX8G2DMxGbibwUqYJLAPlE7sIxOtSqXR5zXjLM1ZAMm3+m6pTYU6lsknqCHddM7
vTTu1U1GhXfcTC8jrEPpJ62F8WTfNiCKELHvVw/L8ZcMYrhnoFVs4EkI3djW8vmq
U39SQ+9kjif/JQsvbZ2BnT/UbY0htv/3Bj7ZZ6KD0XPkhsFDArmcKa7GzxXwGZvC
5y+iBHzy0fsCyWI6WKGw80iSulSsJfFnbcolp4ibt7fUR1Nb9KLQDK3qv7KHRAcB
fBaRkOfmgEHDXfNDTthK5kCe3pGY7NH42JnwAzREYG6nPHgF3bl58ge7/2QwkZTg
XuTI3Iu4PEenfrFFtqr1VV27/qiT/2/2UkyYSveH1km8M4yk5a64mMNFVzmjaZo2
Cp2eRmSlnKjQKNFS5ZOv/fi+ZBCWUcO6X5pdrhlqvcFXurIxZmmJJR9xsp8UhJyE
w3Obsq0LroYAzSXs9zQgYDXETN/Qj9ozrbiwbPDyRX+iz67KcTtvaMbzC5RHc0+d
YCsdJh6F/6uK/tTatbWd1t6X5vWKitPZFILpkRLN7xCCSQZnch6j5BS1Q0OVk4P7
puDkgY/onUdD+ke0lM7O51pD2/BCqHQ9RUcobk6VYHOaOYVVQN+zzp1EnrsghcwO
DjKdybTxb8HP3oAKkJ78BOL3u0Be2aYcYjL+h7ZGsUe+F7Xay5vIG6NoyjgOtPnF
SU2R8fuIr5uoS1YktiaSyo9REpwMZqKhpe0MA3EsjfGBOG1QuZUCZT4N6aQ7Tett
ZHvT2pG02t8hUSc4jPUAQvxEuK1FokHOw7DqwvCdDEClKaqatUpc2T4NhMKJAZEV
cSRNucG4FV1EWiW16z46SEVTNwTQ3FUE8ECrpe+y72fOGVgnM7shYxCzQPq7nyUb
J8ls6k4+S1uRA8Jm+/vbyqFH5hAmQ2pXvcFQoGAvvr0yKTpelq4M8K0DuLFfVkod
ygFLE0cwTQ6fVLoENlmsGHK8Vx3ig+YpDR7c+x5jM1hYece5TE4OFmjDbXSg15kh
G7XwD7v40j+466sBhuqgd5gWNAR2m1c1EiHWrY653lxsHSVEUJvlIIqw8HmB3X7n
INAcPBcmnEVQB65Q2HeYlV/yqMY0jFbPOt9KqU9srP4td0LvIcIYSLIrk3LMFTA3
KVP3DQvXRBMAA3TZDBEXbZHPELN+cHGpJuFIbO6DqnhDJhszVgLjd9FtOZVF2I/S
RltmRZ7X5A3g1eHhrwqMgj8BzeVSw5/yFQaX/jeGeMwFrgVfkssQJ3uFE2QY7qNn
T8iBwSrI3nVOcwQVufAycLgriq9rSgwTxdzvJSuhf+9qA2ut1da5bZGolwsizH/5
Odt3Q8sY5YtuCn35HOFzgbt7IdTZKtJ+LLfbCeTtDghAzZ9ijSjFV8qZ2CpPryQD
w8AjpmSODuL3hhgZQLgLUiS3xIUnhQVYWV7J1xCEIDG9EzEJ7R/neAuax4QiaFgV
k6Wkzd5N8Z+RVjoDuC1KKOvg7iaLHkmrLhx4GCxI6+y7cNV9r/lOvZK7XPtFk0Vn
k89rXGBqnOzlPOd36dr1St51/fbl7yBsX+MRAri5XgDEUGafTEWw8DhchhlQWRRB
MCsNsgEI/vStM/zfcxzqTr3ILRoe5qTtX8TkQ34Aqkp1M5E17/wYEYGWsdQxgx4U
MILoVKszs/3wyJ+mmFoBW8bxlLT3RRREhGJtABF8ew5rBi6LAyOZtM/0je/tH220
kS7z/YIOtlO9siK93oIQkTupcycE0ekOF2E7UuV0gyTetopGkP5XVk7s1sJJHk87
06/Q8doC39WxY1sFK3Qtgv6EnsP6UxeU3VX6YV2uKQgS92dkhiyUK/VfzsloJYI2
qqs8QYyMdzcgcappzy++kgV5jpXwXENuuTOoUGG6H6ThOIgS6rVB+jdCUAdqrSit
Xx2rbEoO0rATuE/VgtJPfV3b5+g6aqbDUdy29HhhgqP2v8TEM/mbTPE52ywp0i9F
0OqU7QEBi7hWSAO4T2BhughRDYcg5RZP/FP3THl6S9FNmcxG7fwXbxmm7HlEY3Bm
sDSeuD+gnbyxbL5EKdRGtz8qctY6bgCrcNldRF+K63GerH2TIsSROwdY9p9DlQ3w
+1jJ1xkcc5V9gnvf0t5mCZ4OethDp3W6Inua6zbdLy3YeL62DJhlnnQjXOo15az8
MArGDXoW0rrU9kaeBK2Vr4cf+mf1G7ZsgTNRSCkhshyShhmopVixMyVRWS6SdfC+
0LXWJOYe8cjHaEciEpyrwBq1wfyy9G6VUzPga4iCllT58nwHSpWWQWoS6Pi/78LJ
Bk5VMQZJnTIzSVAFzMyIILHlQdX3K3bNw3fvQcbhE0uCjsVd5KANXy4qvRsWiKyp
iaMOkK9vXtoocrMp1+Y/hsCoI63i7kRHL076+Diu8Fr28phrqbmGvrQN0saKaX/Z
dzx6akTReizNIjdiUgFkBV5F4TmL2Mg9OPp+Dj3SgmzkejX6y4w48IM4Omeqr3by
SOY6BIAOP+KMOwHL37y03tJhdgPBpAjCcYOsRo2yfb7M4lbcqDZYEKqGbXdL7VPr
t4bJBWJZtRmiFFWOeEUHofAi+D8nZSGjh/uvdwhuK+di0cVQVhodaLG9tf5y1gzp
NTpQamu7eW/nMjlrz5MT7CVBUa6pd/ePkFiJw/iCc9vZJ5z8BFekMtJ+QEoJv0Zw
vo5Bo2qZOqQ+6kHZK8lXd30UX9yuYiLDSaNhtE4vOyzpjxXSwIP8TAxUbnUgDFts
ysv10YdhOfX9plzwA8VZBC2oR1NHK+gluZkDY85EMJ68Wi0dQc1CnHqdamejVRe9
uqno4rQqcix6d5OPF4hUHxNO5GvhQFK+Nit/M+ATgJvvlSqJdk7YXDbFMt9zbIUn
P2qpoKtJ7tRmDW5r1JL3p932pf+w/A9puobR1cth1nIH0xE0uVFrx5HgzEJHrdG/
toCk5VzebzJmLaB3BapoSMNwEdbFwQufE/vDjD5Xx9Ejwhqxal/UqnLLV/guCciy
vNiccepuoBZDQ/b+Ogsb9F5HKH2yY2aB4k3j8QzIwnJI0Pyg9Bnu0rhEWpJCKypQ
VhvmjndnP7DMszwgETxMnRnph09FOBfQ6w4o6+BT5IyGpN2pCWdbKf92yNqrT/bI
R/6QXgPe5QqGdH7pTMf45wuT6OxozsMxVER8fCb3HgaH7+tRlYn74CG0EiuJqQAG
H3+UhXwMgF2O5N/KNnMtp1tkB0DA2ASA1/XGp2Y7Fu5Y0tjTk4HUFAms7LIpHn4x
CR7sesJng9Cb6sSYPI1w4ZkZ1YzY16OXGvGL4W6SmCeUKKCzz+xM73+w1V8OIofb
v8ZEn13ukLvPTWkdnTm1TVfeBg+Aw7z8OixySbOMRZjzoVjFWg5KNJnP+68/wWeh
kUBNM0SIG0nMzGWUm9v/4efp97mfIPtMW/hFwD7V1xEN/FrlLc678DyS2KJZFQFa
A8XzFFkip2fMGhTTccsXx5aTifbtAYScwvNGQ6NhGTfVHNcZ8IdCx6LT5X8IhJys
NYMsJBPGPUp/Sm8VK4XqDVufI1tRmknzVhQsJMPLyfy33M1NZu7W5D1e2QTNFCNM
DNisl+R19u92/nI8CDVQ5IA7wrufk0YMq2jON8E3mXw1nC0Hy9tPXDJ1atB9zQ1T
nXFL041B5fOKZmgMYxrnwU5KSD4aQ7edyZR5SKcAK4CM1yjHhB7K4IEdjM2ZhjPO
qMRPZFdz4N21XLsRsCAKbE3E5yPrd7BLhERmAXW19gMqABr+JJSyz630EFMUpJcf
VOskpBET7C1nFBjDQsGMK2tMjrXEOz7a9Ht0hWFBx65ccv6+e04RohQuc1dTQm7f
OctoqugC7ug+Dr8S/dNRiihGDkkun42LMeUcJlBgkJI1dtEoPlkG8Fe5hW+uc/fV
mxxLeR7gznfqxRQobLGqHyfIczgCle+fgQALTmxlBh2hpV4EFLmIvVPupsE2VT0S
ZYXsObdSlgCEcSmbMH/ym0+v9kMfAzna60oP59coKex/XFOQeWSa0e+d0jl/ae66
Iv955sTVJsfOTg0tlZbgpZ3wrsWBhxlrPCOf9fzvy6ekHVWu7nSDnGVjchzHWxkb
cJgx7kgl8iz8BtuBblfz6uVOT0yU46AsRrFh/hgFxO5LUS0FBS9jeDvE1aj9LYkX
vyWlXEZGkLaub0Jl9QGEg7GjEgKPWbsHq2aMVljHdiyXvyYtoyzZ2vpxqYZHnWuw
4TT51jYr+4pocf9ben3dIYdrcmaCFeY0ppqjjjmx697L7cIIMw2YgiOkcjW7AinF
dvi34Vin9Zi1jX3SfOueiUMXA0V5ndyPswjjSqnkifLeGTfc5cCRQVQneqhKd6tl
v8+LSDxYLPx96XYg+iZEuc2DajADnuspYdi6/fT5mK4MxwF8C8RccE9Ad02V99Sk
koeuzFyG4lfl86WXHy2PPzgopoqEPRXBN0PA8JjMm7nWZJ0SNiqv90xSSnXomAnk
uowQ3oZW2habAOyi0wWQ33gC0a4QcnM4+pGckpB6HgYQQRQ8fJtJ9hNYC+Le28om
Mv/i/tHDQcJoOSYGy7HwTA4R6XW41ZDmJc/ScjIrpZCpUd+Yvsg2qkdBmIkrgoPF
MSRn/mZBg7nePZ7evj6kuldjhfC5r4n0poO2F47J1A3q3CilHInze91fQ4B6+glQ
157prd33LzOyV7lprwbRXWw6Aq44bCbnlibJdouwTreIh6IJJ8+WT5BMZ46VDHu9
fUcGscVC5KiaVdbyGj/lxA2skiOTlqVJnrPt08BwfzmeLnWmNZnsAPSlpyc5O+8s
Myj3gJwU/UyrtYxfKGTJzoD3w5r/uXr7BGhvPpHADKxSS9PJMbIy+nu9CCmo0SFM
CyO23q1p/hARwKndOpVcme+TxDWe7niLsZwGm0Rw7b8gAjo5ggfmdbzpNDX51rdV
HW1l5orsjVPLeJgHz4K1FT1acipZ0SlwHV9JVYJza8Rk8ohmJ6TUbwQk4q8fJqJ8
pHD1SbKE2rbtnEMc5fIzk7eJ2LBfrbMtanvqqwMScxfJJkaRu8MZQVMNrQdwp8i+
KQnbbALgrbmgSg+zkBSyOG3UW+RPq/K2z/uMJeIAXxieV5yK5PLGnpd6DSeKCi/o
cTQx1l465039JSboYV825QaIvP/yYlz+3ZiqewCvmu28bIpOf0d+8ceqFBUKwmZo
w3673D7SzT740qQ5+F7CX+/csKhH/zhfweqEmTwnAqrTueXil9M5ynZjU0jfgPVz
Ro8Tbwpgcj4/rJuoz1GCMGOmatJj3jIBow+gQKWWJ+Bm0BguvK/p1IsQFxfcmBQG
vX09BjP5CzyABrWmSUozlF4iT7CWDPOYQ/l7Uy5hWruPOOOZRkhY08Y4ShJryk8Z
6/65JYkLRiJlIF1Z9r7knFw6b1Zf6eEGr/l2WtKdjTiynNcVO46RM4fkcAdQNSlX
xT+hfTessqhmKyP1oDzENAKzoU3lmJ/uxQGMen4stsZXXX6OknWE2gkt9PedKBo4
us6jYer9i/nXg4bs1lE0j30WdqmEzqYp9MuMrY+0sl+/Vp3eweWSEIoRHLmFMWM8
DAj9S3kZmfA41lG3eeV6+Pr7ZCQqGi3p5IYM4KsqNZHTESEEOYffSB5fP3GgoQXY
j/1oTff0bzwW00lvpSyFOGZ/jBrpD6biUGBQVnt1hxnjUIjzLPoSPp3eesZCLgQJ
mPifuboPunk7idswwHv8rooqeWQmvXvRy9+QyCGzMJUmtVIk22v8YuVdhFj+LG8j
NYn6zhwTIS73NPO5rgiyzUC42ZfJF9PYNzIAHhtcso+95ukJr0JdDXT8GRV6zfh9
3JkD747AZKIrXY6PBQ8f/DVftC2jfP6vrAeGyOb6bpJTzehT/77hHs8L+bh16XjS
FQA1c38NxKe8bC4Z5IVvAXamdvKYib+diGu1WyiWWJcvyeyhg/85Sq1OtGvlbV/9
wl88ILwR6/wMhWOrPl4crW8qoFjHxkFJ7uKyx5ikIKn9FbO7UWdgLhDp09+ru3cJ
iPruVUlHtLPhpKv71gca8RW2DgP5R5NiVQx/RCQ2Bal6M6mjvjJbB4B3q2D71uPb
ObeE5Jx0rE3FkrL4byRlfHN/1EXAT4qk3KwO1aDdf7EA5OXOQMgQozTe6fU9zHrT
yqiUnJTt7/lBRcy5IFATxRKngjLM+PqOolDaaCKtB3GvY/7nYmsqj/lgcLDdYSSX
Tna/bKK+UDYyOrLVMNS+MXSB9UNnh9khVTq9xCio0owZ2IsMR1xU+rbkc0vKcxGr
VWkihCL+3uxw0EgmW36ihb6oT3rJZFya2lsU6Ei/NRu4x/ISoFPPVhYKTygnoSpL
fEQrEIzJqkzm3G5tOJPtjaZBpfL1DPZ9LILe2P7gkB3ZSxFlbfJn8dMSvK3cFUhV
mWOVOYf9sHtsSzKf45/UAm5J9TtxVnMIUHAJk8nPI9jTpasyHI+hrjQd4BRBAe2W
ZbNJhuk+1CXJ2opJgshkvQTmj9cyNODZWh7goZ0gq8cYyG/ZykW7X5SZCGU6ODRn
RBaWH6820+8JioHLl5xTmgDcT03sWj9t9z1WQ9sVdGiJsVKPzuXnmMTCFGA7FAHm
JZB4KwjgWI74M5zNXJCoqPr5ZilI1ed5fVbhf1NgsIr+8clnOB8wmBxqOo9rkykM
3gWevS54JoblUGDfT25c6LOc1IIqs1IceR9h4PaG8osLdkSrh+xnVitqacQTHslF
y+KJXH34YR502HGB/1seA4Xx3IGfjV9ghEK1lGW4ncKTZHIRsEZArxTmmB0HFqrY
JUvHf4YO6j/iSTURG2uLglvN9lOiYnolBxmz3WKOYT1Ss9S6RSNr7fyWs2oaW9ES
71MNpMgvcqWXkEnKLQyeKbz6OAT62pw1v5DRgeVoOdfudKD1JJtfQrrToJI3pfTo
KC1bab63NuYgnXvpDx55uxSS/bDjOx6DfMOqgLdrmMRRiCUooNbV/Zkjf4FSzZBp
v3ATkI8ow6NvkiouT7st/BnLTudLMxTmxN60dRN3z6YfYocvjZCEcy3k07xX0CK3
leTEYwRXBjD8CvZeHqFxcwXB+vmTWHkUtSkB79GpD/1etgkD19nTj4zpSL9Ee5US
0H5M83HtGBMSRBgFGOrcJHUM2j+Gb2d6P2RqMNrjjnLcOsnLMuUZWuERz0/zpWs+
j8Rr2rEbJJwDMo4yf2naDgTQpLJR+f/sZEcW9olkpJT6soTPrMGAo4iPioZZFWeH
RKgSZiU4Oyq3cH0qLPi711EKifW92TiP9fooqQzYBx2edUkNbGZi9CnSMfJalL1G
X4uyh56RaeX8xRNuLcgqn3w28J0a/IK4bHHQnKhSDPAev6zPSm4K2QcFyF5L4Y8E
2SXgA0UjsUzuGO6ZiXXJ5uKhKv65fodhezEcClfIQSEnKMZXwGKDGHHvAsjQukr+
3nyUXvZCyqR1QzteyWg7uoO8a/tFv2yXnKtsy5G8I2qqg4zxYMQ6f0r+z7LasBSQ
NgXSf4NZzCUtII9ec3x7Uj0irGJ1sstsE5sM6hQcxMkkEKJ0Z0lnHsKTu52aDqLy
fWLlx5S3/ukeZtSGvP6m0xIXdn9Kf4408EtruOtXTsJsKVkMNmnjeTrMoql4sq2B
oOyppKbZsy1BR70ZkFEborm7SC9DIKjimYFS+puJBCOeyg+R/oN4kJEmzz1h+h57
fnq3rNTR2ZFgvj1uN8NRB4rL8S31LFInCh2oM0DXWPNX1H5ao/nk0MCNubV2R8VK
YeK7dVkH3w5swweFAUAA/vDpJ5FJ2wVPedbSwGFi+/z66uCMKeRuULvFSNl6xZFY
qbLJm3IBSHksaHeeQc16qjYnF7XVnz614KKNh6u6OWYzjw9Vl/5ShsX+PzITD5ei
wYewoJorgtW0xjs7Mnlfu+4rmIlYlizezrkoV2Dl96GK3bnOw8V6dLKJow1YpriW
WnVOC+64LlZURKPUH6zpm0U/WVZZvxYJvivDcNN+/VARFWr+5isUqmOcL3MwXQ+U
9MT5KGIy15UZLfW4avr1s0NWF5nzc+JsImkvvL1fG47sB5And84u8RKQXK63DKSi
Ek2P+BVHGeMrrUc6HbKjCzfulAwDCb2/9BClkqrF0P8Kxpjr8qe1fBjdiC59f9yF
Z1m0qJoQuLkQxkPRApJXpcp8zSdUIwkKzcdWw/e/vdHy+R+MIJoVUw/u5nlvnxf7
MTj/10BFkDrP/U4VLvExYl0hA+If//hlZvc4ydC3TpxEYcTreT1rj+8ZmJFobR+i
5Eu2useFervTrkCdbjvDiPBXFnoSyFIDMScSI2HQVfInUdMaDmnfiiP1PSB+DBi1
H7Sbq5iqjndGIDHAGc6H1RkvkaWOwL8a9cr1r3+kSbNbfjlNv2wvX1ncob2Te22s
1oZcqAvFdvsHcp/mGLGUeW5TtnvMrl8zf2OMqcEpNW7/ZhV9p4iIOeBYvSNnfx3r
AAybB56l5O/oAr+6ldO6FRFivkx+Q1w7QJrbg05fxnecE9PjbajOmC1+ZCilPrrC
6OytmgxY5jIdFGzAaTyxo8aVxJugnvB+Dp6IYTBauML2kJJ3SiZtdpRpRrWG1vjj
gwPxgwigLVIOKZ8wvQjM5Z50qPLUsfmQUwOgbvS4S0YeoKnlRpaxsXl9732HxYuM
3TXZgZZz94UUdS09ZBlbUzofasvNwHJXNODtlfwWSPQTdvSVn3zH0vkIQBHuFdxv
SAuxbuqu/wFBYq34tTy4OFw8GaQL9GtKQUWUJeaze6ZOPQvmvvOJOyr8mdwbfCk/
pgdb6eZE8wJefAx2f6jIpXdqO1P2aaUiFd1n1NGxCvwsSa6g13yazIDfcu54xo/W
dn8Aa5HyxoYhGW/f2dvSOhy2ssXIWyJEpr09PdY9sZtYpH8wvT1LQp69S/26+i15
IWBI+4S5PmDLXVMN1gX0D9fDe1ZhZlWOg1OfC7+FTT4n1Y6aT42XuBr65j2c14tp
3VQE3qrgP9NNGHk8e4zJLDCZl2PuJKiXy1pp6sD04XngpjYlErHpbnEOnRUS6Tur
X1asCcA45U/6jFvI/pWYF9kudL9NhIFpO7umBm2M8SxkISeoQNtz0w8kRKTYPc41
mwOez31xkE02uevJUa1zk4CgzfDz2LmNR3uqCAS4D63QTWbT9UECWnMfMnECpKM5
lASnzooiagELEe8u1NQlmLijjj9ZBAIDAqQ7cO2ZdsgJt7mdF5i/tYYR4bUwHDyb
0YW6znn2U4BWDGiltNAhKoQshL/umccy0gpc1bAsyHsBMZ01NxJXTlUZhdx5UON3
6EFmEii6M8Bp9na1N38Ekzc7U0O8rmve2y27CEiEBhaQHWSTdsGNtFsX9RHi7LaH
HqP6Xz10Dv3NGGfDs29vPnzpY+YHNjAsN+bHQzPRNbm//B3vM4TIexRw/y0O3uHg
AOwywK9iC0Tjn/SZd94817RL1tCVUEQ8h/5M8T8IHYQx4wwGFpgBwyJbzbEvPbkr
I6w1oC4sW2iFro9t772FJGEBoApvtMM8qg5ajC63KIUdsjA0thSAdZwV4/ag3ocs
/HYx71ch4PLLlvr4mmbMHmJ8no0Cl1FMNokWx08ojIUa+Qp59xXW+4AX6rnm/dCR
4FvpC1UFyhSqSOwudF1MVkPrJvCnSm97EllhaWagJoU20Q46Pnsopr0H+YE50sDQ
MZADadS6Rg1y0Uv20HysAk78AsGbcnWzdijW8Fw6KUT60QiYr7my66i5JSjsW8rw
EhVIeAjJ8jyDIRyaoAKsOTW60wjkTc02eIh6u9jLL1m7Ttqk7AGluzlJJKTW9qbq
XdEch4bPCfrehCyslcFGrkaudhQbY1YUF3BTiKKyEBJeHacjYiKu4XBhnFFW/v+i
R01XKVTEfqnm6iNIXK2kJ5aIGYQjjUeBokgADcMe++NmOxSjjFk+1yJepUuAloPj
MKEXfdCmN5BSLhZzj+kosgmbIcvUpITmimJ7zDI4FnZNR6dMTn69/nPDj3QrKl4w
x1ZBeNO8feIdYcE8t0YqEz9IufsoOdFmUVCQmk0TcNKLoKBh4lDUhMl+dHu4RtyJ
F7JuoHyW4SPRJti1hsSfv1gRrYWwLfaKFAmOcLsezwj3PPbSLA9PooGzJj/AqHQ9
QQ36ymtZr7yyBQ67L0KvXnv2vPYRWsViM6YHvJKNYHCMvnnw5LvcHwoUQsi16JEk
+V9TUsL5cL2slRgUl0yb8zaXwP/4iO7VWgsXynQFbdnSLcnmnRfcHUx2nN4fpLqT
2HftCsgkQyqiOI5LQfwkK+seB3Fs1gaU4JRmfP8b5WrnYV30GnAVuvb6AgWasvti
OPjiBk1Vw+ti8LR0nILEa1fvdLWD164El/aoV13jG5X9lCm/9h6Jp8DoLB/6oWC4
0KDMgU/67IxMDHCpkSfdEe3fAXl1Etwxnmn2+x3qDa3fHaYRywXNZwi0Y3YnpzTG
ENb6FKDsEYrmZZeyJ2/uD7EfbUFnJj9tzdaRflgNdkxYq7DrrvM8n8WejwXC68Ou
aAzAqWYnVU/jWJ17lx3TP6NKLwTJz98gygI8uYJ7HOVre9YuJnskzndIJ0ZqK7BD
kIJ/u8vZwdBMMaeaVr6+sVOG8dDY7exTsg91WyKfDd58Bac07AQhsa2yRuAatJCV
WhioON5MvjEBfvXOuDFrwMgZwm6ZNyOBigwUS/hh7pr+UNoS9sVGdprHAhugaUN3
z0ty3k92ZlA0FApKgvuIdngdwdIDCFK81TiTDF9jLKnvtBzDvEDEHqgGZP+wSLW9
4dFrA4NY76J1ow0rxrkSBXnpDAJnRhUail/e5SC7NE0WxyDM0yOoXQ4AlmdhAPBJ
CYAUVNFoEbNfEQ4/DMMGl6SH9g/xDmvNIOAnFIB5dV6tXNWaJXMeU36rIWRkpOAe
N3AMukdwfURKoJWDwvomrWlZEipLOecF9/yVlFx+KTFT8vE5ZellHqwZ0tFKvKLw
y48Zb69oXS09ZN9BEq6zeATIcm6TYMFbvC2IzCU9Y2q2eJM1cap947YhhgO85ARH
rw/+ma0ZKHayHoMl3Ut+j1ZW8c6g/aqM9KjogVitvxU0nEkI+TxSALCVFIvxUAY3
hQWB1ZkKP/ofHWMW/Bnoi9wHjIPwyJX7Y34/p+VOBU4FEgILZ1BFU8Wbs3GTqbJ2
gvrBI+K5aYXIm41ufommxwhKbMzR0S/gIPjz5MIfhHr3Ao4tWttBroyBhlJYP+xQ
rCh/SnXJjpKpSOsNxXxUg0kDtUCM9n6iN7ciIB7KEzJJPiYIXIK2tdQJTTmWvcjV
um9v2SA8LDZJQd70SP0OhnT3kjSMxbx0pNWxlRkGINFWYqw76dk0eD8G+3qHWsDg
MNe0teFuqoJkPQkS38YJDcCxqcMHBWUfP5zJwplsMd8sHZ5iRzMUAE5ygmU83eaK
qY4p4LkyEa+CZKsnVRbZRhomE8hXYRgu0Aj2e443BxjV61DaMhowkT9Mvxp5Khgw
hVX0QBJV9CCKe+nGLSmxGU3lxFQ4zunghIKDlp6V8oW50JYumEDV/UpVk15wRyjA
DWTc+03WGz0FArFkhIIqFDPbkwrVrxfJwTFw1DUsDt12joYEhjTmvSbCM2CGxwLo
12SaORPFzrqJQ7B/eUfT0BAonvoRSIOs5KTjX/O6nni1pXbCn1W/k7EFNo6EEFlg
xmn73IrmA7wJA+D+3y8LOlK0xF7cJ1v16auG4wbYdxVZMCfMuuOhx4zSTf172VZy
aU2EJ8GjboPy6JLBcX4dZR4hDLDz0OUa3W64ISAyRLtRVspG3BjsZwoefqCiGKxA
V1anN0B66aBuAIVzEH6tbtZy4kxfbd0LaDtnvFMEArIZ7TPUQvur8bJwCRDVLaGx
4E1NIUs6RhnGkbrF4dYuvlpX5me1y95OHl9EBpTh/N/3akH2FtoIJhyY+cwgCT2U
lUC4ePI0ANf72lvFMkbTv+ahcA2g9V/Fzhtl7DJN2AIb9odemMzG4iGxyOWL3y+Z
vqTXauvEyeu+J5hMi9xpmx4/L9PMjUtv9KgNZh9z0gcFw+5SQti+eKFyUBQ8HxXD
QyzGfDsOoQLepZl2FUeD27Jwkn7+axJ/SlAqj6mpp25p0yT8EMHrttLblScAe2HX
zaje922CQAYEuyg5jberU4fGTTqe3PKnV5i9iEkVRK10R33bNzk0bLPuQZFpgxMT
5ZcNDexT3OU8yOXxvZyv5KRQP5I8UMMzUVR3iF5C+2snQxCSWnuurE19lHL4Pyft
zvu7cWaP2PKfJ/Wif+ufJ5Lms+IuoOp5uyyDAyVmHTgRAQtoWqnFZtP4Blh5j9yk
s4T3DTI7OSDYdQen8LgXHVXBGqmCWofz8Qag8B/kXDs8IBSIgf9KSl9f4AzZfU6X
pQy33JwkJqaiFt+2CgDEVr1sZDcalB0ZDFvu2vbjxa/xglKC0D6mzhG0WlghBo3J
FMsbx7yC/cxUtYBv3j07pkW6d0m4jmqqaoGOfE7vNeEjG4RQ5762GWwWyctwD4BY
FKo1QuCtdfFgH52nLyuwCKUUn+KlBWjfaEVPLwllEUKBcE8L/xwXIrLlPs/DtlGp
btZZjZ8E6bNnmE5yo5CJsU09q8M8rezaXqTihojk8lniCukczj+rCnQ+KJMYzRsi
NHUcvwMtA1uJP+T/kodp2kmrjH7WgJYBcIbkC9sZY8kV4p8cdF6sFOq0gGKymWxT
yVRl++6LPjeL8SucXELqTItqjcyXosit4N71r2povQCrQyMY8ffELAT6tIRCRIYU
Sl4Zp8kyiHHBWLUgWO/pf8xI0YmjoRBJmLWv5FO/oChngU4zsuGenl4PR0I7I0Rb
XFGAizQb+8lbD/UfLX4kLEJfpmblg3e085gkE3Iet6O3p6fW++3XPjinwKYXDxmy
J42vFox3iCWwPCuIId2Ge8jHt4unE1+ZGLQIpYr1IzezR3w+/jYV//Nan2uxtEkC
ai2Jn7WbjkqD5RlsKSDFSnNXyUihX3QUkiL6qZDLd6R+97oI3J3TjvpMQe+57BoF
DuNBYZnsq9RZpQIgCX7oCgemyKeFnE9MkM1Ok1MB4KyhJY0Bw1d3KSLnmMZOf2ko
azOkq3Wh1aU3DrSwoogy2y+To4SDT5Xghzh/B+ESuH0rzJlbQGSDaIHGjZebJRqA
/KtOKIfz0+K+lsekORC/4WahpU0UVn562YtQ3xB1SvUiRAjrC7z0flbtwbch9Orx
EjBgKpOlPCOkw+taYQGkdgtg89mtzlRIS4dfmGuZd9UkaOIfjpxiK9LcXbDO6Rqg
NLxZ+7H1tyClQWM2rqJXLJJ/FWI5TPhRMdDp0p8NhH1W2QW2RXyMwdfPwGkyEIGh
OFKjJ6hmpxt4g27EGZ0JhlARoeqfB8dYn0KK0eaPBvoXkcrYijgoycgt+EPUVPVv
QymR1HF4UWWLe3pzbtCxgFGZyK0bqwKoOzBK2YTX5K4Lc28YAKoXrDxRpR6gLo2e
G9II5dQLQ7OfNdqx4kc/oeAq4/6/9AG8VUCWbimkKJYHee5Xz1NzW8T+uG6F/UK2
Ne8jecfUJdvo5xcjf0J7eUcUUh4PtjtqTjQ6Dc/0ANYXr1QyxKeS8yfCuNgTx6DR
HjxCdUYfM67KdBsr8xsbw5iepyVdhRiY7qJiLKvDgywnDIL4ANMn2owqKcmOXsI4
j7OR7qXWmiBhHhNlaEtMgBdnZv5/svAtrSfjyJ2pDBKc+DyrUs5jQkrD01T+Xptk
8WfVBMya1ErYqTpYstVDY080HkNuVSlFRxtZ0ZHzrXTDpiQ6mTtRDSP3IJSo7+x4
2fVSwCXBUn8DblW+cOgFJuXSWbh4S0DDoAAWvPESTX4y2mTi7GAwlrUsznJvVbaP
AXECMPXdJTZEJJwshsWUJlswZZXijps81rtDHCU5540K+MpX1blqe2HP3D6HBHbP
pfmC3cBur0P02mVhHcLjLbQQSPQdGbXvVheZl1p5C22JMRqOLnrRZTcKOf/fCi7Y
dF2c8spmNiQW3lJovhjmfAqvAeqzMInD/yWhL94Ivm0qGVx8GQ6FpDovORXKN34n
YKsOUFFJ88q07qlPm20XvK0xlXLh19S6Mk9L/2NdOlN/ZpLAcHOvdbO8mQGQbhhd
fdhrjvGGxRIhNgSfxO7U4qdLSp9C4X3S2VcRnryZLM1s+EO4XuI2ENo6JX3U8rCx
UQcy5r6zz9FNVyq+fQCbaNksa/154TG5KfEfUwSKApwHhtk6ye7GMet9/3ZTay7+
MFMfHhAwfxPZFoz8XFjiIJkuu0Kc0Vg/A5QttnDQK/r6EL3h33SPCzdBoGX1BAEP
bbTUUyY/PqQ0epqpjgnKrHe9BAgwb6ojmWwicNXe+lIKzB0V3sM15tdmNtMucmu3
cZs8ki0KnIL0tMQsow/W9NrIuTNuDd4glZONGF8XvFhxPdi++wEqreGlISYTz+kn
j3pWfpNTa7fZHKJq9htU+xnmoVckmm9AGgsby1J6yoL4AqA/4+JAyWjO6y/8aVst
b4mCd5iISxbjW6wnGEpcJ7wDTavxblV5gHVfCZu7VedxdIwYsegk0P6b/UK6Xj7e
fLZVMPNTcRSWzTP9wHFMssv4O3SlFLewR0/Er+tKM8KUbgmlPyvV8xNBQkK2Hfwc
X/KInOSwVIqQpvYvXbYhH4J4SpNPBPOorR5QykNtvgMZIxre8W5mVq17LIA3oGvb
MShpY5geIuNCB0qnRAM8j+aqIS87P55ciUzVm/MM2rU8uC1axmlovtfLjRVThQdH
ChMKhblOJDFD/sV9R+J+WF1OiskMREde9hVRbil4wdjjJD7u5gvaQhB5FaTGDCRV
MWYNte9eiWnlIX0jxuKAbPWKbUv9jt0tuJJMdk5fSDHuYps3xzQn5E+ArhBFdtRU
1tySo9pxAudZVMd5XgLl2C/dGwuCxO4U4xhMRyRidJruK9znWtLXL90p6ESpqwGg
A72Up4UuGIYM7nkEGAZt8kjSKzisDHArgmWDZNNvadgBy6RQyY4gcjTrGjPgwRHD
Dz3AfqTYmIwvlqWGa1NYJN8CD7sraddeEJAMapmx9wpqLiWhJkMDwyE6kD0AjigS
HktY0G9WvtMnSGaCi0/rpwx9X7Ecr6doQW0a2UhNWxGa+zP6jRQskTsKiWHPMUz8
/P2uLiv11qlnS9c2ZBKXrwd/f4oYbN3sENyNuI+8xBbFnJBcAKCM62uTXbWB8lr/
/q8NDo5xS3p3x7LjL8qCNaPreKLZoEBcKSDq1VMzpzW1RpdtV6PHozrnK9buUjJQ
QCIKjHHcy3wKbNJrp1AZZ7An6muIZIqJjcoZOvrWwt4QYka6q795PHxUsuCdXJi0
PL2hWXB1IgujJmS//QI+L3WwAjH2RDRavigTZKWYhU7K6OzLwwBnVVu2Z737o/z9
hQjhoog8r6R1lCWzKgtC44dMLDiExYdVKzASmSbRa82DnV54qW6acqba6532mN43
vpOSCRmgEKNZPhDNQMFFpsh9esRinakWEiDmoo8DxMRtVYom6ECHBiIA2oafNVyy
7D4YUtRiM2eEm6uEX4s7LW6oEDPxW9O5Enq6w897HavydjLZUc6wOT+algTlvxWt
2MQIshpZhgSa6XEHyehsolzfe4s8Ku0hQjtRtDS6evJWyTytNmrDBtnMjzKO/9t4
HGf4IZweDCLhlIMUXkou1K0Qhr/ddawjOWHIYNviR0/nzqT2My7z/1w4pduSTqX1
zFxV6MwStIiTTnBOMxJdhQ8mXbRaS3NINKAemjgd9UGtggN9Ra/ao4tOnXqFna/i
EqpHSIWB02fPkdyHXSnRnVtBsH/jBklqzwHhbZwhxpW5x/sH4os0DdhmR4pQwzzF
NrBsc9fxX0WdkuOp9VveNSFnMfde4/hR9lyMIbftC76tvOuCKgjyMiITN3JshAzF
7wxZiMtgYVVknF3eGy6FHRjYOkVLPu+ENukwta67elmVI69tCtv/RltGdpp5Feyq
l1g8pA/tAEKj57tcrJapYLAbNYdrwtGOH3tst623Ylm4jrHLFTFDIOzyp+VTnE9Y
nmgdJYKanvzV0Y3XfecH/9Poa1rWbzWq88w+rUp6BvSd+9ml5TxHDsrc1sEAgNoI
f44658lryVqVBuBm1r0ekk9ptrvfZMqHfaXrj9psRRR4AhRiKuHlAghEL15pNiPs
uXxOdSt3omOYiUd3FuMhRPD3YuVsRMNVg/VQRcE5jMri+4k8BD9BjvVzlKXjwvPG
XAcucO6QirmS8aCqetvZom33SwPCNRGjqUoR1z1ZydWATUDzcg+DZ/MnnMrK8ATD
F6OLuJmLGj4BNJ6tUe7qVZIf6pulPNOaI9g+NpmdcskpENjp/1fGTCfsuCV34fjE
VSQlhxA7uGi0K6ADXkKd0ypY8ceT9E6IeA5C2A8oGLw4UFxuv76uUsyFZ7m77Yty
i5rSAxCSff85+WDaRJ8yE5k7erbHIcCTglhzWdEEH+Y0jPCvOAfzhoSXGPFFw0IC
zmLMJohMUsrv1yYzCdfuJeTe24bBZLl9z899eif4PHslcHyAgIi8jbxnhT2m3Gpd
7scbMZQQlOBUkrCVFBAwM06Ju9V5lsaDFtOrnjGWX5qIC8io4YT18J3kTck+5r2a
LXX5HJBDQxBbr46nTtQ84TXFrwSYR379quMKaHiDXsRz3urpGsyf/p3LlJpBtR1K
fp4cmhyVN0eHcvgywgFmXHRSEh4BACjQf8XF+51c7C8upeuTEKIDP7AL0lRUacPe
TbDywJN748KV/YpINRkgEoT7M5JHyR6Mmk7Wti8xtmU7MapjyRWX2yveNhLnpqUl
yNqKdqPyGS2xQj3/49Rz4h9+rscdUCSr+4cUklRVxaavdFMzaAc6tGVwbx5bDLXh
to+4BzfswPuUwjh+cALjwt53zuV7vIvwc/0lY5sR7VXIk20jrZjtrPgqR5BkelTb
TWLNh/H94aqdUmlssFCFYkLIEz7tCTP6qw+VIzqxV6wskdx8gDVKxrQJ/51JQfo3
2Gh+MU1mviryJjChPnGpsou2ZdhDR729mZIYeMDHdb6zov2yvjZmNkyx+O2uRiZj
h5EKkfBrVftoR0ELc3tRspushZQHMGuLWpfPph02kQFfsDb3OAcLpuWdLVwBq26W
J/2vuIf6H3gfD9Kj5uJcbuyNuvdDYL1buEJn8Fu7QZEx5tWF1WdyqnJZcGZoqeLD
oHIvk0kKpRXD6jbJMzt2D3YvXWtc5bGbhWXc1FUivZEZE0w8pQuXC73D2AfkITiN
ZsRaW7kAlP6rcmxMVYAKEodLAq1A6Dh1jvJbGbNGQ73Q0P2Uf9essyBTs9mxn/9R
zL6PtAwiN5K8B4bYIlnvLAoJbpH0SglJpk/8GyyYNg2700v71mzmtjLVgcrWBd35
pA/TaKPZ5F1zoSfP0Il7RLX1SWMu4errLHPSwtgZDVuxKaVs8WvfkvWyP6UNdML8
h9qCbMGlYLWtSNh72RQLc2g9eEZX/wNXrZmkFU2LYzKzm+/gsKQau60E+PD4Ximf
qpg/nnTLuCGIcLpb4Hk7eiLNq3IbqwtsbWTDegqJssvhrdXaPgl5QM35Q1caZoPh
z7sHMblUOLSrqnfktSO1PBBzfpT+INNIh9i1bPdxSs9Os2ZA+1lk4zRenq3QXphv
YsX67PEBaNNA2hGY+E5UDzH+4c/J5wP/Nvxzv8ArPhdULX9sRW2RivImNdhFswfk
y+yVhUK9pI/TnszPUPZnRIfXpnd0LmHYq7ApmUDHsnZJYverCBuTr8wBkZk0I6+e
GHIRDgpDukzEBQFTd/R2diAyDnHUbf5L412pJM5mxkVfsEJDGGgyEqGKn8LsxRaz
wCMbIdoasHFlXc+2tpRxIMKzlUIPHkxkt1cf62pRYbHa/ehgNv1y1U5klSumsw1x
0UgaGLbDOszENmTPKafqRyyHuQhqk39o8iW6ovZj4EI0k1zmf3CeArWAc8hsUt1+
kqyTGnz5x9b/Z7Hb6JnI9guWEqUwWua6V9PNee+GyNmBwaoWT7ydiBzo7em7FqXv
r0Ul11P1+nemMErF7UUazmAcwFKxrv5YEwy1kndPdC4rRmNqF0N3bAzQ/vY5Xy61
GMiuqkS5G3udMGBissXUghbiWWro/ADfr0uOJ1RNL448te6vgR6P0eqJJfC7h0lW
MM+XaYGtUojaMt6z/OTnFn5thutot+VdzMcNdHzvJOcB5rO7ljehosrZ3q91S36i
l4hA1EJ5gzUgmJwTlErzC7WAqurjG5SEMQWC03TwyCRfGuiYZLOldPQP4+sbCf3b
vEG8KwF73bbV9CTzH+JWY3lHHQBxyLwrtZ4GavYwgzl5V2lCDZSK/qx4clcYgblL
1s96mFGS+Ov2OI9325pVK386aVMdjU06oudnAZC2N87luIGOSsAKnakTP3k3b7E4
87XqZvfwt66Dj80f2cG34pTPYIa5HyL+blPyfkmC7m/Bw+jzwUiJRenVDyOzOknt
7nRNgjhFKESR4vq4dQrYBMs/iRzE1kzpvgPHuIeATDlSv6CW7GpwwqmJYpGhtlMe
Pw2yrJWdhsgg+LOOK+W6W/nBf1Vh8ZBlzpcfLMxmh09iMx3AMFsNpBjgDNX28FUf
Jh6ZRp5ZI2jzFeMZ7LP3Ya2Xx4wQFA/kLRDVs6CG3J9YBsemKPDY+mXJke31JBtc
fMonWry1dXsC6dp3NPHtJaL6hEf96c3nz3oEXnKNooEIAYR5huBx6AyEG6egpbWl
Pg4psE6h0ATZgaaoErytj/5/pbDwDOAUXJToEQvL9jwxq+fT6CKrpBV/tXAqxvnK
FDqLypI2bsgpXxk2drUy7jeVXYK513Pir/Hq5GGTP5SrkgOzodVUVIOHDy1VgQE4
f6VtxyZyWoCp0/JjoOpoeLw4UdwNerMC9LQ0Nvzjl4f1anBnB/nnQSgaT0nihfm0
uHLMipDMThvRAwbj7MfF1pgoULq4VLsKr7SBxCJfHBzFprDHNHvyitVBOKuCntbc
E7y1sjVkD12y86MtX5HITxwDbk3f2tH5vc6YrlmxHJqN2NE7R9qWLA5CB2mdfJ0g
9kp6O2LwIaVSrFzMU9Q25zwyh40roRRj/x/Yxy5JZSw5Yt9gmS9j5UKx+yKIoRyM
fo/qSF+JhoS9ujC/A/H3pi9myPjIyxlOl7+geRjwK0BFOaNfuB4vAI9GbQUSULbt
ZxgidJAo245VLcRML2Wl6swZ/Z5f+t1Z89A8WVR4V0lb32jdL6nuEQscJzHsGdi3
2Y8DWZOVnl3TK4SL71zNBYQBrUC270S5BjLM1+Zvj0v75j1P/8EQSicwmy6xi20L
Oox78lAI8G37zxb4f4zmeP5HUaHLEIvJD5UCj+RqH50jaC4KuTHaAfmISdYRmmW9
7oQktrenqSAq8t/5c8Co7i2VLX9q2owAhIF9F/kg+thM2jVx39kDv5/QlvVRmDWW
G7Y/SBQD+Fm7/9bGylDbA5BOHWHpXw2Xkr1kQ90smni69PfzTooI+zrZRAz2ekMH
mWKJGsZwXlBB3AeliCyfowQ+e1SpLIIZJSXwab9JlDlq1s26D82snWuf7joHy334
a9Pa5ZLimKtUr1Ky+OeiaXSRIN0dArmJOeuugmwJihI8mnjoBfuarw2QmdiKutCJ
ZPjxfDScGIOZnylzsphriyRdaET75MvtgZIl7mgy8FmZy4rTVS4CPpcKcCyU5fk+
ZkaA5Sw6PEGOivRHXFoIxjr9AoDWJoyCc/75+bjI0DMOFvkpAbWc4Pc7jsJFnViG
7X8wVQSqY1H5EdVjwPT6CbaaOB3U6Y31jTfbueZv16+2crcLMV5rk/9YC+cyjYdR
Z373l6p5iDCO1G8BgOWP4OLQH2TGzXy5IdsSIB2hrkyp3p2JI6cGW+q2priwfdWR
inUrLKWRN+KoRrbW5ZmmZRphG+Pn4znreBShxrL9YRybhWQuXjeE06JtzwcU9Dxd
vaSX9SAupbp3F1izARBccauEVOtkOjdgzC9zj11UotMiburVaQtzO5YdgytWEf0k
u/1aevjbAL6o/pvHnxE4yNn387IjS/8xDvh80f6kGH6qVJhnaUZ/lte+EdOkd4/X
eh07dz6tWcFWkAeHyINYuhuu3hYAW8xJ+XsmrrMmwDIgDFvhT3aaNHDru2ygZYKR
mAKnchz8hsyilU1YSdWS1oQrEEzfC4jcz/2b0L4ggPumLyRK4nCu9a3hsikZYYg1
mf1SoFDY0SZG9wkAlCbNB2fKWrWSBAh71WUIL2cCeEAh2ZDPG7TooGyN19R7L7CW
d7qO7nSbKLndWj+4Pi9fj73LJi0zZEulsZxY47YpJuxzXBlIV6JvthIVqR8y4JN7
dRnHLKUzDglTzrhn2WmuVW9/H/l6Vvqgx4uBnNwW3TYPaSRvHIczeGq9OXIQAji+
Amy9sXmngmvEQ+ZzgrqRW0h5hGvKqsADK9XwmPS9IX7xOtNS273CIS+3wF0E8IFu
NrMcwgM+2tCRWTIJbgOe6pviZWgtEjTVBcVlHpLKrz4xQI1ytwch1zIQqCExKY61
QFgotqlHP4r7eUwq+SsotrstZO5VL5wyNxRU/Ut1lyArIZbS5kI/bNdjwchLRiyn
Z1oGJmaJs1kHCfu4vi3zY8lLehxvB5NSXlk2uaD9Ih02JB9w9if2PfHNVioTfUGw
ZNSmTcS0GjfhV1V13YQ3EwUWOofvvkyAsbohk3DTDgjiY3AJ5AApn/cRaXlApzzp
SHtYbczmp2EY/R4cWOb8AwyWQmew2UPXERXu+bMeiotySm75FqGNX2QsXD/HOPW6
pS3L3AxbI9VAgVxR+GUN1cO4XblituO6Pzi974pxEhk9CMtCylFeex3WEP2TZhTz
Op6IggiValYICP8Cffw7X6o76Psi+BaG75IZq0BK4rEsFQ72oHZk6ml/VzkKhfnY
giuX324bi4C21G3aSUbRJ/8sXAMOR7qjutYMU46PSUakp8NA/Pyut/o9TV90ytqj
NP+0KFj1PU89puHKaxCLPNFd3HOoCEmXopeJz5QcLN3OOAVYHaB5kp3RC5x4hRr8
VI6qIAERwmA5MpkCCZWHBdLWtLOqd2SD+XFq5Wqzin4medv4r/MjgpeXqU4V53B4
cwJNPvM2pzk/A5mxHeBBtFg1icLKKqsondLhddfPbrf6PZkwA+DLUVRNoFSveM38
M5jtOoKu9saPHkQYAlQ5WU9rT7FcSR7nqCPN0LFQoTi/Bn9TY/4Iew1JGfO4jTxx
6KSUWgtJrFqApuqWzsj+VQzUYnUFd1Mea2H4DX+7vNAdFoAswOdZ47kxRicrHmjA
W04XtW8eHhUgcaq+kLGZajmElhGJkKv79hSyijHrd/VuxQ1XQEMdbjvW42j0EaNV
6xIvTeRNoJLUKYsAtxTr0yzZAJDsM3Eu2ShU63RtHitFpMlVFEq+OXz4DOPD51SK
vjUpeEDf8asj4XaRMlGdy9EpWDYwocYRjrcoYl9nZYWu1/lbei1HhtZuboWV0jZ+
mwxI3CdAWMNishsDgaps3cbVFpcYermpoX9gsbyvYk9/SaIjm+bIlcD95674dx7s
1WweSzYxZBJlSsecqSYNtdNskTqC0OOYH4aFk65Ce6U9ApA3KpcX7IrEglhlZZdY
hP9MTm7zpIrFfj4Fsrj+hp33KFMwlDsGUA3l6vtm1NBpz5t89h4ummtVw6XJIzaW
z1fJf+O6KiP1Elruq9uZkLCQeE7eGM8/cz/HME1t5YbLAHOKF9hwJ0DZBYd4+7WB
B0DmnHjeBgFFm8xelrSMwVmElSfg+uHKc2lQ7XiHmiX/x8LaxSgOxfS94spCorYz
hvgaUa6UFkwXUMP7Nu1jPDzMG4apb1i0FGimuOtivd1xQdR8k3p/NOzIGzUX3Q5N
R2wNrWlpkfdCHDFfgA492m7rSz4ipgy9/gi0hmUyuQUgqsAJjXMUyqBtDXmuQIue
AVSHKVTvB85wtg+MliB3pKwDDAArePWtfLOdruQN8ml+bmLxmi+xBPjZduLwe4gc
4WRSjIWIF7+B3v+//aXahxKN2Mtr20OZr8TPOowGtNOSDQaVgWxHLDV4Yw7PZElv
u3XhWW9ZLon5A4JPgiCR3IahGitAuTr/MJCcC8pZzwE9/gfrM1jrerz+9X9eVf86
MKRsi3IOQEjHVVhlKcHH7CkkQ90Oibq55F3YcS0SUZ4ZtZvZ3UixyRyGR+uPAyWs
MebFm8gAaQvDZrBreMuT06RiOMVr9laXmHc0xEA4CMia1hSqHoMSHaBZP4govaU8
yCksq6qItjJ+uLAYXznarByeigCCzt/uaMO/NH8UU5dfe3sMruSML0772BUYqirH
7WjCk6Zz3QjENzxbZ/jMVTaXR4mf3JLE8L9H35kHO/UT9KM7Tu4PbJDPTx51nCQt
BGDcnQ6qKO6V1YFB0jBAu2wE0a3bjSk++yLuSFYlnmjgsYTg4uBWXKETrHZEI1Xn
tTMACa8mOFN9cpbPZKx4qdyxv4hhDuTYtxsagDnrrSoBm0Q/R1JMuDUB5y9RG0+L
R7YijqClqUSzMW7fzc773dZna6H0AORxEx5cLoA6UpipWc1qGiwE4UXVaQTSmLUZ
KhJFg0ExmGtXxIb2h1pyOUOgtpwfJe01FxweSicJhO4Q85/G4jikePR3jTqVAuJx
xbciRZ3ajpDAEgvOp2GNqn7NQUDQu+ibsatMtMaj5zYNRVs2GYtyh0DjjpVWF0Da
RZKg8q1dCfJkmYGhpFptUbI0gElliJyp6OglLv+B925gtIpswlqmDzOAdxC81SVp
xBRZW2ZtRW9X2X3kV8wX8tlysedTlo9wK0AsvkHrB4sn8mdhK04VaJdajYBGpZpF
UFBnc+YsWGSi3tkfR4cYfSZ9Q/fjXnlQJzhifi7STA1O6OwnDCyF0mZaCm/oi7pP
iUpT03xLehXJ+zIUIJlTG7xPXOEY2RcPJSmT0T1bEC32Skz9vx85u86/w6njvoA/
D88Z1xXhhW7/F9Ut9zZdVvYyL1oBXTSndaBQ9CLQ+PSghAbl9o2g7qOHjPS1t82/
7mDFeJFmZFfuc4tYeeP2FymjdsjGzZMI95Rf8kojpkIQbPnUCm4bNj6S9rkwTl36
1wA1WH1+CtMvrMy1DRwK2E6xRffCurRSBfBl7mGkEh66DoHT8mn0Mv5VGbA+C3ml
mJxnY4AHfu6XGc/bUEC+4DYy7R+nxgEVG8uxf1ANoy2wsOaab9EV5gUq4rQutoCK
GTR3D2p3qCnNc0F1wnPHiFzRYysmLDGcn696CBbxhtiSwTBVnEzx12iX8b1H8TO2
OIDlIPjCKQYGvuxNQQKCeQXkZp8jVKSADiuu/4g3J3v24u+1/Dm4K51Vg4/RnEjV
gscDyeY1S5iYF3YmNRC3AEbVIFZaakvPZIAyoi4hFdNPMW+Q1tBpzNAS/JJUgnBk
wqBub/JWlsKSR13v+AHvcOumjhwZfwwva5i+QbcXwunkp7CoBUl/HiQpL6XV0xCX
p2rJJUzlL1OCeH1a7+28u9tj9xUpGHvf4NViB9s98IrWoKhrKdeUVFjoP6quQzV3
vJja4PaJ60uBar3SkuoEtKM7Mtrs7JEAdWrOJ9vV6oXuBA4LNY9FOvKTtGP9Ssvy
7lsUCQx3AKKlfMWcb3/YgJZAK08I4m9cdD8lq8MWCLCocXVpRVP8UIiy+Nm5M5PO
t/3L6YCGLoJaXikFRkltUqvzy3oD30dj75x+g68LGafsZYJdA+c6P9LAnw0uzuLg
oRIMWu8rVDWK5eL0Ptynk7zUP+PJLO1ozvBRzYwjDKO83lx1GNFKvkS8aMGsTzq/
D5WwPCGdVXLphtSP7zdJehe2mkzIBYqaM6tY/E+TydOFp7P1Q2TqYYCcsKMTjK9I
gTpX+N9aokiInFYlp6cxIgyrvkgWnyHZ0hGVweyL6G7jCvmDQn/tldb2X3w2ioKU
AP8jyWgN8O5COXm3sbJpoBDYStO+YyD7F2xGtgnoOWN3khn6vW2lDMO0DKvefZF3
etTbqhArPNx7OhQg+oQiriSgsiYDVDLjxLq4vs/tRAhCOx5zvDt61ri6RgXEwCzO
6m5OKBu4JDxwskirG5LsNFbBfRLdHyhNQqo1+8ZyoG0KYwjDHkfHsRvTecAelhcq
njp55p+Fd1LqrG87diEN9AcFFXwLxewGedp3TSb3uAbOT5vJ24QVaF+HOq1i+jUU
d0tsmXV8i9nVrFmMU7BjIgDCsLZD0uhE3EKtdPdNHzpBsIXH4KOa9ho2RT0rIz5d
MItGIR36FHcLZ80Y0Oc2gMBx+juv+5om8xaiONH1KuiKYu8kzWUE3kyTMmorvOjk
XTkfbs3Fpv5Yg6IoK9z2cxMIPRFZ8thJfNUdccmzkh5P47DdrXLV3VPajZLTG0wD
+Ymtnhnmzv1pugUnlWKOu42pcWCHv+eZC/6ZLxM0/SsMCXS73YoZTIdSk6tfzIUm
+trWOBCAoG6aLJP2Q9vSmuHv3VN4RPfHg/C9ov2HsWILJ+SQa+ShLgaG1LJMy+O5
9yHueMLkbYj4D3zWGnBnjbgo8kxmwlqtFykJEJgEQtTkhvDbMocgub1h09PbK+jV
cEnkSHcRNIMnQzJ3mQoZxtpG+nUSJgBSGoQOhJKjNierbmzKj5fuuejMR82uy46s
MbB/V+5IAgLsvmDSdvpQVfIRZrUzGkTKaBcVBEP/eqQDU2oadCxv26yVJz+dcwV0
AhdAvWSL/TzwA9pMzcoH3YMFU9vHic+FHk5tfOZ3zCsO4csd9K6A75Z5NYRUIFqQ
xWC9Uzk+MM6vEf53MnC8N1FU+EDniPJkmrdUmOeHcv20pu1eIHJ2Vl5a93jKsBoS
uIIK5asNqVD1FSizq7d5ZJeJtdjga3ljSO5ZPHR02N3kba/rXWmCgu9J3z6sgqP+
08UnAiLJqbonUhZyhK0HAFs8hfmQ/V4OxO7ll+0wA8t5SnSKvwtCsFt0NBOsmaHS
7ShHWpxGuO67g1OkmzSN/S6nV3Mg0utZ90GA9/AboJO2j6YjqtmOqgT6q7ZWWGm0
kH33K72tmSmzULWU8ssevKVQQrgHsGM/Ti5xuCLgNN71Qx3qlQn/sA2ws/NiKs5V
ryamR/skVjYTnJOjuQa63qiXsz61DUd1iplFcIx/0w+/iuwCq5NSa41kq7Wbk8ii
oavmx4nSnau7NwQlufwO1pkLXAvfiPNcZDbOTI7noy2xHwDPBgcCzGyKtTq8Z5Ik
P55icsKh++W2SRDUWfKSTrKmKMa8QLFyA2g63QR9bNm79HZ4OXX5Mh1ltskXkqrO
xJg9VPlWmJOiHMypMytSgtpt40SrOkVL0XC8XHpuPG6s9TIUqZRCFbXj0hJR6Fbl
GUgeZQ2eaJJ9PgVQE8qlmBTVI1coS1oRI0YvdkAJ2Hx6dzt1TQN+berMM30+U1yk
5wOah/VAYGgolpw1ANi3C+g4mdjZ4tNpRoIzUd84ZZJdvn612KIhCYeunI3TZ+8s
wLgC1jo/sLVWGPlsok4wC1J8rqhr+hT+6MnSQs8Lklj/DDBOKYpsBt7WgfQBgtLd
TmMSKzdLWRKrSI23htfalFAklBLfZ1VHYa9S9LoZb5p0haB3kP/yzo0wGRAW9n+C
rb6A0l0d8IAW+fq0GhnAnJVJAVbjord8oXUK1V9dqFF8RSTvw4X++9XiihHqdZA7
vZiT0hJBH75LJ/I/wysCGRTgpxYuAaIU3jG9ij7b7B+K9ZphZ2s5fM/5OYkLc4Rl
UVlnZVykmwtaUfDPiWg3pyy0YsNWC3HPjEzGVpOqqMt8S9am9UL/7pnE1tBv/EfA
yEukTkjx2YG4Y7mlYUcQNICnxHNRqX9pTeFDJoEU4KeYdW77piJNQ8pY7LR+IqGM
c6c5pcOTxZ+qNyZrXAY7BACP3PY+SrQGtoIwlZKqVHT5nQdSCeqiIAqQ8iOc4Wyj
vkInPbFyfECNStVb8UWv8CbWpEjQ9sEuTBWD2+x3eWGzja2995waDQuqbqgINRdu
f0OGUKopT92jKqMrkoluqW0q5TkJhuamoHjqYyz8Pb32b/wY+CpfJgpSkXeXs8F3
Cd2+2ppXZaq/wn1hRa2x8U+Zrt4jQ0c2Slni/0n5KZuCe8u2aWe5Rs4A0EB+15Z5
NJ4GLzH3wZuwCVLWbBge5BSWOsri8YRVXjfjcSh0TZFA5k0GX6x1tz7vH2pq6Acr
dgo8xbOcbjGdz8Q3sbIMnOlNltNKH2IWcA7BhstNR3mXR3bsS610gPuj3dHgH91t
3gyUFtzf+gbfkPxOZbqZpjISU1CoPoyBQZf0mXroVjkFiqrbqcupBfHjfo1X3j6B
dON2boj7X3j8EjfPpztANdrwo6/DwPdcLvfqeEhZd94yfOLrK6Bt+eS7hgfhFFym
7jbC9/7CTNBskjmRqGTsiVxqtQB6pAS6WSuSnLvt0AVLZRTy0jbac7+sqeZt68A1
2r2KVFox4a+rTnKiXegmyDILDe72EudbZ7uX2eVIqR+pi34F0YIXkutRwBQqgvIh
0+MGTNmKOreZIb2d+LRRPdXhELg+AODINJbo7gQVAAoGKZNSN3mXMOzrUejfNYrk
tzzqZ4HXW30g7X8LSexqLYC+faJRCGwUnOVzAUFiuzwLkKONdwQGEfAsVyb/8DJF
GM7etDPVtZxH2/+U3w1pU9t1goqgWCh+VcuuvAVKDeAWCZqC9EGbKZ/J8vsWCwaH
0qHAMN19EKPSDoqqUhVFq0R8cONLpGl0DUlXg2jwgPmE3uZe7Wapospqn/v+QwcJ
1FUvyd3YMLdZDCsKnYFt0DRpObzNPBBrtmp/P79Q2ITiZ4b9cUnGug4VeDZH9ZF9
CleW081XfpplnuWDVJVJ25b91DdVwJ5dX0otRgcRVKA83+iCaCP4rF8U1TKMz9Et
I4MTgiAMFXalBorh5UGyEmEOk9UqXTZdv78X/XFtJF4OR34aIiVKUw8xuLRP7+lf
nzXS+YjR1z9YViWvC4eKJLIKgYpAyCrZV+A8rr3anGwDa2MqC2yUfv5dcGeIt6eC
rLmtQKONO0ApaMfIJOJ/SE85a94UOhTibwrd3+tKerqhMnyXvXxMQilq3IRk0TFU
8t3l3OCadz/5c4bvqkwasJ/o6yVb4BMpBLnYIMzcf11Y01ehfUvAeYOGCrjh4KU5
WllwfhKM0Vb+dqm2ZJBOpMG2kowNxPtQPrDYWCdOHKBUrq2XedQqlhvsHwiA2ebl
pPxwBZsfXewN0RHFGyIutT1bAfCzhwXzo63AUuSLGPcNnOZ1FuWPkFxQe5Fvs0Kr
+vqOgfjbWzy/U/uSCBrp5znogSXOQ9UGh0AnrdzsiEVIYa1j0zZRqVhcl612rqKj
PrJm8k2C43LKU6qMcyYV6uPMO5pL0qmEmH1hSb6nyLogClGClsdA2mDf77nvg0xx
dv2RJVKiPhozHWl62RO0Rsdh9dyU+gA6gVNvDD0OQ8x6IuUItrvnNP9PIgmt4Tu4
YW5SjsHzX5Jrt4eiDGd+1hX1dI1eHRnXMCbJDPytb3IKMOBCH2tR5+wIODeEl205
6et+Y3o9K9H4ZB/V5cGkYRrkz2zpr26gy8BnDwCYY1mh9BVaEZOQbGzoD75rjc3x
DaUYiib4sJT8AoqO1CrEvHr7c6d38ocRrfDvDUKkKgwN74jjrhZAwkFNcUedN8Zm
ZuPXC+JO+VpC11lRM9XP6SBhqFReCEdSIGu8RG+Lytm2tke0EToTMxKRSxtcdBR/
pJ5OvkDSeHRXM+AJtDouBLr65nU7md2vi8rKtlbHj6jCL787tt+0E9wd1Zn06lPW
iOlU7caFA+lL08gpZSDWOik5iAiodhajsYLLXjZMZx1K69uVfcbYuMXfexHlOrdM
UZrNY/19YPhnNRMp87rCMg65w7OyJ7l7RdBn46+KYvz+m0tFwQoANFL2wMuO91Jp
bGTfCpJewynTn4zGLb288a77YXRyMuoZmTUek2TSSRrgw65nONqGhICxWPequwf3
1QOFzAZ+SPxzCNmeuV0ZuO2Zf02au+Da6+SlJcxSExbqAlDTd2S3DTCKm3h978W9
5m+P3B+neHO6g07dp4a01ZJbsKQOBzctTUVHW2u6D6z+IMP84Ze5vE2VPWdBwGlG
/HUPYCtPhwJ08QDTMVXvsTB1TL9azll+58P70HHIWM+L0SLzjgzi7KURokM7uzwQ
aMeyiL1JcxK59dhPGGHxNXl7ZflPZ39r9JUHSLyGo42OpZoQmPr247s5rNiTmVrc
BhDTX0IDehisrNs2UjKSKXTu+2rVi0I6JPX6INJyisq4Y9V0H+DQZnZjYgbMa7sB
p8AZGPN1yfHA6KCQ+sN7iFoHWQYyjFwWwZtc0lJMqatsNWcCbKXRoK2SSgF4ZAUX
LzsAP8Oma/UO1+H3bzWsBYUBMsxmtiSCd5nyjfacfknRrOFpS/WqzfUqGGNv3dFY
/qukChtnCSRP46UVcSOwASikwR1QZmrAgwNLrBYA+u9pPiGMuMhku/e+1kcAa+M+
g0hjn743LDsk3Nu15DkrPUU9cf3/rhEPzTanVsOMqa6oW2O+bA/dsaXzAoz+EikQ
vKQRSnXExiHHtfo4m5lNvMoCAiqz5/hfIjEb2v9BSyYmjVcvWTgivtnkIWM5SvNA
WGJaiOt3xLj09mSHFYjciafqXVlBeGOEd/MEeCqDaNOGj7WLdQ3+Upp7cmf5+G4O
8rnrbT7jL9vL4G0qdWfqL7ll/81ff61Fba0OIT6a4+j/GLljVfP6Pim+Bkyu6zt+
EJ9B2S+O8W1NJDfjm5BnU1GsaDEpEM963KuS9Vro9dlKmxr1RL72PUWmW932v1IF
50p5pciJvAjuCqoOMoknGIh3GFiQeuMGCANXAlJmf2U5H9Pp5hLq1KTs5o1Drray
4MYM+aDAbeBdEJWUkJS2hwbgUbxoydIuwez+S+XSE/gJbWSYgRXetx/NgCbvQMxG
X2ejYi/utNRMnew2HN1iYsHLPjre5rhH1hyjwjyOho9Gk2g4+mGz8WSTBatm4aYs
5eJYo5f1sMaY/jQF6K8b09LsKawT8vlf+mxTARNpF3HDJnbokXJMREVGjc9jDOnH
vfkYa329rqD66Tuwox0d6Th+EAQk4aEtDWCv8bjoQBTchOfLkmO4oxPhKWoGhgLD
nO1q9qzKrJIYD8cj7M7hkuWMiN6c1fD8L59FEj3/wJiJIdko2Tr9u01y0OtMapau
N+yj2MHmQ+micUXieHbkQJ4pajNDP3cXKvHnpRPo3A3tBJWJH3mMBbi/Us/mL9Vk
yVGBEzSJQ/jSq86W69HFIVm0sCF3wdxI+3fJs4USGPDUOnHHWQN7KU3yN5A1TGk3
H7c0frcVSdSaTIIdyhL16SwHdsoXNu9pVAe6RViRbC3dUZFCZzANCNMJnZw1PA7i
QbhDTu/FV8Uld19m1e2eDaUgEyGe7Mtf6hiTqNk1et11YTz0ErEVS48wwqzgU/lX
7CkKLQfQcpkaHCajApkOeuDd31R1fskS59/CcIcj2JCriUwMUFvWOMbL2hLxENBQ
CROzpRN4lHQsaGA170SUaOJAqZCb+0JFA6/3B4BEakW7+Q+b7TSAV+Fc2moLLnHo
7KiwlaQvTzEqvQdirNlxKAOiNogKGCDZxX+wEd53fgKxOP0s1Yn3/zWuPIUUJ0RF
YbpJiWU0xjshY0GM+TqG28nafcNlASl/98LEuJf4xRuwCChpdVWursbXitkYeOqC
OL/m+UxMylL6KAjhvbl2nl5UipfKOrmOZGu9lNEEZgUwnTxNkTJKVmAILyKZ1AJG
K0JTbDBqiXIcmWaSiYRxIR0HliBO1kJ4ycDzecXebOVksefSteMc9aX2QBx1HZ+P
5t2jD9kKWvYw3K4w1sDQ+UAaTeNRhd/5FqB7H1f/gffPR1Mq6/6Wew9WYMKvx4jP
Hf4eKC1aq0YZiq1ArXEofdvPul8RcVZPMY24D0X8/kS4EDuMjNlljB6YB4XzaI5R
mCYUdQSsRO7hkFxR6Oc4x9A3DJfblhKhGR1PUUp7du5oksdkQBXjfRhC0/uj5T+x
zbfQXBr0FJZSJuum9LvtQGCByugyb5JZuc1COfClMdLbCRMjZUel+Ps+fJlI8M4r
70Z+ieRYxnf7Dk7gDMijoJ4QCYRx0B/yweMwlMfCm7gI35hO9i16uWotcKwKb5aZ
uG3GBZ8ZetE2dNMSbv3F1s7VtOYqNLH4pfUaYFBKwEMkcCv5d2qWNfEeMdxWYdu/
QnkU/aKpr/KOx4WiROfCTv2dHLsAy/6QusK/Lclxgn/7IJPAm/Nl8Q4Q/3rInBGP
CKWqqWF+vHbkrezvSWiXEDM2FDnC3YObOqP31UA1XxaUajLSVr2lksumHA7lO7Ez
xb0aKVUGQ8gZ6wYqgKPXTJ5KaAKIL1Z7Fm2e9FVHYp9YwBX6xdtOfua3/LrhiKup
SmU4byaKMRMSeLfy6auzDiHOpoDc/GQKieWXN5lb9R+NIJXNfGc6ZPra5CEKgNBY
LvsYp7+k61wXh7UUHSg/rmuqs+H29U4j++V3+IELAKbDs/Zpe7QIcR8rbHLUdgU6
WfF0AER0ylnnsHQiaN8qPR0nJxT8RgK08JAREyFtgWm7IIvmXOnzQiw94B/PTMaK
pv8nklL5gZLNW+8CFkJi8UtJ93ximAbyP9/1Vn+XOZYQmszwlxJWzghRLuZEMPf2
wKOQbKl2AKYtyGjGGoBJln7OMfAwZVGmd5kKnFvLy4LMFZgrX3P+VGpJi9PPD8W3
ecpqeUj+idNnOvGc/lroaelYBJwg9YBUQqtO5RBtcjCur3FhOHc1gJzDQ9XiUULE
zT+v6b2yUnaljQ0OGIDV3hQn4Sio9OIF2HmbZ8Z5nlPHjxN37pQKGhNztOXTGSWy
yOAvS/HtTWiR5WA+CpKHoA1jycDVrBIHVgJoN02MJbaInWdk6Oxx7PhV4aCYCs+R
xgKZtalMWZORx1DeND8hWYQpkCaFi7cXJ+Z1Vg6IeXS3hJ4/Xc4xNXNvic7oNQhj
wYIImHiU+SPyZh32pI7D9gHVDC5F9fTmWs49LHmV6nK8/nvE9Fm05SZ678QHhhDR
1xbf2ufyBtVLWlGqTSIzQMQqupq2beHYPYv2RA2aLPPbqa/RMGaV5jJw0QcHcgUB
l6j5OHfAegHDwi7MsNEJEAntOkxMYTrju50lG3LrWgb00902eqYGnSc5GFicGusQ
m4AMVkw1aiQ/RPZtFmshXPfM4wbw2gWwhf2iTmBMPVuT0tQw20zeS6wYIkhK9RHw
UD/iomkDQPJLn2GbBnFDrZsDj5z1JvfET0Yr8/TfmxNpKL1/flLbue8zmx1Pq2Bf
/nPWLaAjjGFzD/USiXLKKjeKVk6RwXhS6COVVWns+Q5xlMiL9rR2nFsd+IT6YdFR
ZnFjXjak9IuuVw0bA1MDz97Wcjawm9Y9a5UnDO5SoFeg2pMHyWiSMUxxE5h6cOMB
uYWDmadgSmxVURLDb1yTmkFkGFHuL0LqQ9Etl9XQqyeHbTIr0qHlo3OUpIsIY41K
zX3QmXHAEDYCdcnZzp2lmf7Wm1Gvn4qnixlIrewMwu6d0ywW2FBudm5/ocqGtGvn
DdeD4KdaTuoC9hEyEbMwFWgWn8DWfjaeu2IAM0z4k5uFT5iPLy4IAluexr911lk4
+VF4pcZFc37LdHO9/4voI0ZiNxFXoQoeMHYU5CqIVc6kYwP2geOgWgPd1eFMD890
xW/DeDxxAFbP8c+HiUVNygqfW9bsEeTp6cQUmmdQRikOufMEOXfznNyZRhfcz+k2
nX8xbdXriLp0JdeWgYnoJ4c26ufRgsr9R7ft5EeDRRJe8gOoaP9ySO8BzUGximxS
UwAaeBYD31bbWxudXG0XdbzKOw4BhQr2B+UMnTz/tGVM9+f/Gc6AEqBvwbjzM/1b
AxOlNUD1T750PpEGMN5T2RTKBqwxcOh4Pbrzatuy4xfeyvpYvi05+q5eyfQSrY2Z
fckDGxploWqvcnW2S6QtkSMh2CAXd1HYGPXMkngoLGFP8z/D4HvpHF8aDqLz4+ww
BVg/O1wGJ+zkHi916FNjc3cfV1iG7GoiwQeiGi/b7uChi/sYepiYuzg5Idj4w+JW
eCaUAZ2ED1T7y2K77Popd5Dz1FJTCtqavKouhaPzPNHEzf7+w3q4lbW4ZYcA02uY
V62M4dobEnFTyJe5YVwTcS4G7XRpbCpO3nFT8wxFULAW0x76H0g/2Mfb+0bWwgbJ
0l06a/k2kNcIhVboVv614+pTFMVFWtxLWDsrdkzJ8mt+1ChMJ5Dmkr2ca2VDp1IR
6iF7dYOjQ9wOHfxh/kVV7OIo5HGGiyoYSWbifC22X7AX6KAjhWN/BMaCbEjH5VD8
jDn/Gd3/qiNM7/2j6lnhXllCja4YZVDo4f9N2UWZoCi7eXivSPov3Nzo6j8BYrV9
y/cHziYnpbqbz8dpMznH0JJzDTN5KJDPJ78rXwOCgvjuQdbYNFf5r2tpkkHyG2mc
jXg8Eh1nRm0JzCwtc27c+vOoYsd4zHYv/jgN9Ict8qNR45UJ4yhKJa9u7RYnW1Ru
vW9lssTL0JL33rkUpnfZYntNoQWKnuHk2u4hckorXSrwekyE4oXmbG7Qq/djNVX5
IwVkE9odAcxk6gMVT/qg9SYi10G7fJHcm+sYqlMMDuJ9thcZ7tWHJ94YRGErZdzM
9bmgnmXXA/azdWVsVhKHagES7A9ao5MwV2Z3FFSEQjWT36h6JFaLPNWUKKHUE1U7
UoLZxuEuiK+kJluF3j3qNHjqNdsxA7+o8arwtZaKC/qNwe9TktuGdEgoTQHDP3kI
qLnburIaGEuV/99qeuszo2L8nq5mVgxtB5PhzVKt9zE+sj5crVqd1x71+Pp5E/9I
7otfmXQb5sLZj/UOZypPW8zXRvaj8O8Z5hluFpY9kTS62/hTpUP0PdXuTD6DkxTq
26S8tRb1btp4ZycQG+s8+Ft5veubDifqkEnRUjUukX9HdZSz5bvPgIML6NeQp6+3
suiYjRquYGjbl5llQiSWtMDaoOmAatpUhm8B3iwPqE36PDU0xoB8i0PJKhqjV0cw
zodoXvUuoPP9IvtIj6WTqOCziqXNz2E3Z4T5waMYVwe5uLDRo1BrQ7Uu1Q0fMpIj
Vdn8eaW7cGXQIQTzlcWYlqQIuXZVceRSrhmJs5YRbSzfc+FIo4kCMkLRgvjVaRjV
zdnv/0ILnUtd3pWTtwS3/JpueXa33VsmuBDqUoZ7ZiM1bIlM3TEI1O+jhG83TXjI
YLGllMV4hqKEdhO9yNYX2DzxAagGf2EwvJOMKlVylWuQUYoc7loFiyHzEpF+bVhR
daP7HXZsWO9pdtcIjwtgVXbHBrE5NZUzHIXzJ8S1DMO0nHMsm6aEWkPat1Ee2+QA
1MGsMA+L5nK1mxRShdbnUIPzUBxjNPSzDeffL+b8UXlqAdtxSxjspiCLP5e3MLWA
tpgjekQ291np70OVsh8JeolveZnQeB3iPN7BN7JXgNueTKEE0oR0fssDPqE1OCzJ
U6vwdt/vLeBean+zoqc9MFaRCU3A7itguuIpfe9Ul35JhgMDcTZuCEgBRu8Fkx2y
X+nXXaGWVPhxYJo41BQRawQxUXYCa5pLKiefhMJBN2p8ruiZTWUInLYsddy4kvqA
h4gt67UDWINlFunNHKrkn9PBvymuwLURF5G3swO0TT/lMJE2sh/qDfFVobQNJsI2
GVOXwNo9hT6YhVU1Y4E/XkuQh0unR96dAPDVzC2lTKbo5aixloO7w6pgKAE8ihTx
uPkv4KuwJFXUofbMGTSyiPDS+l116YtPtFtXI6qILKwvstFWVXHhqPjH5ktOuI1o
pBPXS8AL40aX30zQZKsz6TGkWiOh6m+ub4YMrwO3CnD1VI+MSPCUiN1VbJ5DNcS2
aE0nmWwH8N7rA8qgahDyl5eC4H62KzKLryQbWM9ThEzINnYqdo7h9AFsKFD1Glok
ZjlCN9vObF2kxhDarjQyLy3fY/ifnV70fcVywMbPq2Xv6qZRxqOR1BuQYTNGDPY9
T31w5G2oGc/dEzN+Z5Lt6pyoOHAuVwVV+NCArR9lpXGXXBUi1eSRzbIQ17+XJL3w
Dka6r8t4ea4yNZMkOoC1E5fmQveabm2DrPXpvJnsedP801yL7AaIBk8reP4mg9iC
qZky8KcFxln7Mkd3Y4ARbw8utEjmhhcl+bf92MQrCbHFKomQeiCVIH9chWGogEAP
aGpwxMWhRgEnh9Pil+kTlGURyUYaB/GjcabwaQC7e37kLjsJN/2EMNHfoQX7FwVs
q9f6+AYYPyp3DheXkT7pwkLvBVM0j6X33sLeTJnxKjOZQKKOuiCwOl5jacTS5vTS
ApDm666xJ920P0y62AadClnzxtZXLn3z5IelUlLIxwSeCUVoQsbsDJM17ysOhl1C
dB7q3t9+R/ZGl6A2p3JtjrdLW9xmygbI/bmchb6/yCoNuhWFzXOud0kO5bPzHqvW
YNEo+U8zwufdM57yG2a3Ku3Eh1jk6J4EWF1BVUmmx6AVVGPCme/cErutx+bOtMY1
2JrHgAMTk8WX6o+1L0B1wCVGV73YpFwEkido8ED21lXj3//IGaeNxc7I9x2REkst
cQhXdbLzqwc1oQOpMlLof93sV9K1rAk3SqmjjppwaMEzAZ1+rxhZR1wwPZ31xzck
2fINXYId2IToMhPFBnUq5EkB8TJpMRekvKzUqhvQ78vWpYw/vhTh7GApZwVqRDwy
ePSok7eudDezMvM40bYaBBU8+XqBjlvlUqGeLgE6OpnkXaumjzd3DZzulPpUqDF5
ccwJOSRh4gtJhRHBIEWrSX7156TO6QlLar7DawJzEIe4T4AK3zHKvL+RBs61BZQ7
ylMaecIGEaF81gB2z2s2X6tVXIy3TSTtkxu7atmpOFBriI9U4dIxmXNas8QksTEa
Dv8VcsIPvJFkc5kiueBhMskiiiv/RkY5BZN1zCNoqLRF9/g6DDHBiUNnkj4MN0Z5
Ud3DHhbw4yVNcoHjqIPfuW8Hb3d97QuEmr7n2IaRLI9dwsvd0sGXPGu5FbqECY0N
dpDSajMz4oi0y0DzPg1lGIVbYgK8fUN+vgL9yV1e13xC/M7tFhJzVA1BZorMA1Sq
nKpp+EWK3aO1Cuw77NsI+XKazuCPVsoc90y2/ppGkxHziQpnUxoI1cmhwxqhSqPq
Y3roCr2UFUtpMbVsJwvfIeNQvjLNNer6C5mseVS5Ea978mEVZZdfrdNOnSdaASZO
DdoO0PrSIpXFCOLXINzVRapJ15fe0bFscBZ87Gf5WaCzmFpxQKp9b5IV8QlMH+T3
kqnde6vKhbJkrD1GXqhG/zA5g6bzUj0wMlzGlewN0/Y0xPySeMh1wvM+3jTqoqbc
uhiVID/q2/gbKfh2c123wAnVpn/yXij1rsfPlHhw0rnetjHXdvg0aB/Q+uYjoCpO
AtZIVH8xaVXZ1EZtHllNf4IvDTM4K9A+QdcGft90AayrUdibAyyag5Mb6/H3ItWa
kMAYivv0cstIcLV4/PupNAHof91Zq5O5Dr2jGOWDTFkF2wbL0jmWVZp9XPA8BJhf
lMmNTHj96cqhbI/7Hpjdketz0egRVbdngi3sthLvPwdJwAuAecaUHH52+KiEW/Hg
DP/b2y6xQaxK1P11D4/RfshI+FQuB7QJFixo4xEHuJwMz0QcvkBoBZhDnf84Rzo9
vvGCiNCh3YXzrZep66TIN0d0v7zTxarCJd2h9NdBLd7HsVlHXSqV0twMwx0vwdcx
g/lHOmfJJXU1AtX0wyBgnJ/9Kpwj2irth7xV4N3rSlnnzSavYfbAeRxhd1xOTuRZ
+2HN3eyLsywC8T8uo9nmgDHbqzEKqrIHZWLpiBjG8nASR9IavNae2PVBuLYgRvJJ
sOFzhOzy9yAL1oL+kAztTs3QfjqDptmFaf+ny5xjZEG0nq2pqDxgdKdN5NQr6diE
8f/ZTFd7qFaUXvuKbsY8jb9SO0DJq49GULsYGVpIMnZf9QOKX19KkK9vwx6GUF/N
Yuz+XsMBCbSnvz5W16oUY9c9Ey2ISvJVUuHjHjLUNkkg3OzlKLzecLhVFy9RClig
WeaMjcrkLkIQjqMnXa9opvNOl6MJzVx11GYDHMv4xyRU6jCn3kbVlGd0vb4NvnTm
rNuJLa90SL2GkKQnGqf0WnFVA51ecvtWk5hkAGkAGzrLHXEDD07/gN2hEnF8PG6c
s0njik36qsKJeVVTHRMBn4EwI4jri0r3yG/uIFxjCL7KSIi/mYbDB9cHUAJHDpQ0
jhEIF+l2Div8mHsZcqfa3709EWD86arO2kw6GqJdEbxUjxCiVWd4yoNvhdQX+FzX
niq7jYL9P1aXkBBil2+ZDie++XN5f3CVbmvJDyOfaBm0J4i8Z9Vax1EISlFlQ8jV
3J5kv5LKrS126KCa+2p5x+Wprc2eF07fNc+St/VfD7kjYZJYuYa62TYfWRYLzoMg
OZ4uJivOdJAqt6rIj3MUgZ3FbDfN2Lc59Ke1gTdd6fved8e3JQxoEPZp31rbu4MU
lv3k7fgtJg2dA0Qcg2bdQS6heEe9aFuhXhU7JF5Fsilb2srDXFOBAS8nNJ4p5lJj
fjB15WE8G5HEBk7UvQI2DHG6gVTWcKS6KLGMlSTo/5erZmVq0mPicI1u0lRXYDth
UqM0ai76srZHg6pxZvKoHFX26qrLL+0LFohlLIvhxCriJIfK3mr/cli/ez/LTVsz
jnshasHtSWle6US4Pl+x49yQ3r/R8pmsv+CLhgcO5zNMJLPhaM2MDWJmAvI7DTx5
ZGBiULDzdyztxYYooDXwmyFFc0gyeFLMvLoT6SyyjUVbu+eNkbJknxXzX8M40Znb
+Hd5WDsX9+NouqS54er3WHisPwVHPBFnZ41NaE1otI7xpjADzseEiSOcGCnp4kMf
siZtvBD0N0RJorXdqXS2SgPwJSprA13sjcLmS8J/oanL/AX8eW/UOL3oMKOflmt/
xyuAe1eUFSek0fYlpqFwPVadfS5RydMcAqbeFNQRfiZXnyYyRXKBP+/hDfMd7qA7
wvKUlfNG7/05lJzCSxAXDQT0bwM6CNQWZ6DZ59Ju7vUaNEVWGL8SlWOmsr9qcVPR
cuQ6FFHEwSeHah9Gx/bQP9JBj8QOW4OkimevwGuVFS0MB6/TRM2uUyfrYgs85NwX
sn4xUmaEkWX8y0wxDnd9ohyX2vuPx9bs7OoA7c1ap5fKeVXMunNnzLsUvjKZlBOt
OBLeAeVhNLjs6VS/km5mcpKRcNyFAiklSzc2HuOII7Lb1qw2NzASCCxlaZoYFjTb
+YIxgeRcWe4z9B6jbJLOdL7QtPvjsgYfMNfYAzAoCfH7zm/kruAcdVKe4lD085nM
KHKDxJYGzxxX8DoLXKp+VxsXFsjnJmXAuMZ6x+DMrEufHFaUQqOxTN2UKYcrzLLn
gQ4uy+WzzJEHlXb/38NhYk0bT+mNKhjlgHuOujlxe5Xn/hEtE+iohGn5yKCRQcv8
0Z2AqphCl1PMQUrl98e8xqzdwMsLKpLzg8lsGUdDibXC0mRcFCj+ksgiz2LKCjXc
FnedHXj25brchitvLeicr4Ad5lHwYtG4Fq6xmXKpocNdPbbSgfe8ab1KoWdiO3Gr
a8F+isvX6ot5w8Shjmb7sLSMjB4NaMaublnrJINBKBElT/dl6qVXXpy3xOB4M+Jw
+UjTlwXmgTaGoXLC9SCDGkWro0wm7XdH8rh/xzLcoWB6SdY9n/4s3pxxFDC0ujg+
pfyl6qMJ7FWIFJfALF9I+i879i8c+KyD4xaK/lSCD2L1o5VA/ZMoirAzseRBGmj5
n69ZRbZ3yhuFLsBLi9M4rQmsiPab543qclnn3JVKc8RrkWtX4YF9xUWU6RmNLu0j
rdiXaF+19ixEQAaUWSy11eQUzmH0Zqbcx5ugzW4npA1f2Js+D0x5K6jR3UF6bdPo
EFk/CcZiHHjTR8Hk3NTkUOKucW8cyCJeJypsfpuszKRKslFkwzjFhMgMqk9DHouA
ZYQcyZT+XtfNtocTHi1iaimamBg7q4T+GGzWPw9NcicZ2eEYZC7QqX/DhnT7TpiG
7boD7+iZ24E2GeY2Pn+zSa2WPUqiEDfZ3oi82X0r+1TA1JShlDkem6QyMpj9Ii2/
R8f+TH9lrMqwN9oMFoxhMdl0h7hXIfUoj7FI3zhisZQdf+T+b8Mx62lINN8G1Usu
3rrs6YF929oZ/x/q/8HGDvao4S1G+VEqE6eTyhbng9ewq2sZm36oRJ/a/KSNzXx5
cMkct3kwGOMknguyOo5ehUusf5GlflyMKs4kLC5wJUwh6IMll4eMPSr3nZyB/6+f
H0WhkOBmTTpdOU9K6RBTAg0Aapd0r1JVqaFUeohe6fdWQkHrJtaAtmSW/SmDs/13
JvSaAw2C/pUByp9f5msfux10gR3CwhsImebOTbCycTdHFCahN7PEcs2KS2mx+x19
as1dWjAF6jCf+GjaqXd73d1fANX1wXIV6KwyLt5ZoMa6xTrtp/3b14pwtYDyZcVE
BVNhIlpfAfirQgTBpRpP55KQU2/2GLHbGCZO+sCOeA/5CT31B447BReOVPYjCuH0
cQaf1E3FPq4nQHTY5PtGJ9rzqRYqIqv14fA/64HYGeNnppGUdKvV2ITEKzwPt9FP
lwjwh/ibrRxO1+ydJaROIRAbtayVAzNLslQ/GavGNy71DjOIr5J4HxD43NT2355V
DrrEd9+4ClAPE9D1IwVqEe6/zVqKe51GFQt4KyGd8YDfjp3RMA5orPLUV1dRaF6Z
CF/8Z6aMZGD3fJZiUw8TDawkjycRh1U+Es5+PoeNq/wfL3QI5cYXrmIIp/Jar2qk
p5FxfuGnzV5FnHS+TVCIMsmKRocoXUui6dTkBqPSlxB+RBu2bgOqzmAVCMTsnTpw
1P026xh+oGichnscWLRqCioPlcDgwqHNeYxobnB8Ky4f7ycqQUgwUH6AEIXPfhRm
9FlctRGYvTopFaPWLL/RJC7tbz/6JJd7oeHORi5lFZqO5jMLGIBYMrcbz7UTfbNX
nHSe0uLlb1xpd4Zwx+nVDYkpnYz3OLEAVY8jb0HcgmdEPmLFI04UCnLtzueSqRVi
9aBetlghQdjhc35YamhksI9vOdwc8f6AQm5FfzoAadPOW8ZPjx4lPPK61lK5NIx/
NEOtQCNmfkUAod9yjISSlYx/aPpX8ObuvVVOSJ0ehLYqvFM1xjo0O8ckKZOatFGd
jgJGq4+JCsfAlC5pa+tubE7VF1oQ7/HQi1IhJGj2UFpedE2MKhAPVMQAIJFVZjW4
Qci6UGJrKGW70w8wduxswN9uQjjbi737UD/mqYXGgrk8fYVYXSerUPMiy/lPsomt
RDF2A7JcuwcaFML6fKepeiiGi+GFLitQtvCxDvRedI60o5zvbmpWdt32gcffQ244
2Qe1l5znLoomMllhweg7yz90Ytjf18YvkBVObiIkOMgykesgcPTj4nXGveAGc3N6
fmMGTwzF13tOhuUFs06uGMH5LLbe1FjdLt7HNNieamoaI2nqlXC1JFrTZf5FpDID
xCXDNJ4SgQP3NB1ebAD5c1ssEXm7UwznmCVd//VYqd+NZByXl97R+bQZa/AvNA+B
um/8vRizN0XP3L7NOGChw6dJYV5BKJZzrWzxaEtP1dRTxcyLIHWIq3p6DdhaB1fz
KBfwq1wAVJdm3U41WjEvX4EQqkYXszVnrWVXFdYHW5p2iPmCDk/ecc2S15seguJ2
hV6IpA/PNp3R5jVicvd271vumCEHQ+aRgHLD0fgxOT0QMB1oQmZAVaw20tIC1I17
tY0BKkunxMXQOzD6gNKoSP8diHM2yoha86xHZw7gAI2glI7WMBcwz5VQ8Onw75jS
NDEAMxYtnr1ygSWJlMpAK7V8ihOxDnLIlplZqmJgv8n1SmyErcqrJBTKnxxk49Z5
VhhZxCp2M6+wcDJjHxvMgEJ6cS1EfW4Aiql7H49WDtv5osG/9WZlciYlauJkeMIq
E/QhWA1tKbWW/8NxloORPPqAE1jo3Od1NMi699irvxsvZbuhIjuC5fJ72ZdLrVY4
qxwkhSw6cETOR6mg8asx6ijIAqamLM+qtUamf7sqnSPbk4caN83ptixajZfQKJpg
70fH4RlOclURR5j5h1Z2UsNQCtIOGahvACCdk6O62fuwZ1LOzTza/jrwTShtlq9Z
BeuVKCQzDo53BJJlHT+buTFvdABjiAkSkIPaFjODCw678+W5uyaxDXSPhnkfaq4h
3s6+09Zz9RWZStBTDxXjoWdNtYpHus4jr51H9o5TEOF37T4JQHJlJpjJR/hhImkM
qJklZzAagXIwD00Zkvp+3X02u1v/DhwcLNi1QhPpoFDiJvOTnkKPjwQ41O9hJgLD
bHOryVA9mT1K2hfmQAGBAEO8am5bQGxNz45VkhftUasDxduyU06tjF+N5aCoBWvL
N1sFL7jjnUP0Otf6aOn62/FfmuYRup4+Ob+P+6aagpsr26g38nlCi9GhUzF7J43N
7E/tU0OjJZAcknxBCbjyj7lMEL/Zvbf6jPRwIPBa+sqvFpuFYKpDRAEa3lfqcTRF
0yl11WmUvZlXLCMlyVXF0MLdVx/Eo0B9+gEPckd8RzWoouu/0j0heCgPhx0K4ynE
3luK1bK/4GrWoplk13ZFxYTwfC4gP6eaCMAUVClcbDiw9IxPAV76Uyclhw8dWdsW
vQp4+q08bJST9/gUoSqgEdyL5zfNkqR2YPui2gsCAY9GEDfPsYnefvKfY95VC15/
6w8ZFN5TLIa3R/4UwFWyOEeZrpb4jKNEZYlYMQDfhd4ETK9xoPgNVeC2vnHIAzdx
xddJWGMA5jzS1D4/K+QOI+/xZD5ywog3eVJjGRatx64OK8irNsoC7H1LFbflL/t5
HeMbnO4Qb0X9xnPv11nRbbyWb/jBFeAjfsrglwQCV0M1bD6+gEjvlJqVowTJia8Q
gJCHNMopvkqu5R4AcxB1mSf+QS1EzSSIQOq8UihN7NtzE7L0krLHRXpLTvaJZYfM
O4PXkngst5cW1+UDI3zAvmlAxBSZLjoFbggFFERL/QyqBCJpJorpB5Vtb/qjBjv/
RJ6jNY4owqnyhbamziQpTpsfErCvTM7IDl127TWLanAxZzkgEJpqub41V0XraxxF
gqJRU6x8S43U+PONMphUj9UpXfxSRpSAYBRI4zR0qwZEIPl5BWGfncbiAzcZnGON
yA7/PaRiA/a24+0who+7y6ZMroVxt9mOOIrqtR3KRnuTsyeWeqJF7I3ZokwK9cWk
9CEi8PUWiV792yI9jKsiYXbvm0Ht4zdBAeoZp5l9nCu07YyT3nSFxlbKEPQH4jVg
gd8fy4XgM7JeA1QAa0CKmYyt4cyKv8IleY3XxQCuSyAsy3doQm3OJt/Ltb8wFPRw
r48mIiBY83/goCzF1u8jMPekRcRqofNU/SzOoaiz1fCKgPtvDfPxKgKJioPRi5sS
DfJeI067FEsyTanlxPQjoSf0f1btw4s8rl8rPm/iM/KbJNfuZrRsj7dnNVRXWMGu
2Ak1qLV4o6QZbfXR09CRBlD0lYzqVSOmdezoWXz88/LpB+DJKpAz7mGKyXpYFgJO
nZ874kv3rqZECuEBA29rG3Hv3QFGYMzP6xYaue7r+RrCJVCXkZC5vwG/R3a8OfTM
3441gWWbM1Eg1iWOzj4kw2642Dp9YYJgOJamKGkSaH00dBy0OA70WLyByIYNB8VA
rWGnkTdNql7vQFLKOz5CL3xSCXk8pZ6nhzxOauZSIv2lrHYeYNRNuO2b0PT7TwSR
J21V4eJR6BSjtUm3d3RagRRSWUccnHm2XYdJXNmsZwCs55oQLKbvSSc47BuRZe0P
YedjRi5HAJzhp65JdUcSGnwclW54vSNMyRCi3eBOks2Gfd5l2KwQ6StIeUb/nBiL
F5uFfQldTsVAPFR/ACtt/DzjwzcfDT26KB9zDnZMyDHdiwo+zaVLIV96L4jIxZDJ
dArZpmpVfvtN8+uNXNmVXzsf1WraJT6gYJyw+UMVjMaIUvNR/o2fJ5xiIwPXUs0K
IcuyqoR9oworU3bpWfF3q1ab2utrwEWwbK+E8nEknCyUYQ9KHPsKpf/OAo0ZJahz
U62j1IL8hrSc8u5DZJfRvuFaoGGB7IZgVVEG2ig9E0RNG9T/feHoqSrQuEaz5J0Y
uKzZG0LMdUqTsqUiGa2zJu6Sc2u3lydnij+GO8NZJ52PjvR/QeIVU1X3doNTAnu5
3P8+qNfGj30qnRRFZykeMlZn49PizVw1qa/ZsDYzBoZKJBrZltlDpO6amU6WBDlv
nyBhj4bXe4ekF1+04atVoEvB+pDQCwBkB8bwSeIZ0DwH43nzrFbaoa6pkrArgR41
eUme3IWNI9Oy3JaVdSf/DO7TwWZEOsM1p3KS/DGABcxHw8j5BHjQq1EWjghrIgw9
d3MHRnkyp9ocM+ZvK80L1BZJviBdE7T988qWbNeFmk6y1Md9sDcIENU9ijaluQXW
4MIneMLdr1PSUN2teCOxmDrgqtdS66mYkqv/kIU0ZBbdcQYWvLx2gKnV+FSa4W4P
rrkk+BFSBxXIzpK4QPRMGLLi8R0d332JpqOUc/zi2Qu09rlBr335npADoSEMD5Rn
evHrg7Y1a/7HTUNMLxUR0uldHJ5NUYNWVKrVFecwaa6NsPTJl9odtK0mPq9kc45s
ElYD0GfHClGCV5Fyjx2p9rFvTPi7J9sTXqwuchsMyVdRhES9YByKbHB8nBWiCm7C
t7WOEK9CUK8Lw3xs7tLslROHAZr4kw8aYAUwMb3aBkmnKTFSLf/u600wFcp1VYam
jkrQAKkC5Upu2tAsKuv+rz0dZA6kzKa+yOrFvrGC7PqrFcssGyZdU2z8IunNwxSn
9H7g9o+P79i/t42ihXxgKtiE1AWvB87e2jC3D2B9JCPcgYUlVxvRnvKj/HLVqUoO
ABjyxfJfF2fmlvTGqCoxdPnyKKKPyLExIDvy9ppCau1unufeZXRvPp+LCo4AMtvN
0quU78SrZO5E+N+Lz/i0JuErCpE/tdTpBUQ4kq1g/EU3G9gK7Jq0xgtaQoN6asz2
vrQG+mWc0xiKBFLYTVhrLW/KAY3qc5AmtMfZT4cD9Jv9nH/tjhUDhdd1INjiFp4P
zgM6klvNvRnpBZxj85vQ8QB1pZXxGfyBKduuu6ngn5WaqmFYJHfCddYYyKHVCLNL
jYJ/hhboThJJg3xsYOzAErX3rr6zldzHhN07shzqOtQM5fNOH0702w6rQTI6Dygh
2vo5quOpKYUS571Pml6UlhfsxAaGzbJ47ne+z8wkelrpBCp0+YFi3gLYlMnTxyoc
bsX+29uxr21urf7sIpLuO8flWVndQ2HkoYT1h3d+0QYPqF7BbD2Zh4J+pOBvaFV7
F+EfPiMm9qghUEGBNlE4GvdBc9i4uPpvRAWWMgJUCF7wQUbdigFup9ZwlnoZadCs
1rJ6C+k3W7wcp2hP1E9Crl4D/I9ONo9CYAO8/I5U6YxQxf3Hk3giD78v2AuzlVse
R7BpcIlENtndOZEKYt8sHzKsAB2ff2GcYlueXWm7Fdg9m1vIPeQwrPP7YjExqIkR
7W5UkvED0nHCwI3iiBKjHleknj0Uwp7HFaDBXTN9ZiLNvFwheteoY8lCYsr+KBCW
E8uUlf2BxHfWw36VsRSpqlW3SbKMcywyUDmj7PLGq7go9ZMLcPb60hFmHhJzz0rO
wNs3pRBEQ1mUr83ipJbqLicLfUKW1hrpaqHwtkqJMGo99KSqijKIlhiozo+wHhJn
3EPk23sKzR9F8qShIDhPvsYr6FQJXOoSePLZWfIquWzqof3t8P8BrLvCyVMmZ+bx
XAk3TgJcHlziabIbl/Ktl5BEJo9WIU2PIxr/28sNq1CwoHpP5HGMezRE+0OiWZXn
Fw4zKmwV1lY8islATSr7C4tpnx4sCRGUYVfnv/PO5QjEBOASKLIe9or8UKnxdBH+
XlO+aiCiPw2P1LVTJyN2QMoOIQNw784uX1ZR8OD7MiFC9hoQX8hZ+qawDufxmn1b
ebTZWS6PV5mh3N0I58AP2iclz8DESAUk//o5peHFFXdcMs0cNLRrM0uLWMZj/Pzd
CWgFNRm7Fa5ESvdeY8UFEMLfZpyvwz/DEX7lNTp6zCO4DpPG+1+cUnzPqfFJJHM9
nV/ClrfpM1hDLut4oNaDEP/Q+yCH3IzQkejyhmAHV1SPFNdvU3asmYhGpwHQQLIy
Jo46LsAUDIJtk5oWgXeivdCblDc+3+uuV2gXsUeMxqlik0nzmgaKDu9Kod8AzyDv
NXobog13VpRYkR6orLG9j4IC5/x/eckw5WSSqm+TM7dH6Yje5ionYbJf0f5qGVMG
TmSKIZiQLzHXqosLayXTiPLgGZqMD2AaZAMNMoWyxaYBOuLyz+GaxgT4N1jFA/Nj
493J/9/str1XJfxEhBdu900qQATYhcBVMX7x7aDP5KO62w/UVyhiHqu+/+TQ1kgw
rysWw33rQTxpElJPmaQk3fI3eb5kdz33QghJL751FkDarfe9ieu4JMNA0W6JsH3M
uPyl2CKWMyNYSUfSSIvDLzioQPGdjQ0uIYNU82y5sBw3TXKc9TPNQwMaTmfuKkj1
UJd4W/TxqYT+aMj3iW0Gx8hhAeYOvujYx59o7/ObJ0RKsN5pk0NOGKoHK4cKKm6b
sZHQj8yi7V50dWn21SSjOCF4W3DhxIRbK71EUx2gufYWdEi1YV+K8Hq6kHagzPBv
xW2x/o/eCZ3EMx6T0V759CuQ5tnb3AIkA/bGWNuvaG+H+xqHQ45ArQp3ZlUXQSA1
/JdY/bOwwpTtK5VoLvCBVsPV4bHZOlWLH9PudamJ3c5fAkUxdMAtNCbTKSffn+wu
ACpVAVI1IGF9n5gUiqDuJh5NENZ/njdaHIC3Y7XNbNSVI3TqyZuUCud6GCUZm35Y
sbKi3PQ0TDcxvh8MOmqdjaXxxzaK19PQwgFDaPziBx7uI7NVNTBO/IIpu9JEnRYA
/2VAMm+syxKYdLNVlvS+neSOrr0yJfuMwffnL8Y8rnsUppieohw/yZjQt14Da6gM
gXouZVHJPmgLIBOnXSWPjqCddpDrFuBKI6W/N9RYgz+arqrZ42rvaoEAN5uRlmRP
jPzKCAG5a59/GCVB40jUrmYrdKZqg1UdcIVEaWx7N4QQrrmHCIo0+VA6S7bSZ0y/
FbKvD+MIlJ7MqMnS4gz9nGvqpuQu21GyVmDh+c9jeu4TAPikVm4UT9FbX+GpnVOC
LaL2gz7gzuAysmoMRjvPEr5SXIz0dK3rHo9+Nnx9J+50qgL8xjx+fg/lQYxaxUXa
phJ6W/Dx9cOcBhLWNnkbkrNnUKBm4QPPZn5uj62CAXC+Krd/how4z4e2k6xNhqOH
5nn4KCOO68TlLZb0S03ZrIVevQyKDZYtN2vGheocwnLVFWT4KWCdUhORRNWjVdap
iJmTT1DxkeGsVkf5DO/UrkkVeq/Ae4Zk5ar+P/vLAIAo7o25ixkrrdihi6MbU4e6
XL8YUjYA4PtHeOn0evKSYEQxKMAfs3hbbWy/VhFpMhy//GVdzrR/rfLZWnobwMCs
QH1rqym1Tj+jOPMN1oa9mcRezvWn0Bt7n9esKZIdZqTdY2vOq+pbfNhEjxEFT0FT
gExUCZkymsVEm86OxiGVnHbpurJk+MQTzG0Hsd7zyCrAKonS935P9tzBO709phmz
5XS+htFNcZR15c+e7Qp9KbWsaEFu2eAXm+0bjMYXSek1n+Q2Va/A1LM6SNZ+VsKE
lBEwBVaM+GaFsN7Xht1tfx1FhZo0vRFYrreITpE1ySYEaY9SAw5eV2bbLv3rho8L
IndqzfYrK4Evj3tDGDrN52YqTi8fOpHZF8v2WR0Z1jQZpa6z+ZvR9UTClzenMQlg
YjIEcZzKCFDiRRVvQNqFJNKMu5xYhf+gWngJIzPRBNNZJIG/A91vqM4raf4Vf2Lx
chI1NaiCIGgw/yNLZkorcJun1GB3fPI5FGlE7m9uKiJGcCzzIsn1sk16rH8Qd/BE
bhG+dcYtPrrsYkF9rwwBXFQ37qEpvWGO3zVtgzMmPAPjy0AplCnygBL1rGjCE0wh
ur8fIk8Qhg8JZLiOpXctYyScCVvC9ZfWEn38XDLIu9fwe/obWwbQ23mYv4I0Y2Lx
XhuMWI7no/P5NN8Va0rl1i0jwcOo5QR5+hWUNWHxXDV0xKM9hp4S5T0Gevce8qOG
kOjvlayo2yh6+rlt91MvRv2g48KBhlvL3EeuWmP9+2u7CHMLhoS/0TI0uYss3FWs
jiCp1XAT7jUAmfvTaV8Il/Hx+zPjT52GmjRXB+omI/zorF6cT3qReQNVr9WAmIxr
xiWW+Un4QvOOQY4hQ4ceTkEA+P9x5dKx/rrLrR70P/KY27S1CHd2dwGvGErhFXzM
zUQ5y4f7tWV4X9t+CKb6P99Gy5o6XeIMZqRJZttyeYcgtj31t8/liN4XSYMOlgtx
8z1cpRCvElii8LbWcDtyv2J95p9ZH8ZVTdw48ELIHAS5ZdalAQ3XpPsqzEq/mRex
wFEBVzi+CmQcHmEJXL6MNqK5Ft8sB2uw4nIB9EzaF6lJCdoWr5NPf9q1Q/vVJFOp
cQCbNoLjYFSslp55xzT0AEHVrNYz3JWL81XyCc5CIs32fpj20+ETIlzWVhIitJUN
l4GmA032E8RXeBs006viI6T/zQyVBoT1X0dnvR8LetLjiN1T909ELqCrtEEbbV3T
jyeF7kpgaMZnYrcny+9NaiMd0UcelV10Ybz2+EPCu1vs2SnIJdsjlJYGUkn3DViO
ocn1thhDVlBjnAi7NrYdeMS0Jx53cRtcR9z7+sUBndf5CEQ7P0FjA8V+XEOsEu0T
Jx9CcIyhS/EIifUXAHCaIQ4Q2kKpqaTB+zpYzqZgiF23pV+VMK1aHrTZ1f0nNb9B
J9i+ANzMFMwtkoAhJVZcOQRefxZDbSqZ/QuA0kg1edocUo3fTQqdHa+jnTnXcuci
ARVDVih9y4fiH2KsB2ZOTMLSr/v4puNCaqbqXq2+7BVLW/TNgOZ0F3MiC1NZa23O
nBkXZbHmwVtSwV+sfkct4TaSG3nWvPuvfAWNX/5DH6dLR9UjX70CxZBA9WTjuyw3
Tj79YwjDW/9Ls6Lq/vT5vEzXASfRZSrPgUwQLgBSlT9jYOxIQAGqa/pzRzZac9Zh
7x20+BS280XE8Rq1N5TNnLMGgEFjx3nkGspon6ud2VJEJBbjWZh4SdjJp98x8MaR
mR+0t0uBiq+vDbLLuUjBjquEU3TAzVzXb6/hkKPwHe5MQgch47ci/lOxxiTrkeFS
kZE4TMRwIf4xQ8qVlgoFSVC4JcoJjMw8YaZXkN4L6sjdsGWRpK7gVG6e/TiwyhIg
H26iNL3UXzOz18lRRoNsq5i9PXpUh/mDuXrpLnxnaEwPkxyRHBLSgZp+Ln84mlPy
bZv4R+Ww2+K9pr09oTf0CqGXEc84qkeHtO2BkT83QNnL5ryFNKU04k7IPkKrxhVo
9c87aEi3Mn5nF3RzrrziZjkA9NKB31eqfimh87CAku9l5shnLgZCzyvTZ3oCMSqb
Mj9GOlZ5lioFlJhOJAYRn8X+zLmDHhORUkREbofAPA1jcaNMRjg9EiAQFP+IpixT
t1rtIRFWNnRbkbANmcKV/x0lHqeT7FiZPjHF+/WXebjZlNuf1w/33DSaXE/0zQFf
iIp756qGfThoIHNtUqT4ivKakvd2vjApD3z/2sEp/4wjYOkvSnlz/LZtog5gjJND
zC6APdDJKOlkX7uJ0Rv/NlNbw6D/n83SmKnS/8LUdR5ZvUFr73fvKsKyuTHercVw
XMzJnEtS/1Mh+fWH7FDDcGEwUPuwZfk3u07ifZ8wLqzmYqlFZtnAHFD1AAwn4dHK
aM4sU0VXsjCon10E3xWSLbMZ8z7JvfkNRxOiMTkbNidWxmQKoL7rBrzgcV7XCa6h
dg2CPoQn5QDcgj17Qyk29dzdGp/vCE0ynYsx+y1nSh4Bj6T1OTnutl2QW46vt90p
AKrD0WvHQwVWnjHJ5wzOPdaYQ+73RWpxQD7BgIHyX9wTODWSABYQxijA6uHo2IiV
P343T9+h4mfr+QHlDvuzVDZyJ9Y36LBpmHrOvGxlBXNsU65Js2bHKUMB+E9e5e/B
5lCZzO/K5vwuDyE0RD+697CcKOv5z1ZY60ELxmaIN8JwPldbYUPBBncyJ8u4Fxqe
742rr0KhGgQszpZc//nICN/NHFG6Bn9jAuOKm4x+qb+F+/fXwTd6D6lXgWUq3Enp
mS87jjpDvCj523QShO1HXtN7XZ0rcOkqONsOhNUvCEswHGeXDBXztX0Y4cpB5sTY
jpNf8Zuj+YzTPh46o8npQFTymaZ0pGW/S4ZmHIZs0EVxI24o76FRPqB6WaLfiYEV
ye/WjJS1lCwLPTGEjTA6qQ1BOLv7j9cyWhbhvaef5fUwSS2OPvnFW26vBWkPIhpU
H1xfk9dzxbzmkc4qozBOrjLMeCdtYugmawCS7KZz+WGHx7kIKvCgdOp2vUH6DXGN
6XdtbdoaxUbWnnAC7lmUtPampgyLtz1slEznJcrEI/rmNK5ey/bE1MOnDLrQalO4
MuivBkwTyeq7iPZUhJam3xapI2qgh4ckoClSLRRyJImgIeB5Fq2+C/EgzJQAnwfK
uzakuSJ7USq2sHEi+DhNA02bRt3tNr5EcKu3TqnHDtt6y9VGAgWoS8jQGkg6thnx
2HmI6K9Qy1uIxPMAtefePt72tYDa3UCeN0CBkR8j5JLzbHRWh50RhfL1EYBYU5hG
CHgYlGTUybpZcAorCr7JvNLqLi4NBpZivhkcKhe3vJIe11nTFpafoNVJDGFYtfxE
G59LBnUp0csO/8B4Kv48SuWihmZ+8tOQu26O2NpVAkK0AkDkMpkx/Ty+jJ8JigsR
LJ8NNgdHrdPM9JEpVMoBM6TcnjcwIGpbQ12+Srphx4KOS1CDohMRmzZXOQD5b1hT
b3JNy1KszDLHe3sNjAALGbfGZKjMdbRV6gwPu2jItDHRmXWq9Lk6oo1khPJMJaS3
TmDn6ReuuJpIaK9ampaTvWkmwm6aaReCyLbPdUMPvN9p8D+awlVhlM/YNhf4dQqu
zMiLmiuZ2jbd6QS2mxx43B5pgWNzHBj05f0MjA830OQJn36mxqp+h3dVBR/SQIby
C2PpTi1UMevfpbNmPcISxonNDkvTBTiWxi7vPpDBPT/Lqb/7H/ipbKq2u1Y9SKK7
sYRBM/5nuOnFke6WbqNc8Q4m+l8GkAL7yFo5UQLgvmWbvinHlxQyqckJW1S25+2C
1Db3HasqRIRPmRKhLvwvxp58zZB9aiK525PwX4s9uUTDu94DKeJIc1+H7BcIl9o1
yEfkUME8jid2F4DWQvda6D95JhzHSgxVPfJgMDsQQKukEMy02mF5/PmL8RFhQKwc
MXCIV/6nRbTuYZJ8pQa77K5aUl2A+J3+T+auibcYWsaJ3xr001tRwjBUmhEHrMIX
xhe5Qf9IKkMegiw3gm3AtFgrNiKaMZs7eTC0NTHeoLo+4fiyq5TE+3l7dPnCZihJ
OtmixNSCZWWzHiEwIIs5+1axepzYRIZ9ZF6vFMjvAbJJp56tjRaANRY6xt0G6Nhp
Eu9qqgIkUzVMJ7t0aT+HhEwSAehaAGRQyJEZeomGVcx+bWcC6QY9gkRCOffyzuKx
N21930wL8wCFF3rrZEgEx7Rl9WzHyrGuJtzT1HcRizY/RWEVes7Rga/i3QLZWjrO
8VUNQ/QZpzoXQ43xQtjyszhUtaeCFq3r1uWTii1dIPMHi+0mjT7EtsNUeZV8G0r/
1+fDStpwTlNG13zdKWiin/+nF3ItaQQMe6lObsbrtFPR4YgSzo67iZE7enkIVjO9
7DoISwr29o9uAzA/JfMESVzcvI52Yu1hmxsktKEUukfN9x0OGPjISraxaajWlQ8x
hlX6mzgRV6OkdzjZGE3+g82KEG9kOmqyNXh1WUV4qpaemCZ6YEauCMtev24k3GbS
tt7viaw5lm2kPe9kohBsVA6yrgoDUaw+wmy8E0XGaQBtrX//UGPskODfim2tV03+
w6mmZZ0kGuS6G22tux/Y1zrPi56AQxM7H1GvZ9Zrw0AWyZonJVHKASZsnOsIWZSt
qnGIaH7rI9vuWJcIELqyQ1ELBCT1wiozqPW83A9TxCZXJ/Cn4lqTE7Ia6qS/NxZC
3Z56AQ9bBN1u3IpSU3vdHJ1YP02+TZt4wY4MTTxqe9F1dSdqg7NY32kpSzAnNetf
9i5gG5PEhd6sg8BTNQmSq2Wf+j7Z1fJHSAPH5QiO/UXVtz8pAVIUA+OfAJwl363y
j04eABofm19YHeajMFNiEpSPM4P0blNUCnn3hkEqMAH/Tj0BDBhIvIpjNUvzXR7k
Y+Fu2xP5bfL7Im7i5y24HN7Ke6WVmO8lrSyRbGfRemppkbm2O0Aib8YulIw6f5Wl
Ee+YrmPdKilLj/dMs0M8Yb8D/lva/3ur5GxqDSDjvO5QKbAt33MVOHHXKzz/3tqD
fXAOYfURga8dP9migFHuf892gxRj841UdWWgbkO7E9yiQ8RlNJV48K99bt/7FbVL
Qfv8tECo4gyG7PRey7AF6VNSDQjUSvBfn8Ozzuce7lyGXmJym1kPnAx+k4cekH9l
MWWwIQVxXLgUPC68pdqXveA0gU8K1d88asoMPs3JeWd4vUoWeKzlSBJYUXup5GJN
LVZUyJL4TlGQvDnY6zJxrbrqYzeszM1SO2Y83OSHJri2JspzHsiTiYa9ppgKSdkK
UG8lHToJ3oL1ArO1ToRbAGd+5AYAGfepkGGZG/oL8u10e2ZI70UcWwWRsoGTJfMq
ElxNA52BIXwQ7kgeDaa7/NrllhSe94qzQX1QMuIOc6mbs+sfVGYEWt5oeWsQDKGW
aN9EerSNI5iBakHRjowsG0VBy/gjD39i0Ys3SyW24V64GB1IstQDlTFReYydkZLZ
tLZXLreZ30uzpA+ajEd5LAtNONF5TqfNWuwMukHFxV4ZB+EzSlbNZ8AhIfcly4Rw
kowHXsfqQ7y4qMJ7ZFP1uD40ey+zXwSjE7HZa2ugKigxQ4xY1iN2T4EVQkatXifK
G10Nulgla4IvKn4rzGi4IGpqxZ/1LFbzfa28sacBpTlelJdF0eusubFp48Oc5DE4
X9+RXhEdpEFLuVaSejUHTWxeVU9jJkm3K2h667WwpcR4Jr8TwH5Q/RoMzzce2OZU
mArVoZ5dz/TPl0V6sGTWkMg0TrelcIoAcYTi0/PnbRmvhPxbJ9t+VfNgPlo3bT2V
2eu/lY/yrV2BBPb2cdLYf2Ragq0czAEMeWh4nhkSyMyO6Gp/6svTt2spr5e245pT
hze4UEPYhdgcE71z3mkav/iP+iAu10nuYVQ1Jat9cSmMg/tm4+l6sZOPyNX/jOWb
eqmjyp4IS6KXizgjMDCCseNyY4rPuXIDbZomAC5FKet9MXjHXKar/yNlJ1WtOEJj
BR5UfgqMoGSilSPR2+WrFLxjk+1RFF/WKTICYqBNQcxczj6cTkX3BQ3H6Ra/NIl0
xgFqzdwa/mjhSrdKgjjOipiVws7EvP/AAPddluGL06kaH1fS7ZG5rmtRyaIbCbae
ZA3m01J3zcB8UJaHfPIpbcULF5oq6914/+XsyLuXSPOG+ug65pLAfp7g2STCuEwU
/bZiwSJQq0KM/aBrRsradcv4kV4jrxeWsmjkwLocj2/gyfOMKTgSj3Mo+06hERUZ
cokzimNK+WyAD9tl6ecw1IYXq/6X4VQsmJK2UqfxfeW8k+1oWJQcrSe5RG7J2BDX
l9/0dIq+mkJO2AkuRDU7vWB4HdwILla0L1sb4u7QNnCE4gEDFnaycX+tanExUrDv
6qvxN2UFJo42gURglkUOPkLGAMYX3TmzaxyE3tf3OpR3fMD5TzMEcJWCBw9iGmpa
H1asFMEghyMM6LtGTmqtJ3iKKL2tBFPyvYXl6g7nU9Jcy3Hl/DvA3oXLOPibPfvH
CZ4RW/K/sBv1vHqZx259zK9LxZPnjKdCw/e0TWT0+JiX5EpozhukFnoYs75SjaBk
mKHlPAxrFpsU62aByLKTnWrKvTiRkUIMqBjq2dOeJ3rRnhUD4nw6g8U20Q7CfyyN
rNEoGn+OAe0OPof56By96uErf7J1nJLb+refYCCBHX/x5n8pHFb25Cuy/xfLwSbF
4lEz7+qcnorlT9oFqO4ucZ3A6DKmDe/FRHZ6x6oVeZeqYn1VT5DrFmhWmvg8S3FW
5rHLBIJP2205BL5XAug2BBVDELM7GpMqghAbXVpyoo+614Mx+U3wjM0KV3o58SEk
LLqLGH54d9j2B79xHmO30+xhkPMHFxBmUUtzHJQ5+lMlL5/LzjM1//SqbCK/3oHl
SIjgLmmVLRtuML8Qz6/2ikwki50Xe669mrSaMVo0wrJ4G4+CHpOmfdxZxLNGXX1f
/JhVIjI6IpuBWL0RLn3HStkOhZ2PFBuUyx9RsdRTt11MInpsAe9l1R2qJu9/PP5m
El1xR7HL+SO+Trr16PIPZ01hUfYBM2xr7P3jbV7/0BDvJEK5pt5j0OxFd353P3d9
0H0Mlm98m+wmDZCZt41OcUmHFKeiOeTEFy8E9NxDF6Dq7GVxiIeahrrMm5g60tvB
TiLf+bvv+LhqPz5BB95+VcX2nkKIOYE2KeoXunzwAzNgrkJA4hKCmxJ1qd+l1AuL
w79GzA/WkqXMgxyMLFKRT0rzCDc32ZDdG30XkZOEIVMQ+3vAjoG24C0lGfLEwxlV
ijDySXK0tB4gOM3407I821RY5mmwPE01O32T1KL84uYuJtZ9GfJ8KjV6R4paFx67
ed/3g28p8B/t4YdTZpSiuxWW4pqXaqsPmNVu7BqQuFECbRXx6+NCPBhNHscanc3F
TBckVHNGKngOCU7ckdufilkAELcMDZ2yi7ykk09BZs8jfzZKEJYJS8Bn0AJRJ0rB
zVj5lbj+sHXRN+loEkbeeP2MHkz8m8wRa5HEXHrbcIFKZ7RZgSCv5Tkr9vfQwr++
G10GAkwtTlYiZz/Jknb6XpSOElezB/KKQU/w9vDgNkLDLlszij53JzUxWtheTSak
Hr+ARTxpSMWr/mtaYqHfdDoRNl9Do1X4O9sN3nJtzDyKMtJ/OV0q0AWqpWKKSv/a
T1C7dmAvNLbX+rvRiWgdmwU6VLaJuL2det70d8AyPj/TUn2gPE0cx2EKj3FJ7TqV
BRyNgOKNduIk29UH7QeqjTIyxj89iCRjOM5b3WoO6JeLwOZQuXiLnfQQOcqlMcJj
A38xrwv64OQGEyQTlE/BXKiQgBOE6ksKbJVzdmOsv7F1Q32rGsxYmlXWkb4AY76w
IHm+fqZiqM24PvgHvyLm17xmXT7SvLUTWA+QGKftBtezgqJZ+kyZyN7s0EssBsbF
bkTLzLGn4frAFKQtXIb6syhX/tmT7CF76zLfE54qbO3yrHWvgCxzj20l6swh++gH
lpA5FAeRJ1RwXY8ad2Zd/35AglBSzlj73WFlc4Xs8DH/I3yXBEYxPyyjmHJJz45U
9o7pP9izOjoT3TTGt7NwhnuM35Ils4xUSp+TII77P6+qtdYolgS91y29TOcQgxAb
bTSKcEWbDfzYe/Z3Lo18zaDBa9VXTSFf8c7PYiWmB9hGn7qdYBas9agyBuqZoD68
lVuI+qSWcX9LWjdZneYSLWUtnfu1AIO6YAf89BBN1Yy3yYw9pGBtrp/5czlc1067
OVo1EqOpfuWnxjgBbDbR5J0UhsbID67/Gr1s5pI9AihEvrzTAaIIJc1KWyTVgVnC
eI9UJLNyI77/WSeYIRKaxHtukWjIxjIHONmo4DWKiE/fe4KBNpcN7Cb1gPzWwkWd
aFJQFeiuqk8Cfvj8nRvr5qgpi3U11H9Q4QJ/c4fc0AD9e4aaKdtCDOO0YJ8CBKzH
xmhvoQL4ir+/hHplbb4fbxHeCLt0FrbSf683zowMGbXygdDt6Ey/u4e55XKzTgnV
tcvwyJgFsJlIGVA/de7PazwD8B/2fiBYkBQK+8CHBuVfQZvg8o0pvRt1ZyIbXRLt
KiXn0hCvXQyBinS9rWQC39uA6CELj1O4kd98/y6/sOoTXl7X2cdxTJ71hHTZzer+
RT9ZOR9h4U2FviTfNZv5iFt99SkkZ8GEhI6y214DOB5f2LRq7xe4NTdRWhiavLYv
HCONNaIB+nkKwIwBGJBphq99cKGWDpk+9sp4qznMNHLBmsFbCbRRpkAD5e3qwO4z
oghRwR8ZV6ORc/Vi03sCVWIKRZdSWsalvq0JNzktS3YCmqoV5ony1lTUtm9sSw+P
RF9JzgoCtdtmULRJkSm4nFroXKOx+M/PBduPeo9Drosc090tdFquSg8o8Q56hp9L
BL+6ZErXmuPhte89lqvEPSovwDbM9HFlQZzsZO2KwLVU3Q/nU+STkmfxnRsJL2os
kBFFICejTahzp/JQV5g2fCZwsdvPEsUSPJGvJjcQR3Vt9i+DTzYg3ZAVZnLi4uqq
FrjMy+CVJ0JZ68gZiyUVGh+PCIlBDg3Q5BP1Zxe9bzZYJDbCEaEp6ZR+mzvEYRcD
Yqf71g3kQQ6co1VbHOrGjZYg6KVpLewdx/0AC74UPeoQ9OuKZD9q7RlR12hVgYaq
wrFmq/85sIBOalw1GF0AZyyGxKFrc7BFpZpQjYncl+c0DiGd6dOn2P2QnYnDIwmX
wl8DJlYAU7nNe+aKcp82qqEISm/Y7dgwto6lEGybwCvtaKfimItHrZSXx1Yd4xY5
duLzzrd01h8VyB7ifmGL+5DJXTQJRxe85AsF84dEdpHUXAH5enQkF04S650hJeKQ
Vn8j5PtxYxT+DHfpMKShXPlSjYOn4h/gRPvByqSre81KMj7bITjB7Yg3AxKqxV7w
xhaykLBfAa/hXJnZPQPYWwT4aIj1NAvQzJB4ejLDTnNYLf269cWzqA+kG8ytU7f+
XoV0gJpHBC7MKQNXp26Vpl6Xj3r5SRcVspXOUrGiwwM1cR/F9+u88P0FC398YEVp
SA3C2k02j2CcpsMb92+zjpQed4Kea9+uyo7oU45d1iF0meLMgMT4c1CQYvEVRNO6
15IKkyO+zzZXiEiG840G4wZmcpo/mPHmcVMhokYpFkYMom7dOBzgafRYrX5ao6UA
Hqv2nKYN4R5HYkq7HSSEJxaHOmDb9sVpx6nQwlKkoNeNHrOVPs4DxTWwq18eC5tk
6oo3HVla3mZM3Eab/kGP5RRTcbDptmfBkLrBeQyg2dOfCcVWKJ2Z7PT+9BBpIMxA
9yCcj2bgNyhtJvNyF29vw76pSPohVeCGzC0mqwGkMiSMOlvTb6HxJRpziuIHRicE
mm5HyC2/T7rCMoSCxxr92hqgA8xisrg2SDc7/xSyT6J4aUfP/7gLsl41/AneqzrQ
su+7Nmzbr76wZx8SQntTuFPFy/o7cStIxVQyl2ET5QOpD8pM2XTFCiunlilvAbd+
SDESJEJjYlvj1pnh1snDTHr0XEog4nNQU1jINwNF55NbYsBso4LP8GDZnd99s80F
qrsvYV88HHr+JeOsEZ9R1bOHBUtx1BbjiswVF3S133adVSOBS4Gh05j/L7LZknFE
E2K7NWticrhtREC8fZwk8BT5sgPPXrixmVWLVxlZUZ08heQgyttGTFgJkIuGBazR
pUPCfZrG+xVFJzTg7vFAugZxGnk5xGH5EpTUz3J7vAt3FXiM59dDzDv7Gh7YVqqW
tJi+lBwt5L60UiMRmracUko2DwnCaUyyXlSl6c43zGJmCs263iliPFlZVmqUQBWX
mFRgzzuAap9Ct9+tkBV/QYmRVeIPrnI4InUZDqaMEI+IynpIhkAhQGTm/sokNJBa
jc+jOdq+6eOYdDhaM5/6/CBn+2BVOF/7RyILj4rFFgR9WpGmpfpblzqtGGve4Oh6
bCvDPj1BtrARtjGiZln5y/BLuKtidDlTQniZrVQ4ys51GsejeRZ6tS2hFvrVcEQf
MSE9EG/Lo/tDUd2v47jwe1dnQnW8Cfxmsn3WznKl5YmqUYrXfqOYOMyyOe6LBHm7
wM5RIfcYw4O9+jnGc8ICPCfUczu2+Yk5b7n4oMaS3fhMHw0n0MwCzS0FwgMt3W2T
+E8BlN/ydMM+lw3/n9UJpy7MNX8tmB7KQWYwDBN7uWiAOHTuE/a5OfV1tjSxPN/v
4yiuNEHwTiyq3QsH2Xk32EayHQtIoo0SwvD5gOLxOnVotnjas1WX8k2CTVfJFCBx
seZvEP1li+qfDPvoPk1WAILBRSBJmL5NrAxfDP548fSdXVVZNNA6xMDnZfHm+S0w
QSZqfyPoUk1vOj53oBPORv22yGhNKEIRyKDK1fZP+9QISc6bKunIIk6OZgb+ylE7
GbOGNkZxoxlbw0/MMAUG5J1lOv4J919bRsuVJLtbJwnOzHA4sUW2yLjOhZoMiBmZ
QdMQOm8RHLYD48pQ5kHdKme+JGMF0EPSKdhX/seSRGS8ZareUPSXIzakh/fXd7FW
SHDtr9edMBN0bZdsDY5vUSvHbVNRJpb46GAV4dUpS37p67dXlEmXiO1829cxmiSK
9Szj4yb6E+y9gFp2E6uFeRTB6aRlBQHNYC150H7YHHzPK1Bb37erljQDAAIhrSYs
wqlezu/oKg46LEroGEAnRWceDT9/3QepPeqO3Ir+8voLteQu23j9P622+bbPH67k
s0FDTHSpYEHupA6SGccnqrjr3FRwgGco0d6FWi1T9h6FWPCsjW37dNNfrfwonCDb
feC9JVIn9aqwnRGYsN6N/snhGowJ5oBcFuXkzsfDQtIEfff5961eUyE/bZL9fygq
/1/UYJq2ssQU9QXdrKzoG9BO5NuYVWuHi/C+YL1QpQl+pXKylgEWhPnzN+LqSa11
UymFlwYcZ+wiSYtllDAuLmrZEhZDO8QfxYwqi9X3t4ezD+8MTf5CD8UQaympvhwk
NXvzojj7tj4TtJMf/+uHxie5jLXJ/LC4P408rIKXelpsUCwfm5lWT3+szYqz1qGf
4+DVvjFApzpK95sYoskl0HEG3dbqlYQTNfo1xsfcfU3UHdVR4Vl866Z1ZSkMfFH6
XcGZEyzL7mipmMzOLJKicZEa6U1pHLl2BCzN1tnQol9QxeOs6Rta/fDWAsU2JrIx
L6i0cIR/OFIbBjnlENBXqLOjaEUrQM7xMOI1ED9DXryo00x9kxhS+6ytwOw+KYGu
lmMyBhhxBl1RArkoh1kPR+wR+CmYaC+StI05kdRujmBU3ukOHo2xU1IxDqg6PEhl
Bwtr5XC+JxxD22xlL3VcP82qv3rFORTgVKqK6CLeUe1EuYXtMkGbCs5q71LGVmay
54uLKLeco5Ppu1kcHgjnljf0w42+NaJwEKiRU+ztisyIf9RhDI+yRn5QYbcApTQ2
fYHQOwcoa1E1phPEYegfgrgPXjaYBd3BMxEqQsmNW2dZYgKDRCVIgykGk/WzQtge
4ZJc6rhCXpAx7vMpPxwJ8MEph4V5nvu8hWlLUyCpfi8feGWltVb9c2Ddfjct+K8y
+4QMGMoTqyq6wKb+unRsHCjMkC6WI08Lm7AXcxCM6YACZzNwGFrzgC9TpEFvyQxm
9+jAlOqbcBeFwSpcrgFjclTugtNE6zVT47erQg496tbSF++C8LDKDVX5FvfRbuXl
etpkGzK51+bPonvI6JJdLlAAnq/Mw6Jxp+dfH9dXAqpFPyHBfA5s2a9biAZeO3gN
nulvTJ/4NpxV69A6T2I9snuIRYtzh8NGNDPS382CIFrDTUBH0PzzdlAK4fZ3aZGk
J2PmXzFT0/LpN1/IyVSYsBL2m0ycIxmLyqPTXfd8r7Pp3CspsndrYzlYzQ1TT7nh
7IqPlFKojndreyxIgGUSgWFYK7wgmsmjUUIs6yislNR2Dxs9wBCpiSV2GK/jkdlx
sguni/CIARPi+7GWY07dUCcUucp7Nz4Eqd0Y3Q63uzP/71XkyRr13VBsxdi3668Z
rbE9StaMhi3QWtdFh8+Nq7NyKXNLB9mCLR3zTUmgYn/iSVErfm0wZOb6NpvPVz/O
plInuLkLEiZNBWpmGc3T8No1ksumgwmYt42zsDyA7pETPkiKYOBoEb7GRceQj/K2
hbq6IFUJEhiJdAwxJoxW3GM7mJQTqtQxaFc9zjGyvg7byxFUSSFxpC+rz5yd7bos
FFM0OJSJORfGg7TS/2Ch9K/ugRW+Nbkj5su78NREOtrQioIv6IRqlQHeFwd5mkpz
bykn9RSmZtTcGdDAdxJMV8tcd7S6e8DMi60288HFL/S7VTeV42Nx6HwrGbEYu9yU
FUoL/HtctgGyiTex7zwBG+cpfED43+iobWiSZwmTOXuHUhVYTNFQfOcJFQd3bocC
pGn4+xCeUy2Rtk3OgiodVLvsdjbgiamuEzb1Jb1AI4Zu84Al5Q/8djB+tIH/AwT7
aJMS0w2SOHOR35sXMLWnD4artxPE+OZEzpmZ2tkh4oku/RBNLGmR6pJ4rIddA/Qn
0l28++TQJmSkzW7rpsVo8jeF2TuHQatZh3uRO83o2Ov3DrxKp5EuQ1rISus6t/N+
Ly5B/6AgOoGIxrs0cavtSRXEO94ma0gPSNHlZUHDEeJ24iOBGovB/BVCrC2fC8k5
M9eHRaHvv8WmakMsi9D7GMHyz45Mg05ozCv3zgySq5+wd5j+vH23NVToTqRVJiyz
86xKW3gpbGz0ZcsTEmDsyYVhFbeuxYJ/gi+2n74VrVN0IEE6WR7UCQ+5kFrSFK0P
RPMnyIug5iDsBIcJCWsJpoXHPoiSZoocXCpV4T0/FI208XmY/wjvM0Repc6Eyoju
RIg4Ost1jeEmwLgBQFZxI9JzTfD/dog1hLlZAQP9Es5gtgepWMZ7WezaixJ4iMTS
VqNDpGOSCVxipInCWSQSYZs+djeu/SHkeGSR/NF/WujueIy6V4GizBOINbo5BxgP
KWUYiCAf4ZSNe7rauFeP2fjZoPXYdHdeOBo6fJEa7DK9hRjBlgpsswFnXqzR7/M8
hF3uhh/NUXQFRq5oEicxtkGiz/YricJFX/DLr9Z4+timpK/EWU5cwKGbwebAtm2t
DpfEuRT74nzpPISik25/MQhhckWpd+u3TDarl88Z0WFY/rIgq9P1BEcePsq97XJ4
KByS5c1a774Hy6r5VVMlNrvihSjYtjpMgOQD4jfjbs9hVejfBiW06mSwumCUmck+
XAmVk0oCHY0uHedhktDIkSKk1uUT3kWRJjliedXNILSgWrfkoCfyaDEyKGy+8tTq
Dh6p5rfAuMjaXgpysQVU1EaYZ6Apev1jT8fD9R+6gLaBzb5oOVH9Nr7PepDwbkfJ
5FRS951M+7j4GeudkNpzawDYyUOV77mzT4L1emUIeu7/TSxKltyYYf4u7iKBlWI2
rUdgwvXS8tIMCeNwG67JM0lRBIS25i2cjG5gA+W3utteVbSEOpkAdRkoj7av+OqX
u4IfcBeCRuSMrtr8idBfsdU/c49EhbpuS6M4x5RlfdjhOaQWp+uN0NEqOoYKsK5x
OofVKp8dy0N0IGssfxW4m5HeK7uWpG5SH8V7RL6cBgrXimDZ0539gohbzJSqkZpz
WQFxprh8vRYKr+yPemHgtUp9tGPsyKDPNFE9UnY1bxdCuq+PxdiiGa+lu4KRCVcp
mFp6t5oq28pRwoN/1ax4ubmApX/OweJpvcv70wrzgOcSUt9OdBBXy8CM6EY84k3m
6SbAKuP8iICKT65Qf8Okc8qg62HgiwVSV2PRb5+WdJSpv/OIMtEWNOBvI4AVurpG
cHuCi4pGEbe0HNwg4H3VQfoH77fn2sULAFt6Qlx3zQNpJr2IFFDyECEXjgzs9kcK
XsLGZ8/3IHPgSZpqQoFr4m0CK5yREBs6VLblH7IBC+r2VHcErdClOcNqbu/9xF1f
FwQ7QkKr4PAASTFOICG8t2vmCw3U8dGpFZGjDvnxVHNoH/wzhly4U+FXIwIj/cZ2
afIC8LZn/FROjf48ZRm+ktcoL3qVFGtZLI3N8Pko0DgOQq8/+4Ws67dwqNNGHmg+
TqHcEjzWyaaXSLSN3EvxXnnIJrE5h93ChjB4XmyAHjlYsJQUBWWSUrxXp9Pa5qJU
cXWx9cwyMFyIk6UfusuoPC15RIwSH8LqdPV0sgq5mMcqOXe9ZYEoJzPRKeX9/4vG
mDq1vh4A2rGqVVKZemIQF1g11Lj4gz016tC+p3lcgo6Hhqn638ihTYnolW9aFF5b
LXeXND+7Ujx3u35I+4Gv7KxxRSa4Z/ekUv5whTYOUIgXEXHGKM5+eTQTO7QwjhFi
7ECJtI1dxkt/1J5fjXdEvwlqUlx39ipm9XXXgVE53BQrtMGOaK/KoRpjOZ6Eee1c
rZoqo97kJm9L6r6tGsXvsHFlsvDXh++FPrf9nZVx8ulYk8ia0zeAUM7lKi7V3jtW
KS5SaiKjyUCT03VZ8SDRi/yrXiLqzKGglrE96IGEhCMrvI2qjghl3ZcsGXeQGiyE
n3aMZXxCdDwbim+rmnn8j2DczkWTKBE+05J2JYOqQEanz0+sH4b8PQDOmK/ZXVgh
Qi0Us0vBUA9CFWXOMUXumXQnEhpvIh4vGyQ6Tti0coLRR3CPNIMPhl/RA+7mpmdH
arw/T1gwBweyB/J8T5OkzwZVt855vIqXdbVZQREHqq9eKZkK/mrlr5afc0B4nTkz
MyRiKtKh/s4XUWAWDusd6mu9Zxoe+AcP1F4fmfDV1KqLvBB3+Gy5pVcSgQmEJgoO
WX9rXNAax6rpXusKWH0jBtLL1XlBn6JlNNQem8/bx3Ed+U5m5z/LWJ7MPIGiytuT
5LkFm0UwdCvX8D3JkRcbijFfou0XCFdmNaiApyEmh22Va1rInNo4jSyyXzFC3gCf
5wZ+UIOUggRHr47tD901Yno0+iZX1Wlwz4mkXuZxtXq2L0WJPeez8z4SlkjfOLQp
KutrhvICuWHH+a8WvE34sq5iezEJarR0gzCQNNJbnOYuB0Nns0T5sBDxsNE2K9Ul
7BOAX0SJVzU/OZ2XCeEYSE46dP6ws0g8I/dp0sEyqu21iiK9/JvxZLK8B9WOfi8P
cHq8eKTKbPC3nIhOuq4amNCwDpa2d4Efqh37Xbqmh0vOKvqHsNqSbNQS38uArIaZ
qBpo45MAkq+ac4ESJZJxzI6RRHw/ooDraJIP/hIojkxgf34s+RkZKoEPiJgJhSu+
0F1gAeWBNvPm3GuZfjCRA4lO4qzq7fJvb+U1IpoyQ4buZ25IGclKBOBz6gVwbsEU
sgrygZhcvHR0XkbY58H3B+pja987FyN7LjV0aA9Ysc576KV3F1hdedprQomeVJD1
iRMGsu1a4lR+koChFBfilidF5u6FIdg1XC+er9H/SWuVk4AbP482x7CDNgcrpSHB
MrNez6jSp5bqMO54qaPiW5zizTykWRdocOBt1LPZRU1tXXoXKcnGN64MwZ960qKb
CLdXWklFIKwOaYAekNb/q3QZVibakTdv1TQnimrl2UG/5fToqpNvN2+d4RNfR37o
VBFKNuVnqoG18xAfQ84KClfuevE6KjGmlUwI95saIJxfPEOyegTOWSeCy553uUu7
NCUI+XqBMmsEtVZzJ4Lh0g8gDyZfm28IPZxSGks8vssNjCN4eSH0efwA3HiQZqe5
mOVN7bUlhQ1b4fkV5A476y355vjTW5xATzCW4fFAiyEq85dhj/SBmtBFPMoOxcxE
MarfhUJrE9+lpr9vaY3YhOtpYrjWYIxXn5EdX+Axy6p9/KEG7bbNurC0pzn1oMmO
wSqMbUyQiyDWCFgPw9k1Ib1oJEiilDryUvkYHsX2fsvbLwybSgtuJfoG0Zx05LLl
tn7RBiZftj+WOjFMV484vbGDxdQD6YZlapSRLrflY6HuECLxDbJg6Qvq8/8CJep/
6JbnH6pzWcMgvNDaLZLB4y4NP09THKDrFP5TAhC8n6j7fbOUxwMkoydp8LobtSK/
uGPl+zLSesT/u6K1hG2ABc1UY3Hrrn0KFCJeOfeMyfxOsADQYwB52WHz7ZXSMHbr
TV55RL+SizIRfUOqZULINurpdiCoXJmOSyRGLLrqLElt3TF8HZYsp8sWxTs2ya6J
SNn9I/fSlD3oOP46cM6yaRsweOjUf6pldMd/64z+OIpnAdR5DTiSNIZIM/CG4+pi
zWqD3aTcgxUL8N0b50ll7fc3dLVqYAonSFX2WN5MLSDVG3jDB38Y2yASHAUIIyaG
3ASSPTaU2bXHMPh8O6tsBfFe0+vihv5XkC+tpU3Vq203gXXiZb4z8e+cJ6dwF1h+
e3uE8F5r86E1BjiO2fbZ70STpar1MDjXNFp8BfqG+qy2Yfc49MnYoeXjyJV2QcIL
6whzIQka+dVSWnxPgl02noDK0k1sXC5xCIgwssutl6+6HOQDsfYfhy+yrvE2m2Q7
Yo0c64X6ZFIOzk48Of21pbaTATe/ynJWg+uMaCVzJlAKt0us+AH+f7xkK3HIRLKX
B9FlC8ZhLRo1u/dkQUCCu6FegaHwtZq5g9V5GiOiEA3GiQ5vbX5h4bEvpVkTZnLm
4YIp1NKoOJOwtFcsC1a6Ifq/8uyoe8Xrk8/QXnTB69u5hQa9KSOlAX2DPYsIyo3B
A7RlgaEw6hzCKIX/KJHaGat8ghorJ3LynEyM2ZzMiPjFzQt2KMjoLR8dpay6NuYR
mIWgBNihwZXnu38t7NEY0lr21xY/Fn9HReYlAqRqORPzec5tgPr9ItmCDdbM23KG
ws0zgR1rskDdLdZBrExcEVtAnyqwFHOOy9PdP1Xy+6Ri7qiwctQul+JQfhsPygbf
wNgLtT9lEck+c3rTRcnNCQGcCtUDOUxnv+jjb3mOkRgRcky7G+0/3he7WmchpSe6
B3wy1Az7KLFwVNNaOrIY1TYTo/NV7TvD16hm0riyU8Cs7yljaEm3beuNUSjdFRFF
UjICFZ/lEy8ybXBtJkCHzmeml6Wwdbr67vjnONcCJUNEHpg7RKoIWbC99Tpx9r6Q
tE7AZQAxFLZBGKIqedHfgj8K99Bv95yWsSY3cPgJ2YjxMVtgUKddQDt/vWYNRqxD
ssotShDcDc8wYKKbaCPy1DP5piVqXX8jvxUfLSoj1l2CH6g8TdYw+mCfJal/WsGr
SizauTZFxHKsK1BkqKqY13V0vwVuaf8tzgC8o3NOkCFUy48SFIRA9EBXUdL9rkEL
HmZQ2APCPEVWXB35/Z13fyPMOotVHOM3uiXMqIha+2rk0FRv1j6WV6YDmGH/Joyu
rYYTU1q7p4OLr4Yxbz2aK8A/0aGnHzhLiry2E+b3qNuAga8eOLEkIgd4guhd0Kjr
nVMVMVarA82ihzgA1tGY49EEO/4yJP9E6HxVcDW/o3eLf5PcPX13zVvlRmj561zB
ACL6giEPn5Qrd4napjXm1GLFpysofwV/K7rKqJ7ezwmSapb8C9URKxc2zkuCdshe
OfdQJRkDccx+cQ/HOmKjUYwXDZWPhjtmYaz8DpdgJWk1BptnF+jRkZKh1X4h/XkC
m1+9fEY2lDihzxaIstjiWoEhKLOZqYWLgVIMS4ZqQhM6lQKZRztJUkeFzP32h1Be
gnZSYd3rAW4sfkGG7vDb/FY57a0uS2dGBhfscqXo95dK+OX/zoC9ntPNz79b3YIy
YuDC4csJqhE7D298cT18/ovObMDl4rDwCz5aVrh+7yKJd5z/CPsZtR011b2+Slnt
cITf4/AWW95Q55mFInDwnKuB0VfepsLj9f7Nw+YkFB4SRnZYDxJ/BnkT9Ki2lly/
E7cxBUfnVZXtoPuTmtMCsi2IK8c8KkDXVg+p/4CWKDwERteLbmJez6EUeqzssH1J
ASUycMGSDcU8tWJzYiHZzjWLjbfp3CfFoEiTj2/FtvmOXuXgpvNi61iJLz0QHjUl
EVn82NoJ5kEtesDqe4BlzJKfbj5faR9qtx6nWAegtICf/VtSbqZgELJyiWqRvDRm
LUh6iExx4Una+z3ZthiRrKAfK88bvyaDS0rHwSFer8ahaTZc4ETDzDQMTF3boiEI
Lle3OWN8P3yQF28rlicNwIOY4SexNp7XSkG8OKjounDrWG5DkHpotbVml5xbuwSw
4U8HTFGnD+ZMPHWjxSLD492paBwU216mNUwhgsgcck2nVYL2qsLccuTrUjIkWD7x
SSsLk20kGxz7x5++28FAx0cJTF/NDxO2B4eSMEMZ53jFcbzPurZa4BMb8nVHjpk6
NrAYHKq78xynG/RealXur80fndqzYVRpWT+y/I3cDbGN1Alik7/vJ+oNTlGCsgBr
dFqrajqv42wvcQ9tYIarb+rR4KUknQsN020rur70Ns4G/rUzpduZ/mF1pjQaOJqp
vO9nOj2NHN9s0qmWpjPJmKK7YZfYPTQxbmqpHxz5muMRarBgC+qyMF6JOhwWh1BR
VpeStSn2F7lKfMXwKkedysUei/jYi3pvdkacv27wsHrK0VjGDlSBP+U7hxDq50XE
ETeQ2hMYhnk+KaHkYFkPE1/V1Ti9D9M7cl8mLKCm0EcEtZkNiz4ZPP/PFO9IOfWG
+Ww2wjY7NdFqmexcuna7c0XFrrO0hZeK7TUSmS8FRGCglCfNqjf6DTGd3kBxzgHT
2H3r67eUftPIme1hW2GpRDLCfo/aITV0f02wvuJq1A8tt/0N3cGJh8l1ejxEhwYn
P0475nn/3PFRV0SDlFOwzCh231dIUbjbuUmqYKOxi/Pow1DyiIsQcC9zTxCHQjPC
NZw00T/WlVUofnGREHBqHt6MZ4AxZ03At13zTKibQxXYQGlVYigi4QCLDdgsArag
M/WWL8HmBnmgQV6A8C6IM7T3SxxhI8Xxw2InXcW93Kelh5OJpwk3SU+zs/b0xrIe
P9MB6JEWxT0DQ9d09GJ9t9TKGKYo2NInOjdk7lF0VsvwugibM9AlgHw3216jRuXe
MDXtfloxX5kTky5TbFWfM63zKcdlpAl2gGxfoJdh9ZsuNPk8S9/ueFXvBjcLkOTX
G6ztb/gROv15hVN8CuwONQnFUZe2gGRH07OoOg2Hw7ybmxSMUZb3NeUiLiKnoeEM
fceA+q+72KtAccFLlxikksja9Nk7+c3wvjjfNQOvPi6qackfEdZbzU4mvUN02HXo
IoyRPROvYbZHnxoegVwMihRs0BuKxo31FDDHsZzJfCt3pktpeVpkVPZPCVRCpliP
C+DceYkknh5X4nho8NDyXPBGBQqV2o7z1eyonU+38ToGRzEDcJkVUXpl+GCv8/Y0
N/NsK8LyfwrYyL4xX8Wq55a+JuYmDe93ZSKeVhVt3INXwYQZHAA/J5ZWd4lewx4v
oGK3eF9OUu2y3J4IIClmhedHs26KEI8RHUaB0SFbDCzp+Zgpffck6HZz7F1neH40
0IxmorI6oVtEifVfSylnN+v6OeHrRZysdTjp84NcXEJWjacQuAOGeY9XaeVe9vmM
R6uFF21CeBcybeMqYmPT28NJJhcyxu2/rym4wxyps56rfEysJdjRjreEVZwp4Xjq
JH4mFPgJ0yCmaunLl+//cEpjz77SNyX6LGfpKVeOuc48tFNS6h1x6sS0DieJh0DG
3ioGuIFofs9lCZKd84lhVENe2nYr905yBaie8wpiI+7wKX81O2ce/FK5DDvOgo10
9xQLNeat8Y82PpL4yjuey/jN+sXHp/69jNGKXP+lRtj6Uu3gazIULj56ofshj2aX
DwJQlbaWud0ctGFJGsX4PVfcfEBz9XomfNy6+aHPjUs8/UI+zrgNSQN+B8wPn41v
J8kIGhL8OUuPad4+BfbOfxHz+WImHcLVus1AeSu5EV5Y/klF6+SberAMLC1jVi9D
g7VEom2oOpwYT9isl3tR9atEvSVUe1r92h+5nElfhJ1sheyAv3mTN7iYy/X8Th82
N6ydVPfqhr4mFM0ovp9xLkTXy0RD73rk2ErUAUMEcVmmRbdpF5IXhexrVON9O9FU
TnAiP6Uq7n3dR92xAjuaDimWQ36jtDMTPU5IQ0wPAoBfurbNUf0Xo2cX0ltVfW+v
MlXlo3rBgJBq2oUOid9jR1B7csG8bHFXIslPOhsUMgdwJ8Bx9QzOc5yu9JXTsa5/
iJlFsQkWvjWjNmf9nZYr4WbzlZpUbsRQa+cij6Zux5e2prxywB9XaKXzFf3EbpvQ
60Ka5/88/klVevriP6vP8Bi2bS7nucYRhkprmGWwK2aQeoYZA2rChLb4ibreP3Ex
a9VaRKVcr4JwEODlLgSoASztdVQXW2UQflugc9N3u9m7iMHJ5Wo++CHzhH354dz/
I/BuK7yzr5qo8T68M7Pig6YjOlAXDevY/iGmu00o3VDPFvZaOhr6PV9tHpj3Gqvq
Za5EauzVgMngcCpaICU2QzeLSZ3hSynqUChjn5kt0mrRgmIgIC/B++uDilJ+ayU9
lyLBS5iV2/9GaGjFqksBii+mYY4J67Qey4o9QfMJKqJuEvT2kXQGqGzK+oYzSXA+
JhqfFRkAHIr7WGPT9ZR1alDHALjKeNwq2EYWjhCfJFQeeCGb9Q2DJ5D4vsrJotdk
DoWD6TlFRAAPR4RkHv9COgH1K5P+IAam7SWroBciqg45n+R+G7rcWCpZao2tcJS9
wqk6DaWKrp+IyOByEgTtRPOGZXabeS1pD4xkIYMcURMWRjPrb7CKRUtnZhGQ3F80
qOSDlPBz9SkTBOMyiq0+Mv3bWPVhvX+XObF3Aos+UlHrOduGuYu5nXMvoF5Ver4n
McQcsNU635koALABTjhLbvmvWvY358rE3YRkKQfe8vx6vSJjBuxe47K8RlTvypnf
2uUpJZIl0yaMW5ZvSh2w1MHToQl7RhTRzrX/Rg7rgWr/g1yWZsOJHKMYIRqWhDe6
nEXg19PrdmgB8R72Of0YI76iBZEI28LTudhyYyKD5+uDjmux+AUWtcJIEOFcCxo7
xwNem7nZLRIkO5KUy2zRIqBVUfChLMn/iBoRFAZ2oKqsreLlwDdqEAWa1RoobY/A
F1iw0cRhmL5yy3uPzgZj1WRzBK/tHCTTMbqTDA+QL28JKRmE04EWhdeIciwGGfW1
qqZs7oE4O/6/GBE7LXrh93Mm7GsXPhHummdLfJ/NkYIcs4ftAt3rIfYpktqhwLvE
SyUS19zshu4ASEAf/mpStdOTfE91It1mzsmqp+78DoKs9LoQR9TpThQgtcW5WJrn
6RFswNmX71A0RSUn/lFH2fX3344KxeEtNFeebvBrgS0n3v+EpLEfVzl72mKZpCku
YFlPu3Yxvkt5MDFhrfqjoeaodf8UIIsech8vDu8AznNGKes4KJLTGaM5UL9b7fnz
hxgM/vLIu6PwTIfkj3DWoeH3TUomG0xZkMrWWf65Lo+V1XtCYHyYLf3ycLoDbhaD
uJXtaGXnoiCyF8r3L+WBD90N/LINpNT7W97ylzD3EHPpQTcJLbzHuVPJXYTHWKyG
2etbsBvtuPb7EhdlFPozVqGX86tZXd8vhm+SdAb+Qv203JIhrCN3+9CmTtyzuPZI
13uNZh520Th/mE6CMqmaVpVvmU1RclLA2mio4dy7MgABYrTAiSNxNVe0UC9aDGm1
veANM8J/vZuibtxMBHbo3bnh1TNmRGBGqe087jZhLoXf/Z2xhTdgHmGNH3Skekwr
xgW2R2jVbXCzeGfthpurnzbJUGJDnGmstWs/XfuE/zozulZVXN+hi5UdumAqP6PL
5R3eCfDKZGPk1vVfndI4bBSyJ9Ci5LDCuAt/AbVMPLw6IRCTrqJJnjp/jO0pPe5w
L3XyF3RyJKJjBY5HWOVFtKss5ktpVHMBRzh1Op5CaQrn8cSWpGBdFbrJ1fyMDWYm
XD4SG2Mair5IBbN0CDXOMoSI9RohkL6vyHKt/Qu0zYbuni+yGCrRgexvU910RDDw
ts3VFSVKx7lYef3RsDRIAGNdNm2qNkRpaD1aOEWH5q7WHgGpQZALLYCz1Mha4zTG
hiDIEYfIxJBwa3HKzcIOKTxvxoMXGDNi6FeMJhVnDsvEqP66HEyDdQh2tor9fnvL
zpK4lAgJGpAfDm/hbLzoslPQpSZXBWCGQRY/XE7M76zllKhZX7fzR5NNoIByRIqG
KH8dZBQ/pRR7W9WNZOnepjbQaaPN9C/0UZxKgcCW2S1AfuIbb0G0vvC4V+NwuJZF
L49K4mEVTvx/2woyYlOZ8xHJN68eTcEXCDlSfqgwbfQn21bNppodPCMxGF10ySi3
SE8Pyf15tNKkK7vtU7rc0J3fPDl8oDkbygWyrmzsu+OS5yvKyw8ybr9cQ8BoQGYs
sDiWRZ/h28ZN9DZunuiu6iGq/hgfEfBXYjbFr8Dn7IGMT6p6a8hkQCSdzEg40TxP
/oJqUqwr4++Rtw8clory5AbAbAxdvq3nbvFBQ49n3QgdBZAIxpGa2roh5A/6YayD
p1bL3W2xpPLLnXO8ExxUFoni8rsKsNz+i6xqhCQxfU0CxyQW747qMjeljzokrZa8
xnvhkxoS0wcYtT56fR+xSlY1XY7YPaNuLR2BgEsrCD9WVBWIoduzzcUbY0tJGLi6
XgciiLRsBe7EK6HL+2rd3c3pfNNE77KbHErPB/9QuKk87E/90jib2Bpn6B/ba30f
DgPTQY2dDkjdz4MqduhkOE1Qrt/wHcW1yFb5B95K3dVliEzM3tlk6lCbeb6KLH1f
193tntj8qGRjQBeEWqCn7lqhHt2DJmBUvTP1nS2a7eV22ThOTRZlpDD2qduiTxCh
R0XLIWYHdDkUtUUpaoDANgO9etEH1S7b7lgLb4T72vsNZ96M80cO1YaC18CcZ9eD
Z8eWqPQ8PzUzCI5dNOBelfNpqx7JdxnKaJD7O7uUQMfa1trpYaOu0dAtPRbzBARx
oaO/oEvmr6z0xRKy2PGoemzLClalvGDST2dycVjTvUSCz8uH+lIsrVweOMYFGygm
RSGzfDsCVm7oR9HPqhlctZP/EGiRa6oxjHochdCdsfXj3lMytCEGy99pO+laX6t/
ujnafwJw00onaUIskkLdsJaIOx6JxxCyOhJD/V1cPVdaxFDdGPtXThgZCJJul0vi
aQKvbquHVgIDJvcga9kjg+Npf4k0qlZYWkIL0P8dbbQc4bwYOUztpCZlUV5eIkCF
6bY7u3isPJGjnGmW81scPYAB94+fFO5ObSFX5Ef0yam2ivYjquur8p4PGbN8IJZU
qcktzFzsFWqu269tPAixlPzOCcXS+WTBE2QeMEPfWj+qvmgF822Tk5q+Brk+FZAV
N8gEkfqDcK6Y+zhLY9mpxFtAfXRZ+3Rblj6MX4blW70B0xEr6Fkdy9OMu03QwRtx
jxgTKQuRsi0+Dp2KLThKRnrghSVNyKk1KoLa5wQmMnLtlM3Mt0mEXWtaRN9gS9Iv
+1GWTzlD6l0/VKjYU5zUeayGos0aAXUWT3T52IidoOtWEOmZY24DVnqLO9+nqJtm
+FSZjghvaPftjDGvH5A7lGgzA5yq1/joKxqj2UB1dBeSKHiRLDyYisxjQ0or9pxW
l+e/o8b+BoUnu1WrZfWT0YFofMndZnN3IqU35Tp/hmWH8Pm+Vgw0i/dGpUYcVkZl
w2shsabh8RoLLc83gMkZLNidEM9WkjdvD8foOiwg12cR+HHHqIEKYU929cFwquM+
RlasV89ruT9d1j6CB8ICHy+gmZS9BV3Op/JQpckOxq0lsBQ3HC2O8IfObcq+rhK/
tb3BuuDcXdyqG+eQXvbXXYKYYuH8JqAcKF85GtBt1qxeJkHtmnmOLJJwc3PAZLIJ
PaXPBcobEHjaiHw2QEKwfWYmKOFQuuP0vezj1lZyRXb6q89r/d3ov3ngX5DoR0u3
rOnrLmfHKQdrXvvsEjWetzfuuE9ZihQr0XpuHXyGeWWuH9nJ8ndvVWuDwrH7SBgB
NAcnuIBs7NFCAR2b45TEIv32bpgGbiQCT0+piZkx3hyCd9diglsJn4isqaoF80wp
T4v9rx/nhdMEA4sGPMRm+oPxCigb738+pfnmXwXdzXWBIUs+lIWve2kSq/B7M4ez
mzGL8KZ1FrlzRrjFRYcjJj0pu8Oa4Mjt1bpUlxZ9GH8GNWBB5wHjtygctWSqlVTa
PyLbvnkuSwags2XVZa76tYvCfdn2+obOfIaK16UoI6gUypRBCxPjgjK/oLbEyls9
limlonAYqhtWfL78lZ58jVbD/uLRIJiEdEud7JgswX+CN95kxspUHE/ToX4E08tI
ixncMCw2pVYR2Z7ApRElOrrUGVac27yvQQTbnKSduWwM63w3OHkWfwPXw3pM/fB0
VSMhHidIUKXZ+hIJGa2Wn83dItQIofa7taypwG2+bvjmJF/iVIkBn/RO0Wld3D/D
djD8+JJ8nGDoj3gSvRoogedR0Y5ZqhhAhwjglhIqH29A6VnAlygpfo/052ut2Z6b
WY2+0/KTQzOTpPCIcu3sYSUdiz9EXsOI+SwetsUjSyEUIYrv1faPUt4dAV89bAJw
Isk1eo/pN7GyqVt5ZyNmvNVw0LPAZ2yZSFhFyubJbsp7vvzAb2xEJrMnLGEWC2cl
B87lfyHCh5zdOmhGLQeHtY3Y8sBqF/OBbyJev5iXWF42QJvwZqzeVPgXwxzW+Gni
jaw28MPVXsR1u9IW9S2lyaCtowSVHMkdcqD98AuXGYKGDoyjVpHEzX4SGxYQ93Qa
Ka9YQOyafh7WuQ2gMjyDxXACxm+gecbZZEvZtwgwJsW8ZdWvGl3hz3q8z8J8GxS4
nlNSlVAvo9gCJQ+Jb7ZM+K8GM9gCLtt36QPFLokBmZW2Du+Q7T1POcuXgtIBe/zI
6uKUq/9kp7Zfs9SDF75Gx+0/nJoevmFvE+rKHDePBJqgEqRRfOvyV42EkSwttzfY
MJ9Z81h42oBxSpVFppRy1Hxq+d5O5Hvn0Tz7SB9HHkheQrZImpwQ5nw9kqjv42kb
A0O66U2DU04Lg5tm7/ZhN/m/X0GAAAXqJXQNa/6DykE9EmAwfnY+FOz2Ev4USkox
GkkVSL04++LHN3M5KAvHqQQtYySe0mpoSE564/rtJF478xOv6+tx6jZzJLmGVDNL
HDaC2Ffw5qDThs/u9B5XOlY3Jknb4KRq8arUXhPsD6o+MfYJbQOVJuFJ9liCuC8s
85HY1hA9YGRK7/phHjpppVfv8E0WCYt+CalWeMY2TMFqXKiTxkhxoVEs1YpXZED7
9AnqkOTBGedMYDoS8viTw+PDT3WV1Ro4qR01N7teEzlpdW25PRmlZHMhmFIeFXSC
UmwjATg3RN8qFvXnP5FyPfPfLlQRsJQRIFMPVKO/X6qyBg0PDLhxYYEHwxKtByRk
lGrTwA2kvgaAHMB4Y/VWb+xf4kTmJX1fttHsOfyyAM1r/01qQHpYj758Xw2pDc2S
9TA2zQoumLVIxyqvzEaYhwa2vrd/k7eOZVaqmjqWjFeke5+Hz93fCAsvd60dPkIm
LTCyXcPEvL4AY9n8BNJ6WrbNp/XJ0yXfghy18Unb6nGP+rH5HCJ8aNbzxpUnxxQW
ZUyOdR9xtKV+bl9GcB12bqnUF4MVQffT9C3H9AADVF6dIV1o+3Edgla55DNijcmz
Gw9+VSZHwFd/Sbh70mVeqQlQetZJYv5nsGaBgVs7h+R7A3aUpOrIyll7fCch1Hhh
Q6we7L+PHNXQ9XBARFXSkvkBsnGCDkwIsYtMkk3xlLq9nnghxE7yeripzXR8pN9l
dZDQBLVFhjOMBkkKS4RoRzLdp/1hA+3HMtNIex1B0C35wIw1GlSy9IGG/AWGp33K
8FqrTLSgLk7hnVSNvok60DzxJTq4WMdjfYav7z8XdiVKsskNmPSFA+H3P4w/h8QB
DSG4jv0POF0X/KN43xvIWXUE1yyl9KTD/g+Egx5KNVvo423nIjR+Au4sWbf59KcQ
YEA1NHa1UuR3WZ6BQui9cCAkSmX25JuG+8ofEQ8R075dzvzX/Vs2Nz6ih6AEAmA/
l4K7Inz6+CgjjrN9dZQcZZg9IqwhJovvwv3TWhiwpUTuvQ4LWaUyWOcI4GAwDNxC
CmfFeuuo5zJRwFCt2cmK3qA+wHBHV4VuScMwV+mXl0Ct9PxUDSJ8yOec5PVkPO/j
DRDBr68Zi/1SamOJGbt2ME5SmF5wTEA3uNq14bqZ8KzcIFF3ToUIyFo7NjQf0GjV
IIHP5AwrsvJB89AOf2EABAbm1q5IV6770AZpjmZ6esvRtqzXlUt9oKfL6bNpGghc
KDDNzaGX5xH1yyTumitEip0QM15HnIITBvcN4u02j6wfHxu7hJvKl9Wz40kjhRiZ
vO3yIYqtz2ddYZkN6onxFQGNmg3HJiHL8dARx2ckp83ZHwwpYeeKaGRpJxG3G6Ko
Iqr0U4YdqLYJqXsMalFqv9DcboBXt20HMtW9YhQaXYwxh8RZc08Ke+kF7CHQUV+m
ktNVfCBs0CJV5tgR/lkT4Tl+R1eB8Q6m6m3eOGElNUpR6OIWoWC2PPTGUV/J5LTp
YB/EwHKgzf3CGjIT3ctPGDOl1EoGQt+gh/YLHrJ2DTFZE8DYg0PPq7xqRzWMnfHS
SxN9SsapFh2dp00B5KT7UycCZbN8qXJMSHk17l6iz24ZiViDbe/c6Aw/++2diYbz
L0ckkm97fRhutlD007srHZ9nm/b7Q8m5LS6JnNyuNa+y0NbzyLskOsodKQ6XWfbP
IYPynKwibDd9QjTcxZoivU1rTxQpIooBu4Y+zKxzxQRcxiH5uWyfV3LmgkvyYVQt
qdFg/QC0+ctmev0dIfhBCMq7ns1aSNwcrzNPapIYZt4fPfxdTYt+lVhuIJvcILyl
GXxOXiy7EEyGjKnGoIYdznSdWLc7IvMYmnXHQ0d+vPIlMvbyo/1qUoZFD9q6VD5j
3f7e4lr0PrZ2IaBMDPJtulYBittu2oVTSab9lShRF7G16oEudgFadCvwgGbaCuDo
sl0MlTLKEcT9q7+HOvwqYs0TCto+I3m5eu9l3u8eHGToW/A/2d0EB7qzvB/LI35A
iS29tbHq9Z7/KuzwZIbVVZLL3FDVzi5C6cs3mVu5QHMM6KDyHQO4emSkwxh7jd9H
BZVB2f2ZvU94kLropnPQwX8XioGdDZhMUWMNFI21nHxW9tLs9YUS/LGfRGvxGTp+
DqhegiQ8FK11SyctQqtPKQZW1IorBTHxbaE5tS8aYINhN1kLHAScNEfj72QF3qpW
qk1NrsDSLplycHZaVWoLkOd8nNj+sLNWfLl0U96f42xB2qSzsbAUN1a1H7CAZds4
qDkdGg0OU9Yk0BC/FIHWpGPucxROaOn67i1jxrs+0+yPuV61ilgjGrzYjkjHMP+S
66Z9zpcgDapfS0sownfTeEIb9Zcgae66KDl0JEliC67MBMsQpJs+kITrs9Glxg8H
IHEoaeT6Wa1f3DZfVIgy3+FJlIP3JSKF86L8cYABtjZcv7bE4YSU7HTWO0TnOc3e
QaOyUGuNEtQlxU30eziiIFes54U8kdoj821dXY8otDbymKhqr06Yfr3yLiwk/nyf
4asbt6/0PpnKv1ZbqpQTVsFdNPiCH26v4sARelM1RNRxYPfpiFFB5O4DEmB/qWE3
4oZp2Ko4EkLapVyQl6CTGXeWvPhyMkMmhUcaEPOHJSwvQHSvArKZg+w+UE9acTHW
5urRZ08biaNGObvoHFjkBQRDi8hGHkTmxcJH3IsuvuVvmFvLNp6JHbK5H+aqOqez
bxScUfTlJ1GJqagF7PP/2jqeDn24Lykk8dYwNN9xkRdXpjxf4iO62lfSEI8GXdfk
S+DcnJ8gjhpJSSXINkROAztjOdap9GVO+Wb6XRyg89Arienwv5JnDUZjuK4DEsDF
JB5NCOfMsIjmil69h6zKVxT14NbMxIVLCEHZGSHuSLDw37HLznRYzHlDSYTEbZE/
kcc4BZPzwcM8ojyM4/e16je8lpRr3R4Whanoa4Oqx6I4CKqNGOmQNXGHAgf516Hv
AYREvo6Q6ia3tBBiTeFLGpqsA7J5DZgbqVhXdbXYFeOK99Z2I/+5vVCu8GffYj+P
JeWlPOHaAqO8sohBNNSk/DNwvu4gQyEoFCJ59kttTvNve35YmbY7Kyx587yh6V7Q
8ts5XdrlZkPJzjbFAx6mL0FNpAtp/IDg+TG6dtyTS6aPv+LhrtT9ip+4anBqcS8M
/jDg73lwgLrd60hCwnN64QId2T1z3g45EI96sMU2apZj4RA2OAavg2r/okn1x1AC
xit8epV0vlhOusuv1DNSYQ1Dg4SZrWStm6nv9EnONXXhIdpEbbrRgjqOdLjfdKJY
X+fImu8JnTkhbAD4I3GqScAiaChRP9B3BJf9ct6O5KU8J8MKpEY5WEuwr6dGEEX4
4MBhjbV8Se/l2G0VU85rzee+/neVRyl9n2wCg1wBkdF+OSAyOeJW9S7RgEAWYiXu
h3JUCAjmjmFjT3VT5tCKr4UnLZq++tNc2Jww8qKU4f6/ysg/13G7LI6a+ouX4RxN
I+DSX4hKJwAVIfJTMOKfObUO6sxo3dH78Mj2gScVJxyGEEY4/gPaR/jnDA52Cf2A
RmUJk5eF9jnKt34hYm5s8k7+W3apDMZ+w6RUh84whp5gcpAjzMFrc6ejvUlSanFK
vh/9FGvlF9pSuTMIrUcpp7OSDOUIa0Lt4lfWEo8BLCKVphWi/vllvb3ZezuGL5dI
Aj9AkNST6FJtYnKGpUTwk9LMshriKAn9BQyG6KSkrAF8obPOQDhI1sfAtFBvnVci
Pc0HRuAHf1x/hbPcGmbYee4qbM3XriqLyM41VvAbt5AJQiBqma+wKjuAc5+RMS8O
FWgMLXzx+ffKDGtbvqLoLiWl0TMN2jQy3PZzYtJNuEzKTHABsANoJzyxQaphVKhi
ZG4DEi25WvAZDHHmAk1c97rUFtA8KxeN9szw0mqhSzMR8cbYH8fHSWRw3ZLL1IlY
tTQj9CPTcPKVAz2a6rxIzPxb/TUcfx3TCNuIso+vQDHKbYSaEZTjR6s1cBk/6xaZ
lw9VY+66Hn3ZgJ+KeDTtTbSvoJvYY7PWGkR7OmyZlz9FaOWNiFYSNW7AYklvtrMz
pgzFl3R3RuR9xtsJPywRcmDqHJDu3M7/0N7aabtWkUACiAv8yZopKyC5Y12TTyZg
fzxoZkSrGiIAvanYBhrdlNzoylGiGw0G2TosjHTdwYmXdGwUDYWQ6ri6IYOn07ay
EsvVHznrM1YD7FJUnVTpmasnQELPxXXwoihVQzwanR49Ar1zcVc3vD4h4QFLbbFN
mKp476xwvsbzmE/hFT1Ia/rWhPfHrDm4tNrmwAAHQ/7iMdEgzGZUx/38uIsCQV61
2ran9iDL5MtInalkxOryOUFDscycp2RwyjE55DSsh6VZuRXSbupH6X2epZsUnuzy
0Lvxq4YuFOQ6+9AQgt4TPAOx5lJladTpEuN0lDZNKTlXFCUgRK0q0xyDVGBPO44/
dsNufMAR4Jnnhw+8QkmhyVC8dj9/D/KFiv5x82FEl3RkGfkxu+dJpsoob137teq/
sheCHgQSFZpGmtRnuorv5ljmDimHrI4gHlFtm9vmtM2yHDSGc7clTkeTIi84lLtk
a3DkKDk1UplQ6Yd2rhNnsZV+ehNg6SSAlFQJruOCpltclzGoxatdn/pmWlIS70ga
FbBfNxVcDq4JomthZJUIEKWXkED7yb+ootO55uSLKcyBB18iQSr/eR8doD0jmR39
bMs2O06D+WqlxQkskqVlKtPm7lrOt9eQ80ApLhtkAVZrQTJZ9vG8BwBq0+dU4Ylh
UgF0Bgb+5mFVtVlOf5H/S2g2r6e9wO67+YfVvtu3GHyGTiZZNaTchyKqsiOlPckN
20TmQfX3aKWf9H5IM6WU6SKB77OX9dMAC116DxntF4qNbJ5RkY4cg7jZO3+0Cw3w
PhbJmq1KkmELHlOE/6C0fiIFgjEtu8C3VtSCXNN6vYuwfWzHFIfKwCU8Gx8GKVFG
QXCYHrnslqG59F5hhDT85eV4nkU3sUxR3m+q9vP989abnEX1qqhlB2mO2mS+tpYQ
OLUUuO4Qpk8Q3ZOhgoG6p89zaGcR8J1k5IylUMaVdFV3Q94ulEum06TnPWHEpDh/
ulkNO8GpZpQ0hD6WxhTlFjK7deTuun8QlKU+AWO7BF6M5gbNStVgt0hFY1bAZZ7o
6A3I0pBxyW+w40UQXQ4pDxxAD6dI2Mbgf0p+XaP1PAdzjcY3+RKJmg4ecrZjb/u6
af/a3u7rv3eMPVSUgqRCZQb7UBu5A/gPpOrCKx2dGaRXkKEpshAn1J0Rus8X0jFG
mvToNlZZtxk+cgRsv9aMJMUZIVatLkHUG/p4bTOgrZRtOTZjxff1p0bsP8ouyh2B
qySufCF3V/0UAdRKK5Oe/FPQbFldMKzSZb88zKudxHcHF7k/zdMTsocnt2VWfhKx
hCbVwwYHlAOGC7jrJDInGdREnFmgaMoKCOO+RkzGp9FT3r6cBMSbdvZJRBDeCeb7
HgNwEGsbL5dJzJe6esVMzxIXr3fQyVAjlmq+Vt4IdtLDvx3idscAoMtpUAUAHVxo
RGFO45C/IzrW3ZBeA4aZXqlqU4UqNE0Fu42Tfvalc0jQvU25XzQPrIwEeSk/8sS7
7xgtiIqhPi0MyI8+VjDPdzCWGnKWBYf4dYOYhcng1Bi6GJoClRklMCp/rvyYcAu9
Q2egrl+HhT3GX9QOf5o82ai+qylzPUCaMsbPY+3vO36ZT2RNSLAGYzxEcfO+kicc
A/R8pg2ymsTIUMoZjOcA0SvECOSO5peRqKLP7gKAmQyUFBnC2IdWU9Eo49/lu3Rg
gXh19V6nubX7AQ4HYBkZjbHRZ6Et7r7QOaAtAH/gyCs/DNKaZ2UZk+af292rZoaK
MuvbQjEvzyyW0CKSFZgWeunwl8NO+oEdljpbXLLLDSn/h2KHwV9EyRX/F6ZBwSt0
jrU42aD3x8RT5LZTGkVO+Vo2QGFBI06hS/1c2os7kLffuTnWM8ATTt+TD4LNGcJI
P+rh65ceERiGbSuoztl/+oMLHRdMTT5hCBZuH0z2Sv+6Ee359RKc4WzAOmBqXs0e
qtCJO/guyfXxctbJgwZ4DzI2D4eNntCqqL3PFgQKBzDCi+STHZizLqvPak6cjBWS
U4D6KcQpkxiW4LpAwoEQA13CV4xvnXWqA716eqbHbPEPCEN72OuHvVl/baqBgSYo
kETdpQbEQkF3BDznFyA7IQo93aPIDlfOJtY4Q2d+lfWV68ojGdaVN0B4hA41K6a2
MeU8VSoTAoxYZC6NDVjvB/2w7J6gn5Mm5aVlxgkxgZ9fnfdXpuLmcTQ0fin/gRmj
0yF9y7OxAScfjgFJORvKw/PLECJceo1AJrom7HfIoJUiteWjFkTFQpJxKx36a17+
AQ/i1NINVQn8d15YRzCT8EEXK9LoPTWEx6+OBcRfQlraIwsoFUekVJRJSF/ECjEu
aa0E9wwbZVwPv+npAJkLvMxt7eqcxR8A47R98fgeqxQyTsVbTL+33tc0NOX9m63U
wRsUUjpblsbm7dp1FH2ZJSIv5wHbDYJsaRqkdqeTlqOxmRrZ2Nuykq5iHnBqmZva
dii+3o11wFCgRx7ujc5vuw6AaiUhCoHLdsgrMjR9fYBiGPXKTLaY8Qf8iGKs6Ekb
c6ykrjEDO718wQprY9kchk6wHq9JR4NcmWpsdDn3o0q/lb4nqd1FXVtewPVRDHzK
ftpfm8sHPu24bhBCqRRUdQQ3og6m4K+mw/rWqaSOfmi3WSmkL/RL0IzmYTrdo0bE
eynwWnA5wz6REhJvXk4diH8JioY4MDZNkV9LOE/wA9rcWCqisUbHNGBHQrUbn10z
RDNRCh6IcpSYtLgGQItGObvlZ0gonALQndQRplkCd+lpZK1X0CKMe0Gdrxe5MxPw
TxEqpy/ktKPwTYVz6cny+flOIShGmO00zjqPm+0aItmhXKN2BAU3OTRrUMqqfgdU
zR3pkNeo6e6ZQDHnPlObJKjxGXVk+8iBGFnExa5MXlXKWK7OP8K09C9ERxHZl6hd
W4UwwC8UgTu2zx5ruFsyEvbQdHOgqx8LvHGN4nJgvu6EGic2yKBgA7yvREaw0nO4
QIQw2DJjIq5Ky4I+99JCwwfE+GmnHxzGE05LH8UpDbGcVa566WCHQ5j3hDuI7odR
MVZvxashrHnYrJCLlaP1sAd8ddASxSo1S83hU+6jfGLPTHkVebR5a2dIQ0R4Ja0t
qKW9ghVQ91qRsOgr4fhbXAhP2Fl9RFXCUlGWG5HF8kcZ1Klk6aJG80fdcoJ2CuSz
yj1mFi7YzHML0gFvG+J1qK6pheAmAVE071wqLw6TE6crqwXjOa5RI7uXbvIA10aX
v6G+t3UVBSjnh3MukI4wTTFAemiVaUdgz+TaWs4ItJz8LObAnd2X0FfNQAahlnjd
HmLtoFdePKYqqNWAlyeDRcykEG5P9XnzpamDO+x/R6DVSUDPfhXnf+0HGy5E9DTR
AF4LRB9oPopiaar7QUAYIxbffIdEHEBEldbutbDIgZo2y5MwbEJK9EWbxUjuIUB8
33n29/SPmVsX2uf+LlXl1IXrHqsCYDPmJ9mv0r//q18kpaByumkn7QKWJR+esgZY
wggfvKcSIzOOkQv+SCQ5v8bFu/Oz8vkql+JnkddI4zqFv4B9P8Un2p2/c3ExOAwH
aDO+GQeRFWf3OyIRmto3YiUHn4uHtbnbMyXNPhrq1/STC86q1ajgLkrnGfcjGhl8
FTSVRZ2T35lKf7wEoyxtygdBt9Rj8CEWzDHJm1Is8bZgcusuqPARe/ISnBDSgUw1
bJv04eQ0zg8X406TacyKH6+8EusRcuET8t4XotQrCGof4GVlSFOcCV3Dw9smxMMs
MWjqkMGpDBbVmIXyfO9GqpWUNwgPgTJYfhSiyVUZZzryrJY9n3drLBieYlBZNY0O
ma+KfdcWjq0oeqZOTQyDz13+48t8uMVrIKSHrnQcWvuIAfm2WgIcW6gUvlRKQlPn
csQ3iU8AejMWH2MGeIlAYR4yvaysU/NvwM7tqv1xHEDIGLkS6xJEbSgJyDO31Q67
ZmP5D2e9Pj6ZK8O4QjTLIEiVzg+FnyH/iL+zYIw5/7+6j1hTTIYfNcNfkby45DKL
I/zYeaQfUPefIA7ikHDIDR1lUeqO/qfcElWVTU6NGdLtgeOR9iTYBNPlEgC6avS5
pqrJgWI+6T64eEBdho3dj5VCGaQVaDqKewvpD0x9iMIAOywvscAvgslVVppc53EN
3y7Zx/OS5Hk12SJYTSZBxFEhopxsqILQOdT6fiu3WZzRrb6QRffGzeE3/20c9+kf
xiEmlAUpqzfiktFJxqXwG12H9O8zBjyij77ch1MNEla7uAXQpZqxGD5VPEKyvP/g
TP0EcJIht4CsGrtZRzcD4ilj7PpbYKRzaHQG1DG690NEuV2Np8uEf73/DvGm6AYA
BSu77Fz8uFPMVqUWPpLe7GwM7qrdpikScFc5mQ0G/8wClgB8GcnUjps07wEGlGmF
pQTAkCySQE2ZRAnzJc04vneOUVlnfaLtTFXHkK8IiCBHgiQDPkPf5LJjnG4WKd5w
Zq1K3cmias6+uAgr7yQV2BSGdqh/zxBA8cVZRDH6m89IKrDm97BZ9V/VyT11sd4A
P8h0P23a9JIlG+Z8jBfguNFVg2BeCa6H22YDMbUL6GDQMF86CgJdWf0BvmyHU7CG
j50E52fqYiK1cZ2JIZlHINhgZQ/2A53w1amRTbC7+VeAgvrVKXdxPX+8CbykJ/eS
MChr+VG5rgVf600kmmmtBff45eDwwcFvxwqeUqLETiptBzQZQ2boEYEd4xq658Ht
pEVLWHw0iZXdmRdOlIv2Ja3kEz77vVEQEjLWU8t3TYRu2Ukw9Ze2zOioiHeAU7Oi
NDYXNYIvqd95d7WbdG0Jh+D6UgeJU0nT6FpDFrdq1Zio5k5w9pQBIWoafJJaiKf7
PwaikHAeYr0xEQz16G6jN1lVruJhtgw4xgOyLcdLQOpy/1Nkwrydb8kzqkAFHnmX
SJcQvZNASzmcOpNzAvfyv1JplSp6dll84mWp9RoeDwel+jwpu+TTIsC5wtnjkXfN
fOawuKUb3phRGN/nLZgYhJTm0g1RrEkb1KbA/EZOHlHNzM0b8wIAbPpOJSOgM2Xq
MAm4uDuuAAXov9qYWDKIVYkqcjuPusE7Xe4fj5i1iE6Kx6g4gmAGmkx25yFuEtSI
Cew+tMter3tmSnlsEWz9xF6TE074/7s2oYTDaDbyX1COooUQtX5Rn9x0WwnsACIh
gPd92Z+EZscRtjCkm/U4Pyv07eNu4AZEdHLSCMoSrQS55JLNmU78zVaLOnkzNsHZ
QgmE5SfUqG+YdIsgwM0IJhrF54Ko0Cii0aKy1ynUsAF7ugEMFyC0+LMBmBwJWRSD
MpNKMbkm+tHQD3gNwjrBO9FV5ysB5Fn54jC1sBUF8Yg4RB2t5e3XQ/EHKpE60rGf
9nki+dku8E6VRNym8yvwXb7F1uS24Y7DaC1Bi5lQ6G/TiAezl0JpempbohDrvR8B
jpmXvkXDp9iFE8ObrhHYlAvHwqwxI+hCPB9wLaLt6EZRJuAD6cod+BmOBJx+U8JT
zyrU8OLfQ+rrlbB7l2uoAalkG+YaNKh7XAcL2BzzlnOtL07qa3cZrFWR3xs0mtTn
BgDglC/3AT6NcVMNPomRfXFVi1L+EahKCJjQBu9ASvhewh6XCgUsgxWTbkfUuNNo
+00s8f4HziL8h0jvglzWCxm9p4G/12V/+XhnSJENCHY6DZo+AUeoH2dsL4JSpzGQ
+ey4P9TgvMxBM1buXvmeZoZrHD+Wquvu4ameJAozOar2QbPKaVW6Y7gtZg7gpAeC
M42CX/Al3Vvur5eT3gXBx4jNqPLoEgqNvXrk4c25xnq3SqBeUwSp9UkfLzTl7/cG
mrjb+HRBWVVazadV/BM362dF0ILaZ6Ez6yvpjRVyeSV6lypr51hp6JecNmxJqoWN
13CHd/2ibILpRGW7t3CorF963G2V8wGkL/6ff4I57D5SZVZjFDpR4yypD9mbVW0f
TbfGVkZYa34CU+DRTAJEL3FjjlZPshlv4JoEV3Hb7epjNF3gJ+fWyfWlJSpnT+Mv
bzwTF9oBZu8uHlq3NaWHo0XhIiEK2P7agLrZxLgX4oySHroQdDpgzqIOAw1VTFhW
WaZj84IxeV4HC/4uoH0qOjoEz8rA8ife8LqoPKJEFZbO5gTnR0t2wv2oA34K/DDy
kreJ+K5DehrCtcxKq/Iu87WCuwu3GGS9ZS51lMznZI94KIVNaJy9ZLcik2IePVKQ
j7zET0ezfPdIqrcgFZ1Zf6ZXhQgbk16JznBvrWFMrLIO5qs6XR+D/GY6muEYW7uH
GoxT6T8NTvdPTxui7IjDaqB83QzWp9pHnCGonfEG9Eefv07GfDERQtEJXmCeEZB/
lY0O7IeDmHqsqYlW1pwO+VYVsvLyev9RtaVNIjhS5KSHOb3sr+PY+4RLt5wQAVGF
xfxpD4MYISGb/d1fwS7kSUh6DWUurWhZ02mnag9NN1lIRwK6DuU3Iq1udpx9nCoR
AeAv1Uv08ZFe4cGcJJz57C+91bddYBk8pixxMEyNkIe7tlPnNZEY7EiCb0f+hQFa
ifMRELG2QIk6JGJ1EbyGKf0TDNPktld0KmNhvk7S6gwWDTJ1VIyYz2d8UhkezeSh
OK4By+SX+hDQnyS9an+BIKjj8ERPxXH7XDNtgso8mA7vK+9lp4Gg/kndgryGLYF3
p8hbJHbEcbnGhHWOkIgRoIxBw8tDFWIzNt4IkFh5qJAIro5P9VsRItaDhuJ9YGtH
Q5Uwm0re1l3u6jGGn3XT945JSdBKkiAd8RCXEssOpPGB/vrlbGM+9b1n8LNJLldd
jbWLZvdPtSBI646+5Yn5JoCwJMAcMJ8d8BYA4ypYwBQihHlyOxNA0rw4aqMG1YT3
MenOOrn9/17qB8pZ8OAzVl4okaGhT27evTtXn7UxBVD+GuspoNrOxu8CqsQnjv4O
XotWW6va9hpCizbCgnuNySCbhOb/kQTdcer04ES/PhOEJROkjOE4Ogqz2GecX6FC
HREFfJQhbmKc4c+OvyWd34Oe+bWn4N+SZUXhAz96r3Txzw+lyDicXMwnYNwXA5Rs
iFj55eDThZJzw/gX0qXj2VWPq9opXGItWohNKfreedhAVfLitRvCbetPICUqjI9l
W2Qp7HMHik2CyjO8TkoKVFd/NMVxliYC0IECFyLf1d+1Y0QK0UcyUuMcqVJlsveR
N+sSATyIOFmEzzheperK1t87JtEANeM5S054RpGZWMgFI5RrdwQUD8ix3PdQ3dGe
UNCc9nLZzDzyevy8r0wnxh70rDBLZnTU6ZeYOHgZMZPs3ZRHpse0cQRi3FTxgwaT
180EKlD3ylUMeveAP/O/pnNdTmu6Uk3zot/z9UVEgX6Jjh4cTOiqbr98xlAMwWIr
svsfC+a9BEIF6NPZxxjO1OgVnw+IATMFWE459qKYS1Hr+k0mBb/3u/r99zHvxOsb
NN1zqBvlbcqOfPXi7Xic0nBSvTJLVqX+CpezjMGpa4U1Z3cKjSXSqUUczL3enHOn
0AAOhm2ghFP8DEWYTglrxe+dd5JPBj2mpIRP8MzEe9O/4HJtKtQWyfo+/qTdR9E9
mld6siXQyhmYgtpx/RQKKufmStvlZm0EgwVMW9SHXiL7+Hq3H++hmfFJM7gMVb4z
MIS5pwxG5ynzezMxKRolH6YMVVTrCzcys2QUdRCGF92KkqddR1bE7q67oVvBoTVc
zURXEifP3BShJL2GK3u4s8lxP8tTCwW16TtCadG9bnI/Wh7pwbUKoztGgxXtTklw
pxcqRe97IKoim/PUnplD8LzPnkGxQMuaBSKsNZBG/MG8rqpBQXhCXfE7Zs0eJj30
Ac4+BIOtV6OtkIR5XwfxIGiOO6JymG0X483SNmw9I9NMrvyi5fMK9o5c63Cm56tQ
bpz5Ngskt3H96M3AS4haTfSGE7KZ8uf9OfhLmjIOv51P98Q6FtqeFGjf080wwv7w
Q7hFr8O9CgEmMKnhw1Qo9agxCaANhlK8cPDZNxVTK+PDa+WUK0hrGK1bcoMwsXeq
NHIqIqRoo5kcPIlhm4aEQmGDhatCNiVEoq9A4m16OlPp+zZGejCP6WApQ+6Q+g92
f2wpYD29k8f5md2rcyBnqNsAzL9lRT7OJqz7MfuzQiV1eR81wSEKyU/zYjwucqE8
0ye6hJv48vv6XF1Jk6De+gy0VeQKYAHmTFBI+kNP6EesG2mm47ljbQf/fxkZPDyG
rJ4DTw44Wp5vVnCZ43C2Ob/HcPn62zE1XZwv8hK8NCmZjQ3gPhhOLc1h8co6Hqav
bCvJ/x3BRhK2Rw+AZaYlYuP4wMYpeR/m14IKYwXd51McfhmP0NVfFHjYJrf9r0Fp
rrUN91Jophqdm7vXaQh5dgAd2rByHC7ktRoZ6SoZN4KrOLfY4WsxSURP9O5xOrT4
hdAXzz+XoyU6osdJQLPmmQaViaFYYIEaCTl0USgMj1ARzqN0IIFaCf9YeAg0c9zR
Bie8qrKuKVViHb3Aum+3zpsb04fvdaAebXKb54zSf49RbKht6ZSXkpu8ktYUruQB
waOH/LGqIel+x47rgZ92bjDwIOcW6X6L8BhmqF/n9zAk+fS0PbBx9rnxvk/GRowo
CKHFvWLw3lHWHi65CBejFGnoA8NyiTal3JlKVq+Ltc/9XQ7WjwzeTuQDTYuY3ylH
m6a2mJGZ3bXenJEhHBtNbr9qvmwZa0GGzzch7Dpcujr2ARkP0/AWDVsYEAvyvbT9
qk7iAvGPunSZjGa9iPGJjl7r/Ax2QNDewpmmEFfjYsj6HpncWXsRIynhKd4EfQTw
QZS3V0+G3Ctq5r2c+3yywRnqTAX4gfIZZfKruWEy1ut84ycSaGwcQPbGrGVOe6kv
1k4lIBxVCZyXxd9+u4cosJ5UvDFChV1A3myx0yBOd08hXX/BrvHESpH45zPbFkTr
XHfnxDfLh5LViinhPZrKBd/77lHBjWdl2PLAd6fl/BOxEQB7zB24tcoAFk3EJgX5
A04BN/hnVXt4+YenfU6B3ZgG/l1NqrOuDmbYLs5nGytLwHI0czoHBDFefpVQ8U7M
eWa4kb7AJqmspjO7yTvXyB1Tz7fRiy2rTgZz2X9vN8TEEtjdmn1rS/cLlowLSFce
RFU3HDLon5gHWzdn1B7h/oTuNCwkNcluLpgSzNeXFStKhx4Yv+/pqxxTXIXRFHIW
ZZ6jhJ/mKTMW9zI0P+UHhKD/LG8oNsGPnY2cRcIx3AZRMAt406Bzz8/BuVNgqpDW
K3ooSfKdV+7vVxDXYZRbguqeKOfzO0Xit37jQzdLK4KxD9/O/fjHPal8kTRMfgdf
CYUS1MkRJPd2d9jlCS+mrL/CzIR55ZzMbSTC6UQRa7GNkAp1Nhcd1Nvm9/Ei9EHg
1/eqGcpXY5SAe/QTHg/y3HqQ10Ze1TGBK6llDavr6dAbQBcEzMIqp2XIRhbkLYac
/mHk/S2apItu0P9xwGBGePkTy+Ca7EjvIHcbM7iXvJwGh3p2vEm6fEwBcxvF1I3Q
X+dseoHmdbZKf+iq0aIoq7ZkalpZ3ZDyK5dIzDiqwAzw0ytLe9oKSojS44X2DrjZ
flIaZvTGpC8dBhCqKc1GFnoIIDr6o5Po+wLnT2STYmQGs4fts4x+mo+MYDe3QrLi
MMCoXGHVD+TpF0PiNXgzL2nIW4C/ABA/sJkn0BlPhIL7pAWksRUjP88g4focE6NW
0K2cnwQ2AAnyXmCtsOv5N/03Kmlny+ZdAWK+DlbH1wGdIUKbjfJyAnK+q6tcRvfa
3TZc+ZLBSmPgkKXIyQZz80pn+wzmtxnTJmvGbUczenIBjO5p80moCCu/2TH5e90n
ZO2fAO6IXg4PhCXp+YCK/vxXHN41ppHbQE8j9m4jrdmNfE7ckQ7zHkeGXTz5Ockq
q8q85IYEHN9pMorZl/3R73M59sMT/QYYehX76fFrmPwSkGg6lXVLKjY/+EywGhPv
sG046mOpbmRs/ELIxzVc28M4h1N2N1kUxHwYjBFHe0DV85WEqMVf0mdm3C171kbO
D0TYD+75TlMMRnkKxuyC9DvwJYEGcaef80tURbV76spnnKaQRuLrgC5cOEjnhyq8
EaXyPw+tssBLNu1QJpvO8PlK+/tAj/JwaNawMsdD8fjW8FuaDRyKmjO78HGF/fhR
7fL9u9P+J7mVXIq2Sil83/w6auiucnYbEBTeDzV1P3DTA1hZH4LT/wmIinfRb0iq
PALkOH44G6fctW0a0m27XskOjlguKMz0B8WH35/ATWvxYDybzHVgzYbzg6kQVFQ0
MkqAmXTWImVSQVnY/pdBkHpSAueTxADPTp3hpibLlHOCOAcuiDTImD2iUyB9gAN2
sW4/JIennheOTwvDw5KmvdqMynqoNFOXuxlhT0EaxBHj6YtOdlj+es7CmpQndi+G
oUYBTAgjmeIcy+dTjU8c5YzmYHLOZV5fPfdr1kjP65+5ite8WCahEpi+CUCp00VE
S2WRrcbM5H9zbz+phHQFWLmhSCZcNxE0tebCb1yraOraY4POdhfGBTTfMRwqraXV
X6e8dDiUqTojD18AcQzx8etEJ7Dtd76e/PqT4PfKpYDy5g2/ocfN1WdPltm2vNHK
I+cECppFE0xZk36tTuYKJdCPE6+znViuOLTRG586orSkBs1RrYu04uanpzUfazOR
wMhqaSmK3uJEV0mqJ183H/cY+Ma2QOHylmlzX54ESm9800BPMi0N9/QufBKsC2xM
P5eATTCjcb12TzS1DyvCvdv14NWdTDZ4CGZWq59k5tBNUjFDAGkx3I+vKfb0y/FT
lusYwWCSqpZIMoh1RKXWUVwgDmZHs5c5VW3UzztRknDiOXhTEJhI7vDTQ2LZb2Hf
FQiJI3Ww4DIR0Pj3/LErE+RXKGn3Vpg4vVjgHLe57mUUXW4XQeylz9R735g5Bwkt
uLp8jBjfpwzscxeaTy038p8UdLVHH1lpcerIIAGkcbPNnQZMK57HKQZdGQ1zHqCc
HNWni4Y+RrDUbWdlviZPVr8o1TRNykf/zbbOsULii9Nahsp03A7EFQfQAOW7gCUn
feITc+Mp6C4PglHw1W9NP1sV/i6AYn8iFzAww8ZvmOAkBTRfXRJT6/F4imfAESh0
4iSn5aJDYPM9t3YA7WqxaPqw/lNtcmv2G/chjlPfl9JNULBOrU3+CIMtund4FuRO
yl3PXvi2aTfHnqFy5gj3zCzFlY/HHyo+VViNQ2XWYmtwBx8sI1oJlFiDevV39IwO
B0r0wV1FH5Eg8kqAFoPmRd8Qp011zqkqcgxgopybTSdfHaCbBD2h63wlEPdIzCdS
26L3sN68KlKciV9ZVC6USLP5Q3wpoxo9jOsJ7TBzYl7SfCZF0/hzn6U5PHJgQU1q
3Of1028dfiAm8iQw0n7lEGO76FAkYylHydwnN5tWe+FHmcOfSgttKjcPR1mgS71L
U6xabRYaahYExaerky+mJyUDFFxRKqd6+TVMicuSqJMvzy3gwTANGTX7mhvm48rV
IGu2g28HnT0bUqy7CM4ylVg0dRvdpPzhKrmDPA4S7tW5kigDGJAmcA8VF1GsRG62
H9dVwm5uyCIgvSygJhRXHGqe/fcMBztg/ssSZEKynKsSf8w35X5rWXqtErQVDO/n
kjlkaARMhvVh5bEnb5RLTichOdSwzVDcGFyjY5HXiP2cAlMM6R5LKjT4JQ6TmaRz
ub04Rq+LBCX5ly+qd0qxbTUzqDxTIC22JgscMQlbvGgVKsWa4YmCAR2n2EXPULbb
FVzftAbFbmDHmq7KPaVPWBL4LfyyMTtDzKiiSbmj0TzpprfLz6SAm7pPGSDXJyAZ
adgHTOKa3BvVpFKBy3qt5Z/VOe1DDVeR+oLdxlywSvTYc9I4hO/xIqDlKKLWRoQO
e2qW3wz3dIvbSI7E3gy3g2v1x1CysPXBkCaBdgLa6zKXslehjywOYJRWL6oIb77k
4U1/QRrggWnALIUJ/GWvjwIPW1a1dZ5IKjZwtzHXvLZiMQccB5jrW94Pi9jIfQBj
As3y13mKSxx56Sui/mrxfnW0KPsneLhgNWD2QlcUsi3O/TVyIKOCXYYpX40/13Re
1/SkyDSz5Ju93tO4XpO6Us4fouVin0C75kIcmOzq9G9x5A+j7Zl6OINrGt/ujw1D
Brzfc1kJGFpDG2D4Q7Yqu81fL4Ow0VIyQ2yMndThqYPB301my0TkDfJYc8sL2rGP
EusGZBTCHfHkzSqHWUJlhMDTEGEOYhnwaALY9D2u9XwezHOQpaM5sFmKV3G9mkB6
zWqkLTD765+tpvjFFSICRLTImmxkIg1z5MqtVqQagDZVIUMv2el3iIg827yAolm/
Banq2vWrEbUpJvbIuDqHKpLZfSChmAzpqhqcy35R79tk3TeNzRZ6kVwSU/lLRjB8
au4IXRO4upW+lCokJ1p7b7ARgFUuG6qTQnP6BC/6Kb6Y2wy7vLX8CdwL+2empE/Q
jb2/R7aQn3NbSkYKrTm1yDJnbb1BOolBAUKk0/KPV1PbLohOZn7tbIgeFqy3ATAB
50LWrvbgatr8bwTqn0Epylise4s2gRjYZjF1gGxIyvzyI9h9cJNd5UTKexR2jdW7
iW5XZ03+5nRnXtHC9LkrTpOjgAFFGd+uEBRuOs5xpjdSyyWRsF/s6fLFsxBRETx3
xzx+ibBUhYjk3720hSCl03gVhqkbJwjXZYEC5eTuYGl3SXul5zfi47RlC8Ip8A7Z
u8EQNfA9HFjWeWk9FuFQXp8yGAC1lFftBov9VLuRnX+op+2/16sQZIGiP2E2e9BH
jWvjQVUmilkNunNrgBYwcWbQnSTvMDH7TNAYtqoxB2gJt82WNgVc7PBVE8rOrECd
gugSHDZd/x7ty2rOvgnymMw/1rpL/jVGjP6mnufNb1omdf0e7ZiuP3SeMZQixLJH
pud/MwLRDvP5e2dSX7fmJXV89iRrYnHCfdamRELIlLXc3DJjNFVvMp4piBw8Gv5w
1qzR93ZRYhIHElYqTWlGLKxGMzgOX/HfN/NPNrDBm0/VK2H/i2vnyIUvbUDDkWCj
X/PCssbhSY28+rkfBD5jpzVZpqrYi8Tgk2bpxP8rw5sl9M7zTXWEDoqIIBkpjiG4
G/AhzJNXRMsbH2JPOfHziMOzn1QgUoaqVdfQE3OwxV8TscGEN1ynfRwwnANeSNma
9nHYfzsMb9KgE7d7lPbUJ6/+BtY/Mu/6sL285/Do+RougeeRx7Xo1OBXgAxUHBUi
WZGii4yWsGk7KB1Dxk5BEkWeYa/L662OvwAgaJ+usxSNy2HNoIAlrgR8Q2AWTiKj
0xB+0pJU9kRJIMgJQ5GJAR7tGJAOl9Ew0x/Vs9v7odvLP0wFmKXl+c4bZ5zqrRX1
gi73PKLBwmAax+/G0Jzm04UFUMmTGEukWZaRqvwhD7CSkcG0PAPp/agqrE5MhvHx
GdHHi4NsMQWYG7473Cjp94YIV1XeOie4Io+wB5MSvvbLn9U3kJciEPmEThEnoQEC
dE/t7HRycAuS0q6XHH+yQvQAqEU8HYftS2o2smR8/MXumLA1fzd5yxu79bCkvJ53
PJETKhmjKNEE84i8Ef207kxOl6b5VvRfJWXpADshuoW9uNfunH7eo8oz0Yo5wR3Y
sgHA2VChwKBTMwJ90Yw+vWoBl45hll7CbsQ07hh+fJvAyeNC4OVj4/19B8zgx58Y
l2gYVcI6X5NCBNcG+DNMeGIEKbwfRVPgmgnxKQJz0yeUmnu5UoDD0xTIqpV3cfSf
RXx4WO1wATnYHvB51jcY6hTtIpNAi5YaMNWdenW5UwOqNRnlCq7HhsOETL3K/POf
zI7Z2+sYfCwfANn3DiZxNtH2BMB5pmujT9t8ODt7Wj4NFA56TR+Q+oseOYP27acz
AvZA5zP4o88i3qKmW7t3ipqZ20MgEJO1kI3E6JLheTvM+049Y89K8UZwUav8jJvU
z6WTxMLQmChUss0Rfa7Okt4f5uLZBxytfq/MMGQ1UHAuHOQF+CeNPoWdz1HQ8e/b
6RAnU4Xflwd/TAXG9mhUThiZjFK1lmCK0rIu39xf8pq4uliWzL/NjfLmDgvIOUoI
7p+dXSUg4sXL0EMXzmoEAlaYkdk37d7NvTLFKI86+2yLlpHqehXRxy52NsAonhDS
RxoNjgXMRu28XEQySaYjCtUaEgYbchrzkvuVXd6C+1EMGaP2Dp9dY+MoJgQ5Q4W+
l5mBTbQ72J3SE9sgO9etKV5b06WZ1nvQpCXNpeZAGBGKPIqX67UnfR3dGSrLm2gp
LtQ3xQkXk4YSKcJOlpbbndTUjch1ySEysG2gki32JHNWOwly3WskiICapJ/GsD+V
Oxs9Uzp+150mE24bjc3vzr8ea0iTa7xkRt0OHzKZcYBcCaEJ8+f7mRYGADLEgYP1
2R7Ctl8sZADbPS6cxxcL8JKOL15q/Cknx7pC4PwFUeDG3uqLN/+AjL8K/xRXEBGV
NGrLDWh6LpSZ5dEsK0NxQnwQlzQR+H1ynjvc/EYXbe/qlBKD5E6GQAco4bSTpOtH
RjEAsvv7MWE66T+M1sSDR4wKpmPEkJU96/nEoVYYxrMOr8yIl1rF39EXOH5bnSZt
Pg1RaPBu116dYwKUaJKEZxCHOL+8gjb7+CCN+Y8KBzgOVEoanBsjgGiPGZBBaNzl
aknD5QQDzIqbN8WBASHp0zGkVX20kwY8epllmrFyalb8XF8QCEucCQyfw2u5TSZJ
cMU3QYJD4fbgq1N9Ewxu2G0jZCr/RDDfpcHoShruHd0dtiuc6ajsKV4MNREn1DOF
y16j0Oew8e1iW6CQnnmPbf3dp76cZUpX0vozQY5n5vnw7+EMshEtG0iG7XWCTK/j
/cY+l9WAqWD2n00Fw4xjTa+BW0mjOqyWD+IlgavK4jshJGTi2Lp5Q9260XM6ztSs
crfI/Xsd2s+efAUN1364Gw/ZPkDBGfhTLsEXZY1os0AMoqaxWxIo5jvdTlcDMuHL
wP1rjMZmr6qE+vo1/54Z5wsAjB7qpuWKyC7NI1o/10DWe7NuA0GIRFMZaDFc+s7f
sNb8TDPHi/RCyGUuxA+vZqsDxvq2upeazByn+FndygnAS9e/TzX/sqkcXD+xLZ4F
0BiM8wjGll1+Dtdr34+4mnzhG12H37vAkbqhRQ+lD05MfbUdqCbZBbV3+jJNUBIQ
+0OfeCNgYuTJnvMxXflIjGKu8NZpx9LBaHinOoIMMH+063mJkQlrm1fV7urQ+6qT
82a5w8pN2qpNS2YhSKf+nCOkIyjdb+V48LcNwrtaw/q/239ZNTMh56KNyWN9xQ7H
kCkMZbWb6Hy9p96HVSwwFiVdzKyB66lxqfs55eqQm0rdQv0BrYzBuPdinXRBKrjI
XkGcy85FbsmDmbyIm/nz3YBv68xsk2NlRPjyGIaneclmr3B3LYbZnwAIatn8yrzD
Ww+zg+d0r7KEGMklrBg+N7L1pDqgBKvWHD0pRthqMNtm0VZ1AJv3pZ+FjqbZJiyf
ZkYsp7mTEGPdkEJpNwLRv2V0p73RRvDIjtPL9YasfKjo3xvXVTwY9gVKc3PZpElg
7oqk0fLJQL/W9Bp4WU225lr8OnKkh+DHatVL/0SYrJIvttBJUfEpiZgngcHY7MAS
1wfpF+N+wtrcsf7PmvxBjFBM09mdIAQDjN+T16VrcKFF8o6pMlw6n19n9KEFgdgD
fZU5o0bYzIvZbEFhYWo44+xMjP6AkLg8RnpCS/dBYBBI4aW4UPu39TOI98OD9/3U
iBjCBub5JjLAZXigc/am6/KBb0dMKo6uycQ/QuuqIUblFEkMypV8uVwP01KjlGfS
tmaYAI/nhzy3gFpsND8vFTdqLuqkj27kCb4MJyo4oYLIfrO/zZk0gSQTYzCIr8o3
Xo4R7/l/0i1Y4uEqOnjrteoW+S7s8C0dLr6cHYX4Wt/04PNbdl0KGqYKsO1u0Qmo
VKm8SOGZS5wO6HSjNwvU052qVi/gQGuqV95gjtjHcWC9iERPX3ncc9QCrrjXhlMq
ShGbPWnRQJ/uR/l4XVzJNwJQ+6GiD8+uLM8QqDg97II3UBrtNN7qVbNVPb7T63bu
kobY759172xo3tIJht7EvtRNiJmu85iCiI+MPmgSbConF+HTk9hLxMkJGTJdBaqf
NWzvEkZHcfWSFOhzUhet4/ooXUysCpAG+Feog3UAptMcTmsm4xNWH773RMtCgaog
0UK6BqnF4pikAcFlLHPXdGNOkA3g/3piH5ZZdhRPE+qBUuQR4fC5baOaTi2G9bpr
OET0ZSM0PR318Z6QsXY+HrW3PlyIcLU9kaCUuBQF8PUr3RRwKUaSQq1n8onM98se
RBJNXQgIPdppYr/nDuEC/nAD3CrLpbDFbWaneUymw4tei+w2kAyClsiT00wWBgqW
A/YetBRnmCWeNU2o8LGobgF5OsGfb4qsxSd+bGR5MEjQrX9xK42UJuDeERq+g3Vr
xBk6LqqF1+z1K8qq2yeViP8cIN01ebdSvkt2vJXUQobiwyLAm8Z+67H05Ffj4v9O
1A/1z/DAk/qXG6CUPjzU+ZVyI0tkK5dpTJ5H6+NkJuPpgncVm+liJFd0kNYf3ZiK
/tDpjo4iZdArNhGvoCMsGzLuXsh1VGD1Fvhs2i6TsYDl7Bap1z+0pUSXgfENXM0D
crzctURDCdSza+J01Ysih88KOEY+ml0nRab+Red8iHST3tLBe7PInFlf1L+K2AJJ
L+htJuI7JQKUnzTdOVbitMWws/8IJiHZWyhz6AY3H4sFPKUIpfQaT+mvXgbYOPoz
I9bVlgGFldNGGkOZkul5gsWGVRUuEoa++gmDVIfv0CsMgcv3Sw7IeED1U8pujYGu
Zn0RKqEiQwDiwbqF/ZGegUZDKPfuZEArHa6znCPUdHL/b4R5PG0pNhDImLLMrGlx
3vLA7JRO2UviLoxTYzPRdOKD+ptWXjjNDaqrTpV1v4MHisbKK2U4kYXk6rACPGqf
S5uSPEYRFYEWWzyG9ihRzZme2q0Is9ecqk0rUqGI40yrrVXpl7fknc+VUGHNo2Mc
skqJQwXF7cUeA5MW4IgOMeckyudqYF7rGmZVPLYGnN/RpS6JB3YYuNcJzEohQx+d
J+vARPVXFP5fWPCDTaLI2s4B8zzEZa79wTS4opLvwM7Yq7wGOu95G1BZU7N843Au
k8mD0s/2Yz2B7MzGqk7aaXrttUyUbA1PTSs+Jcxr0vCtdX92tSbemtgrt4Y7VD5k
nzzy5I/Z+a2IHOai1fuGTnx0X9hLKMRf1k63EOBJ5R/I1gfa9I1pNYkzYMzSchhQ
MiZuORbV/E1W+A5iB44scBfR3ixW2w7Otzr6pLcl61I+gYtmPKHbV6//YlY6Wvcw
Qr3rfob/XCQJ9vBVH7TiXiMG4tN+SwpOBLNuU4jGIs12ddd4AtLBrgTzTYxhu0TI
31l46aHRSxl28jD8jAnzk5ZLfdM10H3OcJhX+uHB82N9ku9nSb3/htKs3OD3JCNz
+636VscUxq3bYsGPYLUlshruGYYBfVai5LyUVHhvhUvKJhfVopo+HXidKVhTDoBE
SyU0/fJ0zPvDsrSJ3+GT3I52qyxX3BeYbXIqLO8Z7C0joLNxZYRl75/UqPwzDMR5
ByfYkmvMF7TpXyyU/G6khO6P2Tw+Bh/zZ2258qXkX4NhjVLlQjqOWfmF6veV0u33
eKi+vJk6WeoEn3zHwSvSI9llMnwLxLynFZujXXpG2oDFjb7tdy09XVUjt/8RG4eQ
pxBF4j1jZeuvMMiwP0rnY1ZRGruFbA5mNm7cC5tzd5EpQRmSakAzeIeOwoLcU1Ap
5Ugatg7rj2TSHmx97e5Z786GSuJnY27eO2F2BoOkaoO0ggRvwqdAkDVcSC/Pqvrn
3rwcINpefGLzTd/bSI+zDsyqHfuSfKAoSsnP5b30/YhN/EBEJX+slhDsPrE4adb2
eHyVG8nEMalPFdyK/8l4ERGFZGX61eXrBUz1YDbT6bso0ahLwHrM2NK4acTxbXgi
0ymef8jhnydqaS4QFQkg/gDXBcgEBoNfpH7PvU61csXEmN4GbNAL8STTKnzGv60x
fD9U7NHfmrenVJ6RfkAaQhs+XlmNGQqOl3Ch0DO+BxGCBXykQS4CLiumkJBWopcy
tN8zc6D4CXmNFsxdbOFA/mL8vRtUjRCxfCvXgG2APt9nx9jQXKZt5+XBzkxYJMrn
hCX8cnlHDTe2b15UGJsNXEPotkn5NfdvBMx4xs4sr9mOf/Cj+OPnfE+o93bGglc4
2qUu208hnclNUdSXihs/JikowUBLmG8b6RYLDCaIrV309WOC5gO/1W2vB8KpUKGq
H4hpzmiH8hVtWwAA3DbVViZMEqKnspR7TSEcb0vq/UY0grWej0G3Fssnb+jbingU
hdvkV7pT3qTV5hfrl12wvulWhvnVlUDlmBqzItbPXX2c7UpuIXdXU/AckBL2CDYa
ncubJCBR2VPHYuBCIWzgMlGJ4lXCwc5PYUuTWAnz1466FmYJwvJ2eXQt1cDdThmf
0IWdXQNORuiRTebwnyyq9Z1sBTWFL1Rasoe651U19Y1b8zvWZRQFGz5QJDeSGKil
Swd1uO0MVmdB6QmmCMd9Vi6qTKsT/rc2JRX08w0KThFoRfD3suej958IU4STQqaE
qgZ7r6l0QfLdWH/M/9Kjv0/nzYhEt8yYGo9Y826Ks7UTj7nT7HQl1YPSPEdWOuub
ko2u6pl93HQstGRJg/dj+48PPd4vGyYqlMcqemiABWAlw9dAXPEuEsmXwFny8gzz
afp/aY/4dqS9bDab83p65lUVp1ycx46hshbfnHLZB8WAV8SXoOrVR8I0gm/I3a1X
HbYeMQ2wz9lE+dJYAGm9MiK2Jv6cd3rAXkmbo6nFmGYHiGtGUFarQNtwa5EWn5gM
F7N9OCKGWf44tKIJIj4msRLcI3X59gGmXp+Lng3iIojClbHVhe2UrqkCJb6vMaHd
2mnVvc2jxK7Tsk5r1eFZaYQ4hphfJxyyiPuhJO+sxPVYBv3/Hh5U/XOSoRcIiCc+
iNyQzT2BLwJRAnKg2jjBcC2PN7aNUILNbHYOMzT6AmyGHPLi81GvUeJtywxd/3H/
YHJ5CEwOlYqvAITopnCnOclmwlglprTfh119JBmZsE2BkNhhzti+GB3b4Xypwet8
r7teisATGa7zjdUxaXmocbkiWs8rsrK+SnfeONdcyI8SK3haXkJXxsSQ139eatAH
7TEqOLTNZC8skoQkVhf1RobK/rBSLscbBqON+LdSM4E8nM7L24E1jlSKNEbJfZsg
cw1aj4qJ1P0X3ClEJLDimZwG2E0VxmcDLq/x5ate/ftIwUol4C7FftS+Jr5W4HIz
h9t9QuWrMA8lVKIEZMmG6HVAAdfXeE13bbEqSspkuaLxHBPR4X+sBS+Ti86tdzcs
FtvSy1kubCWVsPTwxqqzH3+NRuosVE72tG/Hy5xDUDUdT/2laYOIOaQuQhJ0H3z+
wPDKNgRJ66CN4NSpf9DZz+pSzuPpFSbof2R1K3o5oDT2nFfFRZFgIeh/FSSoY9E6
1ZLVO6X3vCNACQHIcDbl6Q==
`pragma protect end_protected
